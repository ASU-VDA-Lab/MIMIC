module real_aes_18107_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_0), .Y(n_606) );
AND2x4_ASAP7_75t_L g852 ( .A(n_1), .B(n_853), .Y(n_852) );
AOI22xp5_ASAP7_75t_L g144 ( .A1(n_2), .A2(n_4), .B1(n_145), .B2(n_146), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g113 ( .A1(n_3), .A2(n_19), .B1(n_114), .B2(n_116), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_5), .A2(n_50), .B1(n_204), .B2(n_213), .Y(n_212) );
BUFx3_ASAP7_75t_L g545 ( .A(n_6), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_7), .A2(n_13), .B1(n_121), .B2(n_196), .Y(n_267) );
INVx1_ASAP7_75t_L g853 ( .A(n_8), .Y(n_853) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_9), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_10), .B(n_143), .Y(n_530) );
OR2x2_ASAP7_75t_L g475 ( .A(n_11), .B(n_28), .Y(n_475) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_12), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_14), .B(n_219), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_15), .B(n_224), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_16), .A2(n_83), .B1(n_114), .B2(n_219), .Y(n_577) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_17), .A2(n_46), .B(n_130), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_18), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_20), .B(n_116), .Y(n_551) );
INVx4_ASAP7_75t_R g232 ( .A(n_21), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_22), .B(n_119), .Y(n_174) );
AO32x1_ASAP7_75t_L g574 ( .A1(n_23), .A2(n_127), .A3(n_128), .B1(n_570), .B2(n_575), .Y(n_574) );
AO32x2_ASAP7_75t_L g609 ( .A1(n_23), .A2(n_127), .A3(n_128), .B1(n_570), .B2(n_575), .Y(n_609) );
INVx1_ASAP7_75t_L g153 ( .A(n_24), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_25), .B(n_116), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_SL g165 ( .A1(n_26), .A2(n_118), .B(n_121), .C(n_166), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_27), .A2(n_42), .B1(n_121), .B2(n_122), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_29), .Y(n_162) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_30), .A2(n_49), .B1(n_116), .B2(n_233), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_31), .B(n_532), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_32), .A2(n_88), .B1(n_114), .B2(n_122), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g567 ( .A(n_33), .B(n_516), .Y(n_567) );
INVx1_ASAP7_75t_L g179 ( .A(n_34), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_35), .B(n_121), .Y(n_181) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_36), .A2(n_66), .B1(n_122), .B2(n_581), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_37), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g477 ( .A(n_38), .Y(n_477) );
INVx2_ASAP7_75t_L g486 ( .A(n_39), .Y(n_486) );
INVx1_ASAP7_75t_L g473 ( .A(n_40), .Y(n_473) );
BUFx3_ASAP7_75t_L g500 ( .A(n_40), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_41), .A2(n_103), .B1(n_104), .B2(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_41), .Y(n_489) );
OAI22xp33_ASAP7_75t_L g501 ( .A1(n_41), .A2(n_489), .B1(n_502), .B2(n_503), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_43), .B(n_569), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_44), .A2(n_82), .B1(n_121), .B2(n_122), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_45), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_47), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_48), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_51), .A2(n_76), .B1(n_176), .B2(n_516), .Y(n_515) );
OAI22xp33_ASAP7_75t_SL g101 ( .A1(n_52), .A2(n_102), .B1(n_103), .B2(n_104), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_53), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_54), .A2(n_80), .B1(n_114), .B2(n_219), .Y(n_541) );
INVx1_ASAP7_75t_L g130 ( .A(n_55), .Y(n_130) );
AND2x4_ASAP7_75t_L g132 ( .A(n_56), .B(n_133), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_57), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_58), .A2(n_87), .B1(n_122), .B2(n_142), .Y(n_141) );
AO22x1_ASAP7_75t_L g217 ( .A1(n_59), .A2(n_71), .B1(n_175), .B2(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_60), .B(n_114), .Y(n_529) );
INVx1_ASAP7_75t_L g133 ( .A(n_61), .Y(n_133) );
AND2x2_ASAP7_75t_L g169 ( .A(n_62), .B(n_127), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_63), .B(n_127), .Y(n_536) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_64), .A2(n_124), .B(n_204), .C(n_605), .Y(n_604) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_65), .B(n_114), .C(n_534), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_67), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_68), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g607 ( .A(n_69), .B(n_238), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_70), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_72), .B(n_116), .Y(n_198) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_73), .A2(n_93), .B1(n_176), .B2(n_219), .Y(n_518) );
INVx2_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_75), .B(n_199), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_77), .B(n_127), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_78), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_79), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_81), .B(n_137), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_84), .B(n_534), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_85), .A2(n_97), .B1(n_122), .B2(n_233), .Y(n_542) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_86), .B(n_516), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_89), .B(n_127), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_90), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g494 ( .A(n_90), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_91), .B(n_224), .Y(n_571) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_92), .A2(n_149), .B(n_204), .C(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g237 ( .A(n_94), .B(n_238), .Y(n_237) );
NAND2xp33_ASAP7_75t_L g202 ( .A(n_95), .B(n_143), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_96), .Y(n_550) );
AOI21xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_847), .B(n_855), .Y(n_98) );
OAI21xp5_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_481), .B(n_487), .Y(n_99) );
OAI22xp33_ASAP7_75t_L g855 ( .A1(n_100), .A2(n_102), .B1(n_856), .B2(n_862), .Y(n_855) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_469), .B(n_476), .Y(n_100) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_361), .Y(n_104) );
NOR2xp67_ASAP7_75t_L g105 ( .A(n_106), .B(n_303), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_239), .C(n_285), .Y(n_106) );
OAI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_184), .B(n_207), .Y(n_107) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_108), .A2(n_240), .B1(n_259), .B2(n_272), .Y(n_239) );
AOI22x1_ASAP7_75t_L g365 ( .A1(n_108), .A2(n_366), .B1(n_370), .B2(n_371), .Y(n_365) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_154), .Y(n_109) );
OR2x2_ASAP7_75t_L g326 ( .A(n_110), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_138), .Y(n_110) );
OR2x2_ASAP7_75t_L g189 ( .A(n_111), .B(n_138), .Y(n_189) );
AND2x2_ASAP7_75t_L g243 ( .A(n_111), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_SL g251 ( .A(n_111), .Y(n_251) );
BUFx2_ASAP7_75t_L g302 ( .A(n_111), .Y(n_302) );
AO31x2_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_126), .A3(n_131), .B(n_134), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B1(n_120), .B2(n_123), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_114), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_SL g516 ( .A(n_114), .Y(n_516) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_115), .Y(n_116) );
INVx3_ASAP7_75t_L g121 ( .A(n_115), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_115), .Y(n_122) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
INVx1_ASAP7_75t_L g147 ( .A(n_115), .Y(n_147) );
INVx1_ASAP7_75t_L g176 ( .A(n_115), .Y(n_176) );
INVx1_ASAP7_75t_L g204 ( .A(n_115), .Y(n_204) );
INVx1_ASAP7_75t_L g214 ( .A(n_115), .Y(n_214) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_115), .Y(n_219) );
INVx1_ASAP7_75t_L g233 ( .A(n_115), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_116), .B(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g581 ( .A(n_116), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_116), .A2(n_233), .B1(n_601), .B2(n_602), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g140 ( .A1(n_117), .A2(n_141), .B1(n_144), .B2(n_148), .Y(n_140) );
OAI22x1_ASAP7_75t_L g266 ( .A1(n_117), .A2(n_148), .B1(n_267), .B2(n_268), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_117), .A2(n_515), .B1(n_517), .B2(n_518), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_117), .A2(n_118), .B1(n_541), .B2(n_542), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_117), .A2(n_567), .B(n_568), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_117), .A2(n_123), .B1(n_580), .B2(n_582), .Y(n_579) );
INVx6_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_118), .A2(n_202), .B(n_203), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_118), .B(n_217), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_118), .A2(n_211), .B(n_217), .C(n_221), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_118), .A2(n_529), .B(n_530), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_118), .A2(n_163), .B1(n_576), .B2(n_577), .Y(n_575) );
BUFx8_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g125 ( .A(n_119), .Y(n_125) );
INVx1_ASAP7_75t_L g149 ( .A(n_119), .Y(n_149) );
INVx1_ASAP7_75t_L g164 ( .A(n_119), .Y(n_164) );
INVx4_ASAP7_75t_L g196 ( .A(n_121), .Y(n_196) );
INVx2_ASAP7_75t_L g145 ( .A(n_122), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_122), .B(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g532 ( .A(n_122), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_123), .A2(n_181), .B(n_182), .Y(n_180) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_123), .A2(n_212), .B(n_215), .Y(n_211) );
AOI21x1_ASAP7_75t_L g563 ( .A1(n_123), .A2(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g200 ( .A(n_125), .Y(n_200) );
AOI31xp67_ASAP7_75t_L g539 ( .A1(n_126), .A2(n_131), .A3(n_540), .B(n_543), .Y(n_539) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2x1_ASAP7_75t_L g205 ( .A(n_127), .B(n_206), .Y(n_205) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g183 ( .A(n_128), .B(n_131), .Y(n_183) );
BUFx3_ASAP7_75t_L g513 ( .A(n_128), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_128), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g547 ( .A(n_128), .Y(n_547) );
INVx2_ASAP7_75t_SL g561 ( .A(n_128), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_128), .B(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g137 ( .A(n_129), .Y(n_137) );
INVx1_ASAP7_75t_L g206 ( .A(n_131), .Y(n_206) );
OAI21x1_ASAP7_75t_L g527 ( .A1(n_131), .A2(n_528), .B(n_531), .Y(n_527) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_131), .A2(n_549), .B(n_552), .Y(n_548) );
BUFx10_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
INVx1_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
BUFx10_ASAP7_75t_L g236 ( .A(n_132), .Y(n_236) );
AO31x2_ASAP7_75t_L g578 ( .A1(n_132), .A2(n_513), .A3(n_579), .B(n_583), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
BUFx2_ASAP7_75t_L g139 ( .A(n_136), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_136), .B(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g238 ( .A(n_136), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_136), .B(n_271), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_136), .B(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI21xp33_ASAP7_75t_L g221 ( .A1(n_137), .A2(n_168), .B(n_215), .Y(n_221) );
INVx2_ASAP7_75t_L g225 ( .A(n_137), .Y(n_225) );
INVx2_ASAP7_75t_L g269 ( .A(n_137), .Y(n_269) );
AND2x2_ASAP7_75t_L g246 ( .A(n_138), .B(n_170), .Y(n_246) );
INVx1_ASAP7_75t_L g253 ( .A(n_138), .Y(n_253) );
INVx1_ASAP7_75t_L g258 ( .A(n_138), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_138), .B(n_251), .Y(n_321) );
INVx1_ASAP7_75t_L g342 ( .A(n_138), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_138), .B(n_244), .Y(n_412) );
AO31x2_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .A3(n_150), .B(n_152), .Y(n_138) );
AOI21x1_ASAP7_75t_L g156 ( .A1(n_139), .A2(n_157), .B(n_169), .Y(n_156) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OAI22xp33_ASAP7_75t_L g231 ( .A1(n_143), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_231) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_146), .A2(n_163), .B(n_550), .C(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g161 ( .A(n_147), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_148), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_SL g517 ( .A(n_149), .Y(n_517) );
INVx1_ASAP7_75t_L g603 ( .A(n_149), .Y(n_603) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_150), .A2(n_513), .A3(n_514), .B(n_519), .Y(n_512) );
INVx2_ASAP7_75t_SL g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_SL g570 ( .A(n_151), .Y(n_570) );
INVx1_ASAP7_75t_L g305 ( .A(n_154), .Y(n_305) );
OR2x2_ASAP7_75t_L g357 ( .A(n_154), .B(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_170), .Y(n_154) );
AND2x2_ASAP7_75t_L g190 ( .A(n_155), .B(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_L g249 ( .A(n_155), .B(n_250), .Y(n_249) );
INVxp67_ASAP7_75t_L g255 ( .A(n_155), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_155), .B(n_187), .Y(n_333) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_165), .B(n_168), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_163), .Y(n_158) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_164), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g534 ( .A(n_164), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_168), .A2(n_599), .B(n_604), .Y(n_598) );
INVx3_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
INVx1_ASAP7_75t_L g299 ( .A(n_170), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_170), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g319 ( .A(n_170), .B(n_320), .Y(n_319) );
OR2x2_ASAP7_75t_L g341 ( .A(n_170), .B(n_342), .Y(n_341) );
NAND2x1p5_ASAP7_75t_SL g352 ( .A(n_170), .B(n_328), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_170), .B(n_258), .Y(n_442) );
AND2x4_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_180), .B(n_183), .Y(n_172) );
OAI21xp33_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B(n_177), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_176), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_190), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g380 ( .A1(n_185), .A2(n_381), .B1(n_382), .B2(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_188), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_186), .B(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_186), .B(n_437), .Y(n_436) );
OR2x2_ASAP7_75t_L g459 ( .A(n_186), .B(n_317), .Y(n_459) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
AND2x4_ASAP7_75t_L g257 ( .A(n_187), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_187), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g347 ( .A(n_187), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_L g298 ( .A(n_188), .B(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g388 ( .A(n_189), .Y(n_388) );
OR2x2_ASAP7_75t_L g462 ( .A(n_189), .B(n_389), .Y(n_462) );
INVx1_ASAP7_75t_L g293 ( .A(n_190), .Y(n_293) );
INVx3_ASAP7_75t_L g297 ( .A(n_191), .Y(n_297) );
BUFx2_ASAP7_75t_L g308 ( .A(n_191), .Y(n_308) );
BUFx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g278 ( .A(n_192), .B(n_222), .Y(n_278) );
INVx2_ASAP7_75t_L g324 ( .A(n_192), .Y(n_324) );
INVx1_ASAP7_75t_L g356 ( .A(n_192), .Y(n_356) );
AND2x2_ASAP7_75t_L g369 ( .A(n_192), .B(n_265), .Y(n_369) );
AND2x2_ASAP7_75t_L g391 ( .A(n_192), .B(n_290), .Y(n_391) );
NAND2x1p5_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
OAI21x1_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_201), .B(n_205), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_198), .C(n_199), .Y(n_195) );
INVx2_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_200), .A2(n_553), .B1(n_554), .B2(n_555), .Y(n_552) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g382 ( .A(n_208), .B(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_208), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g407 ( .A(n_208), .B(n_275), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_208), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g208 ( .A(n_209), .B(n_222), .Y(n_208) );
INVx2_ASAP7_75t_L g263 ( .A(n_209), .Y(n_263) );
AND2x2_ASAP7_75t_L g291 ( .A(n_209), .B(n_292), .Y(n_291) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_216), .B(n_220), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_214), .B(n_229), .Y(n_228) );
INVxp67_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
INVx3_ASAP7_75t_L g569 ( .A(n_219), .Y(n_569) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g264 ( .A(n_222), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g284 ( .A(n_222), .Y(n_284) );
INVx2_ASAP7_75t_L g292 ( .A(n_222), .Y(n_292) );
OR2x2_ASAP7_75t_L g312 ( .A(n_222), .B(n_265), .Y(n_312) );
AND2x2_ASAP7_75t_L g323 ( .A(n_222), .B(n_324), .Y(n_323) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_226), .B(n_237), .Y(n_222) );
AOI21x1_ASAP7_75t_L g597 ( .A1(n_223), .A2(n_598), .B(n_607), .Y(n_597) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_235), .Y(n_226) );
INVx1_ASAP7_75t_L g554 ( .A(n_233), .Y(n_554) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
AO31x2_ASAP7_75t_L g265 ( .A1(n_236), .A2(n_266), .A3(n_269), .B(n_270), .Y(n_265) );
OAI221xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .B1(n_247), .B2(n_252), .C(n_254), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
OAI32xp33_ASAP7_75t_L g353 ( .A1(n_242), .A2(n_256), .A3(n_354), .B1(n_357), .B2(n_358), .Y(n_353) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g343 ( .A(n_243), .Y(n_343) );
AND2x2_ASAP7_75t_L g379 ( .A(n_243), .B(n_257), .Y(n_379) );
INVx1_ASAP7_75t_L g443 ( .A(n_243), .Y(n_443) );
OR2x2_ASAP7_75t_L g317 ( .A(n_244), .B(n_251), .Y(n_317) );
INVx2_ASAP7_75t_L g328 ( .A(n_244), .Y(n_328) );
BUFx2_ASAP7_75t_SL g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g467 ( .A(n_246), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVxp67_ASAP7_75t_L g454 ( .A(n_249), .Y(n_454) );
INVx1_ASAP7_75t_L g468 ( .A(n_249), .Y(n_468) );
OR2x2_ASAP7_75t_L g348 ( .A(n_250), .B(n_328), .Y(n_348) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_252), .B(n_348), .Y(n_370) );
INVx1_ASAP7_75t_L g401 ( .A(n_252), .Y(n_401) );
BUFx3_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g435 ( .A(n_253), .Y(n_435) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2x1_ASAP7_75t_L g404 ( .A(n_255), .B(n_405), .Y(n_404) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_256), .A2(n_427), .B(n_432), .Y(n_426) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx2_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_264), .Y(n_260) );
AND2x2_ASAP7_75t_L g336 ( .A(n_261), .B(n_278), .Y(n_336) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_261), .Y(n_466) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g368 ( .A(n_262), .Y(n_368) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g350 ( .A(n_263), .B(n_324), .Y(n_350) );
AND2x2_ASAP7_75t_L g421 ( .A(n_263), .B(n_292), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_264), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g349 ( .A(n_264), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g428 ( .A(n_264), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g277 ( .A(n_265), .Y(n_277) );
INVx2_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_265), .B(n_281), .Y(n_338) );
AND2x2_ASAP7_75t_L g398 ( .A(n_265), .B(n_292), .Y(n_398) );
INVx2_ASAP7_75t_L g526 ( .A(n_269), .Y(n_526) );
NAND2xp33_ASAP7_75t_SL g272 ( .A(n_273), .B(n_279), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_278), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g373 ( .A(n_276), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_276), .B(n_356), .Y(n_448) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g280 ( .A(n_277), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g409 ( .A(n_277), .B(n_324), .Y(n_409) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
OR2x2_ASAP7_75t_L g354 ( .A(n_280), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g311 ( .A(n_281), .Y(n_311) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g337 ( .A(n_284), .B(n_338), .Y(n_337) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_298), .B1(n_300), .B2(n_301), .Y(n_285) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_293), .B(n_294), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_288), .B(n_297), .Y(n_300) );
BUFx2_ASAP7_75t_L g318 ( .A(n_288), .Y(n_318) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_291), .Y(n_288) );
INVx1_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g344 ( .A(n_291), .B(n_308), .Y(n_344) );
INVx2_ASAP7_75t_L g360 ( .A(n_291), .Y(n_360) );
AND2x2_ASAP7_75t_L g402 ( .A(n_291), .B(n_324), .Y(n_402) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g377 ( .A(n_297), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g424 ( .A(n_298), .B(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g455 ( .A(n_299), .Y(n_455) );
INVx2_ASAP7_75t_L g394 ( .A(n_302), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g303 ( .A(n_304), .B(n_313), .C(n_330), .D(n_345), .Y(n_303) );
NAND2xp33_ASAP7_75t_SL g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_306), .A2(n_384), .B1(n_400), .B2(n_402), .C(n_403), .Y(n_399) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NAND2x1_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g381 ( .A(n_310), .Y(n_381) );
OR2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
INVx2_ASAP7_75t_L g446 ( .A(n_312), .Y(n_446) );
AOI222xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_318), .B1(n_319), .B2(n_322), .C1(n_325), .C2(n_329), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g400 ( .A(n_316), .B(n_401), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_316), .A2(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g439 ( .A(n_317), .B(n_383), .Y(n_439) );
OAI21xp33_ASAP7_75t_SL g413 ( .A1(n_318), .A2(n_339), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_SL g384 ( .A(n_321), .Y(n_384) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g389 ( .A(n_328), .Y(n_389) );
AOI22xp33_ASAP7_75t_SL g330 ( .A1(n_331), .A2(n_334), .B1(n_339), .B2(n_344), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_336), .A2(n_346), .B1(n_349), .B2(n_351), .C(n_353), .Y(n_345) );
INVx3_ASAP7_75t_R g460 ( .A(n_337), .Y(n_460) );
INVx1_ASAP7_75t_L g378 ( .A(n_338), .Y(n_378) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_341), .Y(n_395) );
INVx1_ASAP7_75t_L g405 ( .A(n_341), .Y(n_405) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_350), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g423 ( .A(n_350), .Y(n_423) );
AND2x2_ASAP7_75t_L g451 ( .A(n_350), .B(n_398), .Y(n_451) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g445 ( .A(n_355), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_417), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_399), .C(n_413), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g363 ( .A(n_364), .B(n_375), .C(n_385), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OAI21xp33_ASAP7_75t_L g376 ( .A1(n_366), .A2(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx1_ASAP7_75t_L g416 ( .A(n_368), .Y(n_416) );
AND2x2_ASAP7_75t_L g457 ( .A(n_368), .B(n_446), .Y(n_457) );
NAND2x1_ASAP7_75t_L g415 ( .A(n_369), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx1_ASAP7_75t_L g437 ( .A(n_374), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_376), .B(n_380), .Y(n_375) );
INVx1_ASAP7_75t_L g429 ( .A(n_383), .Y(n_429) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_390), .B1(n_392), .B2(n_396), .Y(n_385) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g425 ( .A(n_389), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_391), .B(n_421), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_395), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g464 ( .A(n_397), .Y(n_464) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
OAI22xp33_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_406), .B1(n_408), .B2(n_410), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_418), .B(n_444), .Y(n_417) );
O2A1O1Ixp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_422), .B(n_424), .C(n_426), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp33_ASAP7_75t_L g433 ( .A1(n_420), .A2(n_434), .B(n_436), .Y(n_433) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
O2A1O1Ixp5_ASAP7_75t_SL g444 ( .A1(n_424), .A2(n_445), .B(n_447), .C(n_449), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_428), .A2(n_433), .B1(n_438), .B2(n_440), .Y(n_432) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI211xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B(n_456), .C(n_463), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_460), .B2(n_461), .Y(n_456) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI21xp5_ASAP7_75t_SL g463 ( .A1(n_464), .A2(n_465), .B(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
CKINVDCx8_ASAP7_75t_R g480 ( .A(n_470), .Y(n_480) );
INVx5_ASAP7_75t_L g854 ( .A(n_470), .Y(n_854) );
INVx3_ASAP7_75t_L g861 ( .A(n_470), .Y(n_861) );
AND2x6_ASAP7_75t_SL g470 ( .A(n_471), .B(n_474), .Y(n_470) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_474), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NOR2x1_ASAP7_75t_L g846 ( .A(n_475), .B(n_500), .Y(n_846) );
NOR2x1_ASAP7_75t_R g476 ( .A(n_477), .B(n_478), .Y(n_476) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
CKINVDCx11_ASAP7_75t_R g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g868 ( .A(n_485), .B(n_858), .Y(n_868) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g497 ( .A(n_486), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g843 ( .A(n_486), .B(n_844), .Y(n_843) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_486), .B(n_861), .Y(n_860) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B1(n_501), .B2(n_835), .C(n_838), .Y(n_487) );
NOR2xp67_ASAP7_75t_SL g490 ( .A(n_491), .B(n_495), .Y(n_490) );
INVx4_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g845 ( .A(n_493), .B(n_846), .Y(n_845) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
BUFx2_ASAP7_75t_L g837 ( .A(n_494), .Y(n_837) );
NOR2x1_ASAP7_75t_R g835 ( .A(n_495), .B(n_836), .Y(n_835) );
INVx5_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_SL g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_723), .Y(n_504) );
NAND4xp25_ASAP7_75t_L g505 ( .A(n_506), .B(n_655), .C(n_682), .D(n_713), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_507), .B(n_621), .Y(n_506) );
OAI21xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_557), .B(n_585), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g743 ( .A(n_510), .B(n_632), .Y(n_743) );
AND2x2_ASAP7_75t_L g750 ( .A(n_510), .B(n_751), .Y(n_750) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
OR2x2_ASAP7_75t_L g659 ( .A(n_511), .B(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_538), .Y(n_592) );
AND2x2_ASAP7_75t_L g616 ( .A(n_512), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g625 ( .A(n_512), .Y(n_625) );
OR2x2_ASAP7_75t_L g633 ( .A(n_512), .B(n_589), .Y(n_633) );
OR2x2_ASAP7_75t_L g654 ( .A(n_512), .B(n_617), .Y(n_654) );
AND2x2_ASAP7_75t_L g663 ( .A(n_512), .B(n_546), .Y(n_663) );
INVx1_ASAP7_75t_L g736 ( .A(n_512), .Y(n_736) );
AND2x2_ASAP7_75t_L g739 ( .A(n_512), .B(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_537), .Y(n_521) );
INVx2_ASAP7_75t_L g652 ( .A(n_522), .Y(n_652) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g760 ( .A(n_523), .Y(n_760) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g705 ( .A(n_524), .Y(n_705) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
OR2x2_ASAP7_75t_L g632 ( .A(n_525), .B(n_618), .Y(n_632) );
OAI21x1_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_536), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_526), .A2(n_527), .B(n_536), .Y(n_590) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .B(n_535), .Y(n_531) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_537), .Y(n_814) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_546), .Y(n_537) );
INVx2_ASAP7_75t_L g626 ( .A(n_538), .Y(n_626) );
AND2x2_ASAP7_75t_L g664 ( .A(n_538), .B(n_590), .Y(n_664) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g618 ( .A(n_539), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g620 ( .A(n_546), .B(n_590), .Y(n_620) );
INVx1_ASAP7_75t_L g706 ( .A(n_546), .Y(n_706) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_556), .Y(n_546) );
OA21x2_ASAP7_75t_L g589 ( .A1(n_547), .A2(n_548), .B(n_556), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_SL g764 ( .A1(n_557), .A2(n_765), .B(n_766), .C(n_768), .Y(n_764) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_572), .Y(n_557) );
OR2x2_ASAP7_75t_L g712 ( .A(n_558), .B(n_696), .Y(n_712) );
INVxp67_ASAP7_75t_SL g774 ( .A(n_558), .Y(n_774) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g608 ( .A(n_559), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g640 ( .A(n_559), .B(n_612), .Y(n_640) );
INVx3_ASAP7_75t_L g642 ( .A(n_559), .Y(n_642) );
INVxp67_ASAP7_75t_L g650 ( .A(n_559), .Y(n_650) );
INVx1_ASAP7_75t_L g660 ( .A(n_559), .Y(n_660) );
BUFx2_ASAP7_75t_L g686 ( .A(n_559), .Y(n_686) );
OR2x2_ASAP7_75t_L g709 ( .A(n_559), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g748 ( .A(n_559), .B(n_710), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_559), .B(n_578), .Y(n_796) );
INVx1_ASAP7_75t_L g822 ( .A(n_559), .Y(n_822) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OAI21x1_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_562), .B(n_571), .Y(n_560) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_566), .B(n_570), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g801 ( .A(n_572), .B(n_640), .Y(n_801) );
INVx2_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g641 ( .A(n_573), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g727 ( .A(n_573), .B(n_674), .Y(n_727) );
AND2x2_ASAP7_75t_L g744 ( .A(n_573), .B(n_673), .Y(n_744) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_578), .Y(n_573) );
OR2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_578), .Y(n_696) );
INVx1_ASAP7_75t_L g763 ( .A(n_574), .Y(n_763) );
INVx1_ASAP7_75t_L g776 ( .A(n_574), .Y(n_776) );
INVx3_ASAP7_75t_L g611 ( .A(n_578), .Y(n_611) );
AND2x2_ASAP7_75t_L g666 ( .A(n_578), .B(n_596), .Y(n_666) );
AND2x2_ASAP7_75t_L g687 ( .A(n_578), .B(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_593), .B1(n_610), .B2(n_613), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_586), .A2(n_721), .B1(n_824), .B2(n_826), .Y(n_823) );
INVx3_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OR2x2_ASAP7_75t_L g735 ( .A(n_588), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g769 ( .A(n_588), .Y(n_769) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
BUFx2_ASAP7_75t_L g645 ( .A(n_589), .Y(n_645) );
INVx2_ASAP7_75t_SL g669 ( .A(n_589), .Y(n_669) );
AND2x2_ASAP7_75t_L g689 ( .A(n_589), .B(n_625), .Y(n_689) );
INVx1_ASAP7_75t_L g740 ( .A(n_589), .Y(n_740) );
INVx1_ASAP7_75t_L g729 ( .A(n_591), .Y(n_729) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
AND2x4_ASAP7_75t_L g721 ( .A(n_592), .B(n_703), .Y(n_721) );
AO22x1_ASAP7_75t_L g809 ( .A1(n_593), .A2(n_662), .B1(n_810), .B2(n_811), .Y(n_809) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_608), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g628 ( .A(n_596), .Y(n_628) );
INVx1_ASAP7_75t_L g637 ( .A(n_596), .Y(n_637) );
INVx1_ASAP7_75t_L g688 ( .A(n_596), .Y(n_688) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g612 ( .A(n_597), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g599 ( .A(n_600), .B(n_603), .Y(n_599) );
AND2x2_ASAP7_75t_L g808 ( .A(n_608), .B(n_718), .Y(n_808) );
AND2x4_ASAP7_75t_L g675 ( .A(n_609), .B(n_611), .Y(n_675) );
INVx1_ASAP7_75t_L g710 ( .A(n_609), .Y(n_710) );
INVx1_ASAP7_75t_L g784 ( .A(n_609), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_610), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_610), .B(n_828), .Y(n_827) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
AND2x4_ASAP7_75t_L g636 ( .A(n_611), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g755 ( .A(n_611), .Y(n_755) );
INVx1_ASAP7_75t_L g674 ( .A(n_612), .Y(n_674) );
INVx1_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
OR2x2_ASAP7_75t_L g775 ( .A(n_612), .B(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g802 ( .A(n_616), .B(n_645), .Y(n_802) );
AND2x2_ASAP7_75t_L g810 ( .A(n_616), .B(n_652), .Y(n_810) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g752 ( .A(n_619), .B(n_702), .Y(n_752) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g623 ( .A(n_620), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g730 ( .A(n_620), .Y(n_730) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_627), .B(n_629), .C(n_647), .Y(n_621) );
OAI322xp33_ASAP7_75t_L g667 ( .A1(n_622), .A2(n_659), .A3(n_668), .B1(n_671), .B2(n_676), .C1(n_679), .C2(n_681), .Y(n_667) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g677 ( .A(n_624), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g733 ( .A(n_624), .Y(n_733) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx1_ASAP7_75t_L g702 ( .A(n_626), .Y(n_702) );
AND2x2_ASAP7_75t_L g741 ( .A(n_626), .B(n_705), .Y(n_741) );
INVx1_ASAP7_75t_L g834 ( .A(n_626), .Y(n_834) );
INVx1_ASAP7_75t_L g812 ( .A(n_627), .Y(n_812) );
OAI211xp5_ASAP7_75t_L g832 ( .A1(n_627), .A2(n_711), .B(n_754), .C(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_634), .B1(n_641), .B2(n_643), .Y(n_629) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_630), .A2(n_708), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g646 ( .A(n_632), .Y(n_646) );
INVx1_ASAP7_75t_L g670 ( .A(n_632), .Y(n_670) );
INVx1_ASAP7_75t_L g751 ( .A(n_632), .Y(n_751) );
INVx1_ASAP7_75t_L g780 ( .A(n_633), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_638), .Y(n_634) );
HB1xp67_ASAP7_75t_L g831 ( .A(n_635), .Y(n_831) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NAND2x1p5_ASAP7_75t_L g767 ( .A(n_636), .B(n_748), .Y(n_767) );
INVx1_ASAP7_75t_L g718 ( .A(n_637), .Y(n_718) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2x1_ASAP7_75t_SL g679 ( .A(n_639), .B(n_680), .Y(n_679) );
INVx3_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_640), .B(n_675), .Y(n_699) );
AND2x2_ASAP7_75t_L g762 ( .A(n_642), .B(n_763), .Y(n_762) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g661 ( .A(n_645), .B(n_646), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_651), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g815 ( .A(n_650), .B(n_672), .Y(n_815) );
INVx1_ASAP7_75t_L g828 ( .A(n_650), .Y(n_828) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g732 ( .A(n_652), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_653), .B(n_678), .Y(n_722) );
INVx1_ASAP7_75t_L g765 ( .A(n_653), .Y(n_765) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g692 ( .A(n_654), .Y(n_692) );
OR2x2_ASAP7_75t_L g821 ( .A(n_654), .B(n_822), .Y(n_821) );
O2A1O1Ixp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_662), .B(n_665), .C(n_667), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_658), .B(n_661), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g754 ( .A(n_660), .B(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g799 ( .A(n_661), .Y(n_799) );
INVx2_ASAP7_75t_L g792 ( .A(n_662), .Y(n_792) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_663), .A2(n_714), .B(n_719), .Y(n_713) );
AND2x2_ASAP7_75t_L g779 ( .A(n_664), .B(n_780), .Y(n_779) );
BUFx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g747 ( .A(n_666), .B(n_748), .Y(n_747) );
AND2x4_ASAP7_75t_L g761 ( .A(n_666), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_666), .B(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx2_ASAP7_75t_L g678 ( .A(n_669), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_669), .B(n_692), .Y(n_691) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_669), .Y(n_817) );
AOI21xp33_ASAP7_75t_L g719 ( .A1(n_671), .A2(n_720), .B(n_722), .Y(n_719) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx3_ASAP7_75t_L g681 ( .A(n_675), .Y(n_681) );
AND2x4_ASAP7_75t_L g806 ( .A(n_675), .B(n_694), .Y(n_806) );
INVx2_ASAP7_75t_SL g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_689), .B1(n_690), .B2(n_693), .C(n_697), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g803 ( .A(n_685), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
BUFx2_ASAP7_75t_L g716 ( .A(n_686), .Y(n_716) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
OR2x2_ASAP7_75t_L g825 ( .A(n_694), .B(n_709), .Y(n_825) );
AND2x4_ASAP7_75t_L g717 ( .A(n_695), .B(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI21xp5_ASAP7_75t_SL g697 ( .A1(n_698), .A2(n_700), .B(n_707), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
AND2x2_ASAP7_75t_L g786 ( .A(n_703), .B(n_736), .Y(n_786) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g798 ( .A(n_717), .Y(n_798) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g807 ( .A(n_721), .B(n_808), .Y(n_807) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_724), .B(n_770), .C(n_813), .Y(n_723) );
NOR3xp33_ASAP7_75t_L g724 ( .A(n_725), .B(n_745), .C(n_764), .Y(n_724) );
OAI21xp5_ASAP7_75t_SL g725 ( .A1(n_726), .A2(n_728), .B(n_737), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI211x1_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B(n_731), .C(n_734), .Y(n_728) );
OAI322xp33_ASAP7_75t_L g771 ( .A1(n_729), .A2(n_772), .A3(n_777), .B1(n_778), .B2(n_781), .C1(n_785), .C2(n_787), .Y(n_771) );
NOR2xp67_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
O2A1O1Ixp5_ASAP7_75t_SL g829 ( .A1(n_732), .A2(n_830), .B(n_831), .C(n_832), .Y(n_829) );
INVx3_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_736), .B(n_760), .Y(n_759) );
OAI21xp5_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_742), .B(n_744), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_738), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
AND2x4_ASAP7_75t_L g738 ( .A(n_739), .B(n_741), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_749), .B1(n_752), .B2(n_753), .C(n_756), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_761), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
HB1xp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g790 ( .A(n_763), .Y(n_790) );
INVx1_ASAP7_75t_L g797 ( .A(n_763), .Y(n_797) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g777 ( .A(n_769), .Y(n_777) );
NOR4xp25_ASAP7_75t_L g770 ( .A(n_771), .B(n_791), .C(n_804), .D(n_809), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR2x1p5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx2_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g811 ( .A(n_790), .B(n_812), .Y(n_811) );
OAI221xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_798), .B2(n_799), .C(n_800), .Y(n_791) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_792), .A2(n_805), .B(n_807), .Y(n_804) );
INVxp67_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
OR2x2_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g820 ( .A(n_812), .Y(n_820) );
AOI211xp5_ASAP7_75t_L g813 ( .A1(n_814), .A2(n_815), .B(n_816), .C(n_829), .Y(n_813) );
OAI21xp5_ASAP7_75t_SL g816 ( .A1(n_817), .A2(n_818), .B(n_823), .Y(n_816) );
INVx1_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NOR2x1_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
HB1xp67_ASAP7_75t_L g830 ( .A(n_821), .Y(n_830) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .Y(n_838) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx10_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_850), .Y(n_849) );
CKINVDCx16_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_854), .Y(n_851) );
INVx2_ASAP7_75t_SL g859 ( .A(n_852), .Y(n_859) );
INVx4_ASAP7_75t_SL g856 ( .A(n_857), .Y(n_856) );
OR2x4_ASAP7_75t_L g857 ( .A(n_858), .B(n_860), .Y(n_857) );
BUFx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OR2x6_ASAP7_75t_L g866 ( .A(n_861), .B(n_867), .Y(n_866) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
CKINVDCx20_ASAP7_75t_R g863 ( .A(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g864 ( .A(n_865), .Y(n_864) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
endmodule