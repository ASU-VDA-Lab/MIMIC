module fake_jpeg_17583_n_190 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_5),
.B(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_5),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_34),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_20),
.Y(n_75)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_32),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_37),
.B1(n_26),
.B2(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_21),
.B(n_7),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_45),
.B(n_28),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_57),
.B(n_60),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_32),
.B1(n_31),
.B2(n_37),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_58),
.A2(n_68),
.B1(n_71),
.B2(n_74),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_52),
.B(n_28),
.Y(n_60)
);

NAND3xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_22),
.C(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_74),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_86),
.B(n_11),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_33),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_67),
.B1(n_12),
.B2(n_10),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_33),
.B1(n_23),
.B2(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_16),
.C(n_23),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_81),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_23),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_42),
.A2(n_23),
.B1(n_21),
.B2(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_39),
.B(n_20),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_38),
.B(n_17),
.C(n_35),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_17),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_17),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_50),
.A2(n_17),
.B1(n_19),
.B2(n_10),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_19),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_88),
.B(n_92),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_96),
.Y(n_118)
);

INVx5_ASAP7_75t_SL g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_60),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_9),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_112),
.B1(n_83),
.B2(n_85),
.Y(n_121)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_57),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_81),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_111),
.Y(n_128)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_109),
.A2(n_80),
.B1(n_83),
.B2(n_107),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_66),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_76),
.A2(n_77),
.B1(n_63),
.B2(n_78),
.Y(n_112)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_111),
.A2(n_72),
.B1(n_77),
.B2(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_115),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_102),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_91),
.B(n_93),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_109),
.B1(n_105),
.B2(n_95),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_87),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_122),
.A2(n_127),
.B(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_129),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_125),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_80),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_106),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_90),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_114),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_137),
.Y(n_148)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_108),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_122),
.B1(n_127),
.B2(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_136),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_97),
.C(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_145),
.Y(n_155)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_117),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_145),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_149),
.B(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_143),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_128),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_153),
.A2(n_160),
.B1(n_135),
.B2(n_133),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_159),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_144),
.A2(n_118),
.B(n_115),
.C(n_119),
.D(n_113),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_113),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_166),
.B(n_169),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_140),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_168),
.B(n_171),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_150),
.A2(n_147),
.B1(n_137),
.B2(n_142),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_149),
.B(n_132),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_147),
.B1(n_131),
.B2(n_146),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_173),
.A2(n_165),
.B1(n_157),
.B2(n_167),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_166),
.A2(n_160),
.B(n_153),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_178),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_177),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_160),
.B(n_153),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_179),
.B(n_182),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_177),
.B1(n_134),
.B2(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_164),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_172),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_184),
.B1(n_183),
.B2(n_180),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_186),
.Y(n_190)
);


endmodule