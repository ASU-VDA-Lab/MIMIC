module fake_jpeg_31695_n_350 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_18),
.B(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_19),
.B(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_48),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_32),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

HAxp5_ASAP7_75t_SL g53 ( 
.A(n_20),
.B(n_30),
.CON(n_53),
.SN(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_53),
.A2(n_28),
.B(n_3),
.C(n_4),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_55),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_29),
.B(n_9),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_58),
.B(n_61),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_30),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_30),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_40),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_37),
.B1(n_33),
.B2(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_68),
.A2(n_78),
.B1(n_87),
.B2(n_88),
.Y(n_121)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_71),
.Y(n_131)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_41),
.B1(n_22),
.B2(n_39),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_73),
.A2(n_74),
.B1(n_83),
.B2(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_22),
.B1(n_39),
.B2(n_37),
.Y(n_74)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_1),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_63),
.A2(n_37),
.B1(n_33),
.B2(n_39),
.Y(n_78)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_33),
.Y(n_80)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_80),
.A2(n_91),
.B1(n_106),
.B2(n_111),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_39),
.C(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_82),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_40),
.B1(n_35),
.B2(n_32),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_26),
.B1(n_21),
.B2(n_23),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_64),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_25),
.B(n_36),
.Y(n_90)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_90),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_28),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_60),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_96),
.Y(n_150)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_60),
.A2(n_38),
.B1(n_34),
.B2(n_27),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_99),
.A2(n_110),
.B1(n_50),
.B2(n_28),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_65),
.A2(n_17),
.B1(n_27),
.B2(n_11),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_50),
.B1(n_67),
.B2(n_28),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_49),
.B(n_1),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_114),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_46),
.A2(n_17),
.B1(n_11),
.B2(n_16),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_46),
.B(n_56),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_100),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_116),
.B(n_135),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_120),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_56),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_137),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_80),
.B1(n_106),
.B2(n_114),
.Y(n_172)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_127),
.Y(n_180)
);

NOR2x1_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_128),
.B(n_14),
.Y(n_188)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_106),
.B1(n_80),
.B2(n_91),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_103),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_77),
.B(n_2),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_10),
.B1(n_14),
.B2(n_12),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_138),
.A2(n_100),
.B1(n_85),
.B2(n_91),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_109),
.B(n_4),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_80),
.Y(n_162)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

OR2x4_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_106),
.Y(n_170)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_107),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx6_ASAP7_75t_SL g148 ( 
.A(n_100),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_151),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_153),
.B(n_163),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_74),
.B1(n_73),
.B2(n_114),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_156),
.A2(n_104),
.B1(n_144),
.B2(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_115),
.Y(n_202)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_146),
.B(n_90),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_170),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_168),
.A2(n_188),
.B(n_121),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_81),
.C(n_109),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_143),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_91),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_181),
.B1(n_189),
.B2(n_128),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_119),
.B(n_76),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_117),
.B(n_112),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_186),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_84),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_182),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_146),
.A2(n_75),
.B1(n_98),
.B2(n_93),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_131),
.B(n_112),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_86),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_187),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_75),
.Y(n_186)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_132),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_146),
.A2(n_98),
.B1(n_93),
.B2(n_70),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_177),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_190),
.Y(n_230)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_203),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_193),
.B(n_199),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_194),
.A2(n_157),
.B(n_158),
.C(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_124),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_166),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_200),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_115),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_205),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_202),
.B(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_140),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_155),
.B(n_152),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_223),
.C(n_174),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_165),
.A2(n_148),
.B1(n_139),
.B2(n_122),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_207),
.A2(n_216),
.B(n_217),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_139),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_208),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_189),
.A2(n_145),
.B1(n_151),
.B2(n_141),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_209),
.A2(n_210),
.B(n_188),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_116),
.B(n_132),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_181),
.B1(n_172),
.B2(n_184),
.Y(n_225)
);

NAND5xp2_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_149),
.C(n_135),
.D(n_123),
.E(n_147),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_133),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_214),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_186),
.B(n_123),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_160),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_175),
.C(n_160),
.Y(n_235)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_183),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_219),
.A2(n_222),
.B1(n_178),
.B2(n_180),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_163),
.A2(n_130),
.B(n_127),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_239),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_225),
.A2(n_247),
.B1(n_193),
.B2(n_212),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_197),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_201),
.C(n_195),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_232),
.C(n_250),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_221),
.C(n_202),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_235),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_236),
.A2(n_238),
.B(n_242),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_170),
.B(n_162),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_203),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_158),
.B(n_154),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_245),
.A2(n_217),
.B(n_216),
.Y(n_269)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_180),
.B1(n_104),
.B2(n_157),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_192),
.A2(n_209),
.B1(n_206),
.B2(n_204),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_249),
.A2(n_251),
.B1(n_198),
.B2(n_191),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_213),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_213),
.A2(n_215),
.B1(n_212),
.B2(n_220),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_260),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_254),
.Y(n_279)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_258),
.A2(n_244),
.B1(n_248),
.B2(n_251),
.Y(n_281)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_194),
.C(n_190),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_259),
.B(n_226),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_230),
.B(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_261),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_200),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_264),
.B1(n_268),
.B2(n_270),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_218),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_272),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_225),
.B1(n_247),
.B2(n_244),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_227),
.B(n_229),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_238),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_240),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_269),
.A2(n_242),
.B(n_5),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_248),
.B(n_222),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_154),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_273),
.B1(n_266),
.B2(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_241),
.B(n_236),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_227),
.C(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_274),
.B(n_280),
.C(n_285),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_289),
.B1(n_292),
.B2(n_252),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_232),
.C(n_249),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_286),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_284),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

FAx1_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_244),
.CI(n_245),
.CON(n_286),
.SN(n_286)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_252),
.A2(n_242),
.B1(n_219),
.B2(n_178),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_242),
.C(n_129),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_257),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_262),
.B(n_269),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_258),
.A2(n_10),
.B1(n_11),
.B2(n_15),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_270),
.B1(n_278),
.B2(n_275),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_277),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_297),
.B(n_299),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_302),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_268),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_304),
.Y(n_319)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_253),
.C(n_273),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_305),
.B(n_292),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_265),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_259),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_291),
.A2(n_256),
.B(n_263),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_306),
.A2(n_289),
.B(n_286),
.Y(n_314)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_288),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_307),
.A2(n_288),
.B1(n_276),
.B2(n_261),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_308),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_309),
.B(n_318),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_280),
.C(n_290),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_312),
.C(n_317),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_287),
.C(n_281),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_313),
.A2(n_306),
.B(n_295),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_314),
.A2(n_300),
.B(n_6),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_305),
.B1(n_294),
.B2(n_308),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_286),
.C(n_255),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_4),
.C(n_6),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_296),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_325),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_328),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_311),
.B(n_303),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_312),
.Y(n_331)
);

INVx6_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_303),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_318),
.B(n_304),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_329),
.B(n_310),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_6),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_337),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_327),
.A2(n_319),
.B1(n_310),
.B2(n_7),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_319),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_335),
.B(n_338),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_333),
.A2(n_323),
.B(n_325),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_339),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_336),
.A2(n_323),
.B(n_330),
.Y(n_343)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_343),
.A2(n_334),
.A3(n_322),
.B1(n_331),
.B2(n_335),
.C1(n_326),
.C2(n_338),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_342),
.A2(n_7),
.B1(n_334),
.B2(n_340),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_347),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_348),
.A2(n_341),
.B(n_344),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_346),
.Y(n_350)
);


endmodule