module fake_jpeg_25855_n_99 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_99);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_30),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_11),
.B(n_0),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_24),
.B(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_14),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_46),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_43),
.B1(n_22),
.B2(n_14),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_28),
.B1(n_18),
.B2(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_25),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_47),
.B(n_51),
.Y(n_61)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_48),
.B(n_52),
.Y(n_55)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR3xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_53),
.C(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_64),
.B1(n_65),
.B2(n_20),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_26),
.C(n_23),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g72 ( 
.A(n_60),
.B(n_62),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_26),
.C(n_23),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_12),
.B(n_18),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_12),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_67),
.B(n_68),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_59),
.A2(n_26),
.B(n_40),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_2),
.B(n_3),
.Y(n_79)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_41),
.B1(n_50),
.B2(n_49),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_61),
.B1(n_22),
.B2(n_58),
.C(n_21),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_30),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_75),
.A2(n_23),
.B(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_79),
.B1(n_15),
.B2(n_3),
.Y(n_87)
);

AO221x1_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.C(n_62),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_13),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_72),
.C(n_75),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_79),
.C(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_72),
.B1(n_21),
.B2(n_15),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_81),
.B(n_5),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.Y(n_92)
);

XNOR2x1_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_21),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_93),
.B(n_4),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_83),
.B(n_7),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_95),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_92),
.C(n_96),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_4),
.Y(n_99)
);


endmodule