module real_jpeg_8469_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_206;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_0),
.A2(n_1),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_10),
.B1(n_23),
.B2(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_0),
.A2(n_25),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_1),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_20),
.Y(n_21)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_2),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_9),
.B(n_33),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_23),
.B(n_46),
.C(n_47),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_5),
.B(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_5),
.A2(n_6),
.B1(n_38),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_5),
.A2(n_6),
.A3(n_23),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_31),
.B(n_34),
.C(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_6),
.B(n_34),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_6),
.A2(n_8),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_10),
.B1(n_38),
.B2(n_50),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_9),
.B1(n_26),
.B2(n_38),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_6),
.A2(n_26),
.B(n_34),
.C(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

HAxp5_ASAP7_75t_SL g25 ( 
.A(n_7),
.B(n_26),
.CON(n_25),
.SN(n_25)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_9),
.A2(n_23),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_9),
.B(n_23),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_9),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_9),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_9),
.B(n_47),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_50),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_87),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_85),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_69),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_14),
.B(n_69),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_57),
.B1(n_58),
.B2(n_68),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_52),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_17),
.A2(n_59),
.B(n_65),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_17),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_17),
.B(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_17),
.A2(n_51),
.B1(n_59),
.B2(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_17),
.A2(n_51),
.B1(n_55),
.B2(n_78),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_17),
.A2(n_51),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_25),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_23),
.B(n_24),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_26),
.B(n_31),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_26),
.B(n_63),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_40),
.B2(n_41),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_35),
.B(n_37),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_31),
.A2(n_35),
.B1(n_37),
.B2(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_31),
.A2(n_35),
.B1(n_54),
.B2(n_67),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_31),
.A2(n_35),
.B(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_32),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_38),
.B(n_48),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B1(n_47),
.B2(n_49),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_44),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_47),
.Y(n_56)
);

AOI211xp5_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_75),
.B(n_80),
.C(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_52),
.A2(n_53),
.B(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_55),
.A2(n_75),
.B1(n_78),
.B2(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_55),
.B(n_109),
.C(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_55),
.A2(n_78),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_59),
.A2(n_66),
.B1(n_84),
.B2(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_63),
.B1(n_64),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_62),
.A2(n_63),
.B1(n_74),
.B2(n_100),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_62),
.A2(n_63),
.B(n_100),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_66),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_81),
.C(n_82),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_70),
.A2(n_71),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_SL g71 ( 
.A1(n_72),
.A2(n_76),
.B(n_79),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_72),
.A2(n_103),
.B1(n_104),
.B2(n_198),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_72),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_75),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_73),
.A2(n_75),
.B1(n_96),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_73),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_96),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_75),
.A2(n_96),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_75),
.A2(n_96),
.B1(n_131),
.B2(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_75),
.B(n_109),
.C(n_135),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_75),
.A2(n_96),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_75),
.B(n_163),
.C(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_75),
.B(n_99),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_76),
.A2(n_79),
.B(n_187),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_77),
.A2(n_80),
.B(n_110),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_96),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_78),
.A2(n_96),
.B(n_157),
.C(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_81),
.B(n_82),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_203),
.B(n_208),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_193),
.B(n_202),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_124),
.B(n_180),
.C(n_192),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_111),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_91),
.B(n_111),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_93),
.B(n_98),
.C(n_102),
.Y(n_181)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_103),
.A2(n_104),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_106),
.A2(n_109),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_109),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_118),
.B1(n_134),
.B2(n_137),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_109),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_118),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_153),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_120),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_112),
.A2(n_113),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_114),
.A2(n_115),
.B1(n_152),
.B2(n_157),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_146),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_120),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_179),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_172),
.B(n_178),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_159),
.B(n_171),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_149),
.B(n_158),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_138),
.B(n_148),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_134),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_145),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_152),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_174),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_181),
.B(n_182),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_184),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_190),
.C(n_191),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_187),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_194),
.B(n_195),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_201),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_199),
.C(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_204),
.B(n_205),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);


endmodule