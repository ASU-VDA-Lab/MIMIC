module real_aes_8114_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_434;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_404;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_279;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
AOI22xp33_ASAP7_75t_SL g855 ( .A1(n_0), .A2(n_185), .B1(n_373), .B2(n_704), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_1), .A2(n_257), .B1(n_387), .B2(n_845), .Y(n_844) );
CKINVDCx20_ASAP7_75t_R g826 ( .A(n_2), .Y(n_826) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_3), .A2(n_16), .B1(n_315), .B2(n_376), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g372 ( .A1(n_4), .A2(n_109), .B1(n_327), .B2(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g479 ( .A(n_5), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_6), .A2(n_18), .B1(n_547), .B2(n_560), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_7), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_8), .A2(n_124), .B1(n_362), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g476 ( .A(n_9), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_10), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_11), .A2(n_127), .B1(n_340), .B2(n_607), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_12), .A2(n_173), .B1(n_417), .B2(n_578), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_13), .A2(n_118), .B1(n_432), .B2(n_570), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_14), .A2(n_49), .B1(n_546), .B2(n_547), .Y(n_545) );
AOI222xp33_ASAP7_75t_L g731 ( .A1(n_15), .A2(n_121), .B1(n_219), .B2(n_327), .C1(n_414), .C2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_SL g815 ( .A1(n_17), .A2(n_55), .B1(n_575), .B2(n_816), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g460 ( .A(n_19), .Y(n_460) );
AOI222xp33_ASAP7_75t_L g579 ( .A1(n_20), .A2(n_85), .B1(n_139), .B2(n_376), .C1(n_524), .C2(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_21), .B(n_288), .Y(n_287) );
AOI22xp33_ASAP7_75t_SL g749 ( .A1(n_22), .A2(n_168), .B1(n_604), .B2(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_23), .Y(n_451) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_24), .Y(n_507) );
AO22x2_ASAP7_75t_L g296 ( .A1(n_25), .A2(n_86), .B1(n_292), .B2(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g799 ( .A(n_25), .Y(n_799) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_26), .A2(n_119), .B1(n_696), .B2(n_698), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_27), .A2(n_203), .B1(n_340), .B2(n_387), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_28), .A2(n_144), .B1(n_435), .B2(n_438), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_29), .A2(n_133), .B1(n_360), .B2(n_462), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_30), .B(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_31), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_32), .A2(n_269), .B1(n_345), .B2(n_348), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_33), .A2(n_157), .B1(n_483), .B2(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g520 ( .A(n_34), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_35), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_36), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_37), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_38), .B(n_303), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_39), .A2(n_198), .B1(n_330), .B2(n_578), .Y(n_814) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_40), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_41), .A2(n_803), .B1(n_804), .B2(n_832), .Y(n_802) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_41), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g710 ( .A(n_42), .Y(n_710) );
AO22x2_ASAP7_75t_L g291 ( .A1(n_43), .A2(n_89), .B1(n_292), .B2(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g800 ( .A(n_43), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g448 ( .A1(n_44), .A2(n_131), .B1(n_328), .B2(n_331), .Y(n_448) );
INVx1_ASAP7_75t_L g403 ( .A(n_45), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_46), .A2(n_143), .B1(n_685), .B2(n_686), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g746 ( .A1(n_47), .A2(n_179), .B1(n_316), .B2(n_330), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_48), .A2(n_259), .B1(n_378), .B2(n_379), .Y(n_377) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_50), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_51), .A2(n_84), .B1(n_546), .B2(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_52), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_53), .Y(n_701) );
AOI222xp33_ASAP7_75t_L g856 ( .A1(n_54), .A2(n_147), .B1(n_161), .B2(n_321), .C1(n_376), .C2(n_646), .Y(n_856) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_56), .A2(n_60), .B1(n_354), .B2(n_820), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_57), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_58), .A2(n_123), .B1(n_565), .B2(n_629), .Y(n_628) );
AOI222xp33_ASAP7_75t_L g672 ( .A1(n_59), .A2(n_194), .B1(n_255), .B2(n_309), .C1(n_594), .C2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_61), .A2(n_71), .B1(n_360), .B2(n_362), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_62), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_63), .Y(n_587) );
INVxp67_ASAP7_75t_L g840 ( .A(n_64), .Y(n_840) );
XNOR2x2_ASAP7_75t_L g841 ( .A(n_64), .B(n_842), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_65), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_66), .A2(n_263), .B1(n_440), .B2(n_486), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_67), .A2(n_151), .B1(n_315), .B2(n_417), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_68), .A2(n_187), .B1(n_345), .B2(n_670), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g748 ( .A1(n_69), .A2(n_208), .B1(n_345), .B2(n_440), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_70), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_72), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_73), .A2(n_199), .B1(n_704), .B2(n_706), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_74), .Y(n_591) );
AO22x2_ASAP7_75t_L g583 ( .A1(n_75), .A2(n_584), .B1(n_608), .B2(n_609), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_75), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_76), .A2(n_232), .B1(n_438), .B2(n_604), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_77), .A2(n_162), .B1(n_645), .B2(n_646), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_78), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_79), .A2(n_105), .B1(n_607), .B2(n_822), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_80), .A2(n_238), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_81), .A2(n_227), .B1(n_575), .B2(n_576), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_82), .A2(n_149), .B1(n_340), .B2(n_348), .Y(n_382) );
AOI22xp5_ASAP7_75t_SL g482 ( .A1(n_83), .A2(n_148), .B1(n_483), .B2(n_484), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_87), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_88), .A2(n_137), .B1(n_376), .B2(n_646), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_90), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_91), .A2(n_211), .B1(n_361), .B2(n_390), .Y(n_389) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_92), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_93), .Y(n_683) );
INVx1_ASAP7_75t_L g278 ( .A(n_94), .Y(n_278) );
AOI22xp5_ASAP7_75t_SL g513 ( .A1(n_95), .A2(n_514), .B1(n_552), .B2(n_553), .Y(n_513) );
INVx1_ASAP7_75t_L g553 ( .A(n_95), .Y(n_553) );
INVx1_ASAP7_75t_L g364 ( .A(n_96), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g383 ( .A1(n_97), .A2(n_209), .B1(n_345), .B2(n_384), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_98), .A2(n_134), .B1(n_570), .B2(n_572), .Y(n_569) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_99), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_100), .A2(n_190), .B1(n_416), .B2(n_417), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_101), .Y(n_631) );
INVx1_ASAP7_75t_L g276 ( .A(n_102), .Y(n_276) );
AOI22xp33_ASAP7_75t_SL g386 ( .A1(n_103), .A2(n_167), .B1(n_356), .B2(n_387), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_104), .A2(n_145), .B1(n_309), .B2(n_328), .Y(n_741) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_106), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_107), .A2(n_245), .B1(n_429), .B2(n_849), .Y(n_848) );
INVx1_ASAP7_75t_L g450 ( .A(n_108), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_110), .A2(n_156), .B1(n_330), .B2(n_667), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_111), .A2(n_244), .B1(n_607), .B2(n_726), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_112), .A2(n_221), .B1(n_309), .B2(n_315), .Y(n_308) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_113), .Y(n_760) );
AOI211xp5_ASAP7_75t_L g823 ( .A1(n_114), .A2(n_431), .B(n_824), .C(n_829), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_115), .A2(n_171), .B1(n_355), .B2(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_116), .B(n_303), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_117), .A2(n_180), .B1(n_337), .B2(n_340), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_120), .B(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g643 ( .A(n_122), .Y(n_643) );
INVx1_ASAP7_75t_L g325 ( .A(n_125), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_126), .B(n_379), .Y(n_648) );
INVx1_ASAP7_75t_L g477 ( .A(n_128), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_129), .A2(n_233), .B1(n_356), .B2(n_390), .Y(n_722) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_130), .Y(n_767) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_132), .A2(n_262), .B1(n_384), .B2(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_135), .A2(n_261), .B1(n_565), .B2(n_696), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_136), .A2(n_253), .B1(n_438), .B2(n_565), .Y(n_850) );
AOI22xp5_ASAP7_75t_SL g755 ( .A1(n_138), .A2(n_756), .B1(n_780), .B2(n_781), .Y(n_755) );
INVx1_ASAP7_75t_L g781 ( .A(n_138), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_140), .Y(n_633) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_141), .Y(n_733) );
INVx2_ASAP7_75t_L g279 ( .A(n_142), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_146), .A2(n_150), .B1(n_432), .B2(n_570), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_152), .Y(n_808) );
INVx1_ASAP7_75t_L g419 ( .A(n_153), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_154), .A2(n_230), .B1(n_331), .B2(n_578), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_155), .Y(n_759) );
AND2x6_ASAP7_75t_L g275 ( .A(n_158), .B(n_276), .Y(n_275) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_158), .Y(n_793) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_159), .A2(n_229), .B1(n_292), .B2(n_293), .Y(n_301) );
INVx1_ASAP7_75t_L g422 ( .A(n_160), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_163), .A2(n_251), .B1(n_384), .B2(n_486), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g810 ( .A(n_164), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_165), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_166), .A2(n_210), .B1(n_661), .B2(n_662), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_169), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_170), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_172), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_174), .A2(n_271), .B(n_280), .C(n_801), .Y(n_270) );
OA22x2_ASAP7_75t_L g397 ( .A1(n_175), .A2(n_398), .B1(n_399), .B2(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_175), .Y(n_398) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_176), .A2(n_267), .B1(n_440), .B2(n_441), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_177), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_178), .Y(n_728) );
AOI22xp33_ASAP7_75t_SL g353 ( .A1(n_181), .A2(n_204), .B1(n_354), .B2(n_356), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_182), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_183), .A2(n_191), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_184), .A2(n_676), .B1(n_714), .B2(n_715), .Y(n_675) );
INVx1_ASAP7_75t_L g714 ( .A(n_184), .Y(n_714) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_186), .A2(n_218), .B1(n_540), .B2(n_541), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_188), .A2(n_254), .B1(n_337), .B2(n_607), .Y(n_606) );
AOI22xp33_ASAP7_75t_SL g752 ( .A1(n_189), .A2(n_248), .B1(n_340), .B2(n_348), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_192), .A2(n_225), .B1(n_431), .B2(n_432), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_193), .A2(n_222), .B1(n_416), .B2(n_417), .Y(n_415) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_195), .A2(n_246), .B1(n_292), .B2(n_297), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_196), .A2(n_260), .B1(n_327), .B2(n_330), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_197), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_200), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_201), .A2(n_223), .B1(n_428), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_202), .A2(n_249), .B1(n_593), .B2(n_594), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_205), .Y(n_638) );
INVx1_ASAP7_75t_L g447 ( .A(n_206), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_207), .A2(n_215), .B1(n_563), .B2(n_565), .Y(n_562) );
INVx1_ASAP7_75t_L g517 ( .A(n_212), .Y(n_517) );
INVx1_ASAP7_75t_L g473 ( .A(n_213), .Y(n_473) );
AOI22xp33_ASAP7_75t_SL g753 ( .A1(n_214), .A2(n_250), .B1(n_602), .B2(n_661), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_216), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_217), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_220), .A2(n_247), .B1(n_390), .B2(n_438), .Y(n_671) );
INVx1_ASAP7_75t_L g852 ( .A(n_224), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_226), .Y(n_599) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_228), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_229), .B(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_SL g743 ( .A(n_231), .B(n_379), .Y(n_743) );
INVx1_ASAP7_75t_L g412 ( .A(n_234), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_235), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_236), .B(n_378), .Y(n_854) );
AOI22xp5_ASAP7_75t_SL g488 ( .A1(n_237), .A2(n_268), .B1(n_348), .B2(n_489), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_239), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_240), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_241), .A2(n_252), .B1(n_379), .B2(n_665), .Y(n_664) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_242), .A2(n_620), .B1(n_621), .B2(n_652), .Y(n_619) );
INVx1_ASAP7_75t_L g652 ( .A(n_242), .Y(n_652) );
INVx1_ASAP7_75t_L g407 ( .A(n_243), .Y(n_407) );
INVx1_ASAP7_75t_L g796 ( .A(n_246), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_256), .Y(n_499) );
INVx1_ASAP7_75t_L g292 ( .A(n_258), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_258), .Y(n_294) );
OA22x2_ASAP7_75t_L g555 ( .A1(n_264), .A2(n_556), .B1(n_557), .B2(n_581), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_264), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_265), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_266), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g271 ( .A(n_272), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_276), .Y(n_792) );
OAI21xp5_ASAP7_75t_L g838 ( .A1(n_277), .A2(n_791), .B(n_839), .Y(n_838) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_615), .B1(n_786), .B2(n_787), .C(n_788), .Y(n_280) );
INVx1_ASAP7_75t_L g786 ( .A(n_281), .Y(n_786) );
XOR2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_365), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
XOR2x2_ASAP7_75t_SL g283 ( .A(n_284), .B(n_364), .Y(n_283) );
NAND2x1p5_ASAP7_75t_L g284 ( .A(n_285), .B(n_334), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_286), .B(n_319), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_302), .C(n_308), .Y(n_286) );
BUFx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx4f_ASAP7_75t_L g379 ( .A(n_289), .Y(n_379) );
BUFx2_ASAP7_75t_L g576 ( .A(n_289), .Y(n_576) );
AND2x6_ASAP7_75t_L g289 ( .A(n_290), .B(n_298), .Y(n_289) );
AND2x4_ASAP7_75t_L g355 ( .A(n_290), .B(n_323), .Y(n_355) );
AND2x2_ASAP7_75t_L g358 ( .A(n_290), .B(n_342), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_290), .B(n_298), .Y(n_410) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_290), .B(n_342), .Y(n_471) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
OR2x2_ASAP7_75t_L g307 ( .A(n_291), .B(n_295), .Y(n_307) );
INVx2_ASAP7_75t_L g313 ( .A(n_291), .Y(n_313) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
AND2x2_ASAP7_75t_L g322 ( .A(n_291), .B(n_296), .Y(n_322) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g297 ( .A(n_294), .Y(n_297) );
AND2x2_ASAP7_75t_L g343 ( .A(n_295), .B(n_313), .Y(n_343) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g314 ( .A(n_296), .B(n_301), .Y(n_314) );
AND2x4_ASAP7_75t_L g305 ( .A(n_298), .B(n_306), .Y(n_305) );
AND2x4_ASAP7_75t_L g361 ( .A(n_298), .B(n_343), .Y(n_361) );
INVx1_ASAP7_75t_L g406 ( .A(n_298), .Y(n_406) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g312 ( .A(n_299), .Y(n_312) );
INVx1_ASAP7_75t_L g324 ( .A(n_299), .Y(n_324) );
INVx1_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_299), .B(n_301), .Y(n_351) );
AND2x2_ASAP7_75t_L g323 ( .A(n_300), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g342 ( .A(n_301), .B(n_333), .Y(n_342) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
INVx5_ASAP7_75t_L g378 ( .A(n_304), .Y(n_378) );
INVx2_ASAP7_75t_L g665 ( .A(n_304), .Y(n_665) );
INVx2_ASAP7_75t_L g745 ( .A(n_304), .Y(n_745) );
INVx4_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x6_ASAP7_75t_L g339 ( .A(n_306), .B(n_323), .Y(n_339) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g405 ( .A(n_307), .B(n_406), .Y(n_405) );
INVx4_ASAP7_75t_L g456 ( .A(n_309), .Y(n_456) );
INVx2_ASAP7_75t_L g506 ( .A(n_309), .Y(n_506) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx4f_ASAP7_75t_SL g376 ( .A(n_310), .Y(n_376) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_310), .Y(n_421) );
BUFx2_ASAP7_75t_L g593 ( .A(n_310), .Y(n_593) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_310), .Y(n_732) );
AND2x4_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
INVx1_ASAP7_75t_L g424 ( .A(n_313), .Y(n_424) );
AND2x4_ASAP7_75t_L g316 ( .A(n_314), .B(n_317), .Y(n_316) );
AND2x4_ASAP7_75t_L g328 ( .A(n_314), .B(n_329), .Y(n_328) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_314), .B(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g578 ( .A(n_316), .Y(n_578) );
BUFx2_ASAP7_75t_L g667 ( .A(n_316), .Y(n_667) );
INVx1_ASAP7_75t_L g705 ( .A(n_316), .Y(n_705) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x6_ASAP7_75t_L g363 ( .A(n_318), .B(n_351), .Y(n_363) );
OAI21xp5_ASAP7_75t_SL g319 ( .A1(n_320), .A2(n_325), .B(n_326), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_320), .A2(n_371), .B(n_372), .Y(n_370) );
OAI21xp5_ASAP7_75t_SL g739 ( .A1(n_320), .A2(n_740), .B(n_741), .Y(n_739) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g414 ( .A(n_321), .Y(n_414) );
INVx2_ASAP7_75t_SL g454 ( .A(n_321), .Y(n_454) );
INVx4_ASAP7_75t_L g504 ( .A(n_321), .Y(n_504) );
BUFx3_ASAP7_75t_L g524 ( .A(n_321), .Y(n_524) );
INVx2_ASAP7_75t_L g807 ( .A(n_321), .Y(n_807) );
AND2x6_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AND2x4_ASAP7_75t_L g331 ( .A(n_322), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g536 ( .A(n_322), .Y(n_536) );
AND2x2_ASAP7_75t_L g347 ( .A(n_323), .B(n_343), .Y(n_347) );
BUFx4f_ASAP7_75t_SL g580 ( .A(n_327), .Y(n_580) );
INVx2_ASAP7_75t_L g595 ( .A(n_327), .Y(n_595) );
BUFx12f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_328), .Y(n_416) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_328), .Y(n_528) );
BUFx3_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_SL g373 ( .A(n_331), .Y(n_373) );
BUFx6f_ASAP7_75t_L g417 ( .A(n_331), .Y(n_417) );
INVx1_ASAP7_75t_L g537 ( .A(n_332), .Y(n_537) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NOR2x1_ASAP7_75t_L g334 ( .A(n_335), .B(n_352), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_344), .Y(n_335) );
INVx2_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx5_ASAP7_75t_SL g384 ( .A(n_338), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_338), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g680 ( .A(n_338), .Y(n_680) );
INVx4_ASAP7_75t_L g775 ( .A(n_338), .Y(n_775) );
INVx2_ASAP7_75t_L g845 ( .A(n_338), .Y(n_845) );
INVx11_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx11_ASAP7_75t_L g490 ( .A(n_339), .Y(n_490) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx3_ASAP7_75t_L g429 ( .A(n_341), .Y(n_429) );
BUFx3_ASAP7_75t_L g483 ( .A(n_341), .Y(n_483) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_342), .B(n_343), .Y(n_474) );
AND2x4_ASAP7_75t_L g349 ( .A(n_343), .B(n_350), .Y(n_349) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI22xp5_ASAP7_75t_SL g463 ( .A1(n_346), .A2(n_388), .B1(n_464), .B2(n_465), .Y(n_463) );
INVx3_ASAP7_75t_L g486 ( .A(n_346), .Y(n_486) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx2_ASAP7_75t_SL g431 ( .A(n_347), .Y(n_431) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_347), .Y(n_551) );
BUFx3_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx3_ASAP7_75t_L g432 ( .A(n_349), .Y(n_432) );
INVx1_ASAP7_75t_L g469 ( .A(n_349), .Y(n_469) );
BUFx2_ASAP7_75t_SL g541 ( .A(n_349), .Y(n_541) );
BUFx2_ASAP7_75t_L g572 ( .A(n_349), .Y(n_572) );
BUFx3_ASAP7_75t_L g607 ( .A(n_349), .Y(n_607) );
BUFx2_ASAP7_75t_SL g693 ( .A(n_349), .Y(n_693) );
AND2x2_ASAP7_75t_L g462 ( .A(n_350), .B(n_424), .Y(n_462) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_359), .Y(n_352) );
INVx1_ASAP7_75t_L g634 ( .A(n_354), .Y(n_634) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx6_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
BUFx3_ASAP7_75t_L g437 ( .A(n_355), .Y(n_437) );
BUFx3_ASAP7_75t_L g602 ( .A(n_355), .Y(n_602) );
INVx5_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g438 ( .A(n_357), .Y(n_438) );
INVx3_ASAP7_75t_L g484 ( .A(n_357), .Y(n_484) );
BUFx3_ASAP7_75t_L g544 ( .A(n_357), .Y(n_544) );
INVx4_ASAP7_75t_L g564 ( .A(n_357), .Y(n_564) );
INVx1_ASAP7_75t_L g750 ( .A(n_357), .Y(n_750) );
INVx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx4_ASAP7_75t_L g571 ( .A(n_360), .Y(n_571) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g440 ( .A(n_361), .Y(n_440) );
INVx2_ASAP7_75t_L g459 ( .A(n_361), .Y(n_459) );
BUFx3_ASAP7_75t_L g670 ( .A(n_361), .Y(n_670) );
BUFx3_ASAP7_75t_L g726 ( .A(n_361), .Y(n_726) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
INVx6_ASAP7_75t_SL g390 ( .A(n_363), .Y(n_390) );
INVx1_ASAP7_75t_L g441 ( .A(n_363), .Y(n_441) );
INVx1_ASAP7_75t_SL g698 ( .A(n_363), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_392), .B2(n_614), .Y(n_365) );
INVx3_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
XOR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_391), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_369), .B(n_380), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_374), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g709 ( .A(n_376), .Y(n_709) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_378), .Y(n_575) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_378), .Y(n_650) );
INVx1_ASAP7_75t_L g817 ( .A(n_379), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_381), .B(n_385), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_L g632 ( .A(n_384), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g547 ( .A(n_388), .Y(n_547) );
INVx2_ASAP7_75t_L g662 ( .A(n_388), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_388), .A2(n_773), .B1(n_774), .B2(n_776), .Y(n_772) );
BUFx2_ASAP7_75t_L g565 ( .A(n_390), .Y(n_565) );
BUFx2_ASAP7_75t_L g604 ( .A(n_390), .Y(n_604) );
INVx1_ASAP7_75t_L g614 ( .A(n_392), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_509), .B2(n_613), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AO22x2_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B1(n_442), .B2(n_508), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_425), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_411), .C(n_418), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B1(n_407), .B2(n_408), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g500 ( .A1(n_404), .A2(n_501), .B(n_502), .Y(n_500) );
BUFx6f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g446 ( .A1(n_405), .A2(n_447), .B(n_448), .Y(n_446) );
INVx2_ASAP7_75t_L g519 ( .A(n_405), .Y(n_519) );
OAI22xp5_ASAP7_75t_SL g758 ( .A1(n_405), .A2(n_409), .B1(n_759), .B2(n_760), .Y(n_758) );
OAI221xp5_ASAP7_75t_SL g700 ( .A1(n_408), .A2(n_518), .B1(n_701), .B2(n_702), .C(n_703), .Y(n_700) );
BUFx3_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_409), .A2(n_423), .B1(n_450), .B2(n_451), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_409), .A2(n_517), .B1(n_518), .B2(n_520), .Y(n_516) );
OA211x2_ASAP7_75t_L g727 ( .A1(n_409), .A2(n_728), .B(n_729), .C(n_730), .Y(n_727) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g495 ( .A(n_410), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B(n_415), .Y(n_411) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx4f_ASAP7_75t_L g646 ( .A(n_416), .Y(n_646) );
INVx1_ASAP7_75t_L g811 ( .A(n_416), .Y(n_811) );
INVx1_ASAP7_75t_SL g707 ( .A(n_417), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B1(n_422), .B2(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_421), .Y(n_526) );
INVx4_ASAP7_75t_L g498 ( .A(n_423), .Y(n_498) );
BUFx3_ASAP7_75t_L g531 ( .A(n_423), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_426), .B(n_433), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_430), .Y(n_426) );
BUFx4f_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g687 ( .A(n_429), .Y(n_687) );
INVx1_ASAP7_75t_L g637 ( .A(n_431), .Y(n_637) );
INVx2_ASAP7_75t_L g627 ( .A(n_432), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_434), .B(n_439), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g690 ( .A(n_440), .Y(n_690) );
INVx2_ASAP7_75t_L g508 ( .A(n_442), .Y(n_508) );
XOR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_478), .Y(n_442) );
XNOR2x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_477), .Y(n_443) );
AND3x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_457), .C(n_466), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .C(n_452), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_454), .B1(n_455), .B2(n_456), .Y(n_452) );
OAI222xp33_ASAP7_75t_L g708 ( .A1(n_454), .A2(n_709), .B1(n_710), .B2(n_711), .C1(n_712), .C2(n_713), .Y(n_708) );
INVx3_ASAP7_75t_L g645 ( .A(n_456), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_463), .Y(n_457) );
OAI21xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_460), .B(n_461), .Y(n_458) );
INVx2_ASAP7_75t_L g540 ( .A(n_459), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_472), .C(n_475), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_470), .B2(n_471), .Y(n_467) );
BUFx2_ASAP7_75t_R g825 ( .A(n_471), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g640 ( .A(n_474), .Y(n_640) );
XNOR2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
NAND3x1_ASAP7_75t_SL g480 ( .A(n_481), .B(n_487), .C(n_492), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g561 ( .A(n_483), .Y(n_561) );
BUFx2_ASAP7_75t_L g820 ( .A(n_483), .Y(n_820) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_491), .Y(n_487) );
INVx1_ASAP7_75t_L g831 ( .A(n_489), .Y(n_831) );
INVx4_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx2_ASAP7_75t_SL g546 ( .A(n_490), .Y(n_546) );
INVx3_ASAP7_75t_L g661 ( .A(n_490), .Y(n_661) );
NOR3xp33_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .C(n_503), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_496), .B1(n_497), .B2(n_499), .Y(n_493) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_494), .A2(n_587), .B1(n_588), .B2(n_589), .Y(n_586) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g853 ( .A(n_495), .Y(n_853) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_497), .A2(n_765), .B1(n_766), .B2(n_767), .Y(n_764) );
INVx3_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g598 ( .A(n_498), .Y(n_598) );
OAI22xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_505), .B1(n_506), .B2(n_507), .Y(n_503) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_504), .A2(n_643), .B(n_644), .Y(n_642) );
INVx4_ASAP7_75t_L g673 ( .A(n_504), .Y(n_673) );
OAI21xp5_ASAP7_75t_SL g761 ( .A1(n_504), .A2(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g613 ( .A(n_509), .Y(n_613) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_554), .B2(n_612), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_SL g552 ( .A(n_514), .Y(n_552) );
AND2x2_ASAP7_75t_SL g514 ( .A(n_515), .B(n_538), .Y(n_514) );
NOR3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_521), .C(n_529), .Y(n_515) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g588 ( .A(n_519), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B(n_525), .Y(n_521) );
OAI21xp33_ASAP7_75t_L g590 ( .A1(n_523), .A2(n_591), .B(n_592), .Y(n_590) );
INVx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_SL g809 ( .A(n_526), .Y(n_809) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g712 ( .A(n_528), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_531), .B1(n_532), .B2(n_533), .Y(n_529) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_535), .A2(n_597), .B1(n_598), .B2(n_599), .Y(n_596) );
BUFx2_ASAP7_75t_L g766 ( .A(n_535), .Y(n_766) );
OR2x6_ASAP7_75t_L g535 ( .A(n_536), .B(n_537), .Y(n_535) );
AND4x1_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .C(n_545), .D(n_548), .Y(n_538) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx3_ASAP7_75t_L g568 ( .A(n_551), .Y(n_568) );
BUFx3_ASAP7_75t_L g685 ( .A(n_551), .Y(n_685) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_551), .Y(n_849) );
INVx1_ASAP7_75t_L g612 ( .A(n_554), .Y(n_612) );
AOI22x1_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_582), .B1(n_610), .B2(n_611), .Y(n_554) );
INVx1_ASAP7_75t_L g610 ( .A(n_555), .Y(n_610) );
INVx1_ASAP7_75t_SL g581 ( .A(n_557), .Y(n_581) );
NAND4xp75_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .C(n_573), .D(n_579), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_562), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_564), .Y(n_629) );
INVx2_ASAP7_75t_L g697 ( .A(n_564), .Y(n_697) );
INVx1_ASAP7_75t_L g827 ( .A(n_565), .Y(n_827) );
AND2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_569), .Y(n_566) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx4_ASAP7_75t_L g625 ( .A(n_571), .Y(n_625) );
AND2x2_ASAP7_75t_SL g573 ( .A(n_574), .B(n_577), .Y(n_573) );
INVx1_ASAP7_75t_L g611 ( .A(n_582), .Y(n_611) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
XNOR2xp5_ASAP7_75t_L g618 ( .A(n_583), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g608 ( .A(n_584), .Y(n_608) );
AND2x2_ASAP7_75t_SL g584 ( .A(n_585), .B(n_600), .Y(n_584) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_590), .C(n_596), .Y(n_585) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AND4x1_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .C(n_605), .D(n_606), .Y(n_600) );
INVx1_ASAP7_75t_L g682 ( .A(n_602), .Y(n_682) );
INVx1_ASAP7_75t_L g787 ( .A(n_615), .Y(n_787) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_653), .B2(n_785), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_SL g621 ( .A(n_622), .B(n_641), .Y(n_621) );
NOR3xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_630), .C(n_635), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_628), .Y(n_623) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B1(n_638), .B2(n_639), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_637), .A2(n_639), .B1(n_778), .B2(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_647), .Y(n_641) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .C(n_651), .Y(n_647) );
INVx1_ASAP7_75t_L g785 ( .A(n_653), .Y(n_785) );
XOR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_717), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B1(n_675), .B2(n_716), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
XOR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_674), .Y(n_656) );
NAND4xp75_ASAP7_75t_L g657 ( .A(n_658), .B(n_663), .C(n_668), .D(n_672), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_SL g663 ( .A(n_664), .B(n_666), .Y(n_663) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_671), .Y(n_668) );
HB1xp67_ASAP7_75t_L g822 ( .A(n_670), .Y(n_822) );
INVx1_ASAP7_75t_L g716 ( .A(n_675), .Y(n_716) );
INVx1_ASAP7_75t_L g715 ( .A(n_676), .Y(n_715) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_699), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g677 ( .A(n_678), .B(n_688), .Y(n_677) );
OAI221xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_681), .B1(n_682), .B2(n_683), .C(n_684), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_691), .B1(n_692), .B2(n_694), .C(n_695), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NOR2xp33_ASAP7_75t_SL g699 ( .A(n_700), .B(n_708), .Y(n_699) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AO22x1_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_734), .B1(n_735), .B2(n_784), .Y(n_717) );
INVx2_ASAP7_75t_SL g784 ( .A(n_718), .Y(n_784) );
XOR2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_733), .Y(n_718) );
NAND4xp75_ASAP7_75t_L g719 ( .A(n_720), .B(n_723), .C(n_727), .D(n_731), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AO22x2_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_755), .B1(n_782), .B2(n_783), .Y(n_735) );
INVx4_ASAP7_75t_SL g782 ( .A(n_736), .Y(n_782) );
XOR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_754), .Y(n_736) );
NAND3x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_747), .C(n_751), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .C(n_746), .Y(n_742) );
AND2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g783 ( .A(n_755), .Y(n_783) );
INVx1_ASAP7_75t_L g780 ( .A(n_756), .Y(n_780) );
AND2x2_ASAP7_75t_L g756 ( .A(n_757), .B(n_768), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_758), .B(n_761), .C(n_764), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_772), .C(n_777), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .Y(n_769) );
INVx1_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
NOR2x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_794), .Y(n_789) );
OR2x2_ASAP7_75t_SL g859 ( .A(n_790), .B(n_795), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_792), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_792), .B(n_836), .Y(n_839) );
CKINVDCx16_ASAP7_75t_R g836 ( .A(n_793), .Y(n_836) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_796), .B(n_797), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
OAI322xp33_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_833), .A3(n_834), .B1(n_837), .B2(n_840), .C1(n_841), .C2(n_857), .Y(n_801) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NAND3x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_818), .C(n_823), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_813), .Y(n_805) );
OAI222xp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_808), .B1(n_809), .B2(n_810), .C1(n_811), .C2(n_812), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_821), .Y(n_818) );
OAI22xp5_ASAP7_75t_SL g824 ( .A1(n_825), .A2(n_826), .B1(n_827), .B2(n_828), .Y(n_824) );
NOR2xp33_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_838), .Y(n_837) );
NAND4xp75_ASAP7_75t_L g842 ( .A(n_843), .B(n_847), .C(n_851), .D(n_856), .Y(n_842) );
AND2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_846), .Y(n_843) );
AND2x2_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
OA211x2_ASAP7_75t_L g851 ( .A1(n_852), .A2(n_853), .B(n_854), .C(n_855), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g857 ( .A(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
endmodule