module fake_jpeg_29359_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx12_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_19),
.B1(n_33),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_14),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_12),
.Y(n_48)
);

INVx5_ASAP7_75t_SL g49 ( 
.A(n_40),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_50),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_0),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_62),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_61),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_34),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_71),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_59),
.A2(n_40),
.B1(n_42),
.B2(n_37),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_72),
.B1(n_6),
.B2(n_7),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_40),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_66),
.A2(n_38),
.B1(n_34),
.B2(n_21),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_76),
.B(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_54),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_5),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_1),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_81),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_92),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_91),
.B1(n_71),
.B2(n_68),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_8),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_25),
.B1(n_30),
.B2(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_72),
.B1(n_71),
.B2(n_79),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_R g100 ( 
.A(n_94),
.B(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_95),
.B(n_90),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_75),
.Y(n_97)
);

MAJx2_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_85),
.C(n_84),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_101),
.B(n_102),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_97),
.A2(n_83),
.B(n_93),
.Y(n_103)
);

AO221x1_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_99),
.B1(n_94),
.B2(n_96),
.C(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_9),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_10),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_10),
.B(n_22),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_108),
.A2(n_23),
.B(n_24),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_104),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_28),
.Y(n_112)
);


endmodule