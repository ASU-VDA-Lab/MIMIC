module fake_jpeg_28190_n_39 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_6),
.B(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_0),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_10),
.B(n_0),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_5),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_19),
.C(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_2),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_20),
.A2(n_13),
.B1(n_14),
.B2(n_11),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_28),
.B1(n_13),
.B2(n_17),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_28),
.C(n_15),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_26),
.C(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_37),
.B(n_25),
.Y(n_38)
);

OAI311xp33_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_35),
.A3(n_36),
.B1(n_37),
.C1(n_34),
.Y(n_39)
);


endmodule