module fake_netlist_6_4653_n_1775 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1775);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1775;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_26),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_47),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_83),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_36),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_103),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_28),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_55),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_49),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_39),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_3),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_10),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_38),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_85),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_17),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_138),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_31),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_87),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_37),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_23),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_140),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_116),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_58),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_43),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_128),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_37),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_55),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_54),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_48),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_27),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_101),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_108),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_14),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_23),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_89),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_49),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_9),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_124),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_142),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_62),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_152),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_150),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_48),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_44),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_69),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_79),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_21),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_74),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_15),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_20),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_36),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_21),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_46),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_104),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_77),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_70),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_94),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_148),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_41),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_3),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_119),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_30),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_42),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_80),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_43),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_93),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_1),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_100),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_38),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_34),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_73),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_31),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_97),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_27),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_14),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_40),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_9),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_0),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_105),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_90),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_120),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_4),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_76),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_15),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_133),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_53),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_53),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_114),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_41),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_141),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_99),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_88),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_39),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_20),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_61),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_11),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_35),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_131),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_113),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_35),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_81),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_107),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_44),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_143),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_54),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_98),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_11),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_45),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_2),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_134),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_92),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_71),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_16),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_135),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_24),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_16),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_32),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_33),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_109),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_226),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_159),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_226),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_211),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_226),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_178),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_226),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_155),
.B(n_0),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_159),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_161),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_180),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_164),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_305),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_249),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_165),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_165),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_1),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_200),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_4),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_155),
.B(n_5),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_214),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_166),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_163),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_240),
.B(n_5),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_163),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_263),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_240),
.B(n_6),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_264),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_174),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_175),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_168),
.Y(n_342)
);

INVxp33_ASAP7_75t_SL g343 ( 
.A(n_276),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_182),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_184),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_189),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_189),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_168),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_188),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_171),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_196),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_251),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_190),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_171),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_177),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_204),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_251),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_185),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_183),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_206),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_208),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_183),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_212),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_156),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_213),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_216),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_221),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_191),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_229),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_198),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_235),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_198),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_237),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_306),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_366),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_308),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_359),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_325),
.B(n_196),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_262),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_347),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_347),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_332),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_352),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_332),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

INVx6_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_334),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_324),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_326),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_333),
.B(n_270),
.Y(n_415)
);

CKINVDCx14_ASAP7_75t_R g416 ( 
.A(n_341),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_336),
.B(n_277),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_325),
.B(n_258),
.Y(n_418)
);

INVx6_ASAP7_75t_L g419 ( 
.A(n_313),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_327),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_351),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_327),
.Y(n_423)
);

BUFx8_ASAP7_75t_L g424 ( 
.A(n_335),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_L g427 ( 
.A(n_321),
.B(n_157),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_328),
.B(n_193),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_356),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_321),
.B(n_193),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_357),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

CKINVDCx11_ASAP7_75t_R g435 ( 
.A(n_311),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_361),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_361),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_364),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_359),
.B(n_249),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_315),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_369),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_372),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_372),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_380),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_388),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_316),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_418),
.B(n_196),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_428),
.B(n_318),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_419),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_L g453 ( 
.A1(n_440),
.A2(n_320),
.B1(n_309),
.B2(n_353),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_380),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_331),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_389),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_348),
.C(n_307),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_397),
.B(n_337),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_419),
.A2(n_343),
.B1(n_335),
.B2(n_313),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_388),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_419),
.A2(n_329),
.B1(n_199),
.B2(n_173),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_431),
.B(n_339),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_431),
.B(n_340),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_419),
.A2(n_329),
.B1(n_199),
.B2(n_173),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_382),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_419),
.A2(n_290),
.B1(n_248),
.B2(n_256),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_385),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_434),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_388),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_419),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_350),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_440),
.B(n_354),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_395),
.A2(n_242),
.B1(n_222),
.B2(n_207),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_415),
.B(n_417),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_417),
.B(n_362),
.Y(n_478)
);

INVx4_ASAP7_75t_L g479 ( 
.A(n_405),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_379),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_385),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_389),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_379),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_399),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_379),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_416),
.B(n_317),
.Y(n_492)
);

INVxp33_ASAP7_75t_SL g493 ( 
.A(n_381),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_392),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_435),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_399),
.B(n_363),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_395),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_434),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_390),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_383),
.Y(n_501)
);

INVx6_ASAP7_75t_L g502 ( 
.A(n_405),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_379),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_390),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_427),
.B(n_365),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_424),
.B(n_367),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_424),
.B(n_368),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_418),
.B(n_374),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_418),
.B(n_196),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_383),
.B(n_373),
.Y(n_511)
);

OR2x6_ASAP7_75t_L g512 ( 
.A(n_400),
.B(n_258),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_400),
.B(n_377),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_395),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_434),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_395),
.Y(n_517)
);

INVx5_ASAP7_75t_L g518 ( 
.A(n_395),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_424),
.B(n_378),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_395),
.Y(n_521)
);

INVxp33_ASAP7_75t_SL g522 ( 
.A(n_424),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_416),
.B(n_330),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_434),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_395),
.B(n_196),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_387),
.B(n_258),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_434),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_395),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_443),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_387),
.B(n_210),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_387),
.B(n_344),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_403),
.B(n_210),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_403),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_387),
.B(n_287),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_401),
.B(n_287),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_438),
.A2(n_222),
.B1(n_256),
.B2(n_304),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_443),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_401),
.B(n_160),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

INVx4_ASAP7_75t_L g542 ( 
.A(n_405),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_438),
.A2(n_268),
.B1(n_248),
.B2(n_304),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_443),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_443),
.Y(n_545)
);

INVx5_ASAP7_75t_L g546 ( 
.A(n_405),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_409),
.B(n_185),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_424),
.Y(n_548)
);

INVx8_ASAP7_75t_L g549 ( 
.A(n_401),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_445),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_445),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_409),
.B(n_377),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_401),
.B(n_376),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_445),
.Y(n_555)
);

AND2x6_ASAP7_75t_L g556 ( 
.A(n_401),
.B(n_196),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_410),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_445),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_405),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_438),
.A2(n_246),
.B1(n_242),
.B2(n_279),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_445),
.Y(n_561)
);

AO22x2_ASAP7_75t_L g562 ( 
.A1(n_438),
.A2(n_279),
.B1(n_268),
.B2(n_272),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_438),
.A2(n_246),
.B1(n_207),
.B2(n_233),
.Y(n_563)
);

CKINVDCx16_ASAP7_75t_R g564 ( 
.A(n_410),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_445),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_446),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_446),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_406),
.B(n_259),
.Y(n_568)
);

AND2x6_ASAP7_75t_L g569 ( 
.A(n_406),
.B(n_259),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_406),
.B(n_345),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_414),
.B(n_192),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_406),
.B(n_358),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_446),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_446),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_406),
.B(n_370),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_414),
.B(n_421),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_421),
.B(n_349),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_379),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_446),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_396),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_384),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_422),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_396),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_396),
.B(n_187),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_402),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_402),
.B(n_202),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_384),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_402),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_407),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_422),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_407),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_426),
.A2(n_288),
.B1(n_290),
.B2(n_302),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_578),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_578),
.Y(n_597)
);

BUFx5_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_477),
.B(n_405),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_474),
.B(n_371),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_375),
.Y(n_601)
);

BUFx12f_ASAP7_75t_SL g602 ( 
.A(n_512),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_455),
.B(n_255),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_513),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_484),
.B(n_259),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_484),
.B(n_259),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_582),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_585),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_534),
.B(n_592),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_513),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_585),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_466),
.B(n_232),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_488),
.B(n_291),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_495),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_488),
.B(n_234),
.Y(n_615)
);

INVx4_ASAP7_75t_L g616 ( 
.A(n_452),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_534),
.B(n_407),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g618 ( 
.A(n_452),
.B(n_338),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_592),
.B(n_407),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_449),
.B(n_459),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_562),
.A2(n_294),
.B1(n_272),
.B2(n_273),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_587),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_426),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_498),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_532),
.B(n_299),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_570),
.B(n_573),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_473),
.B(n_540),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_484),
.B(n_259),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_553),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_473),
.B(n_407),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_509),
.B(n_407),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_509),
.B(n_407),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_557),
.B(n_408),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_511),
.B(n_209),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_456),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_522),
.B(n_231),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_517),
.B(n_192),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_484),
.B(n_259),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_557),
.B(n_408),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_495),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_584),
.B(n_447),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_408),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_447),
.B(n_408),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_517),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_579),
.B(n_429),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_454),
.B(n_408),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_505),
.B(n_280),
.Y(n_648)
);

INVxp67_ASAP7_75t_SL g649 ( 
.A(n_471),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_553),
.Y(n_650)
);

AO22x2_ASAP7_75t_L g651 ( 
.A1(n_451),
.A2(n_267),
.B1(n_195),
.B2(n_201),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_453),
.B(n_281),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_481),
.B(n_282),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_590),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_454),
.B(n_408),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_460),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_554),
.A2(n_284),
.B1(n_285),
.B2(n_289),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_579),
.B(n_429),
.Y(n_658)
);

OR2x2_ASAP7_75t_L g659 ( 
.A(n_501),
.B(n_430),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_461),
.A2(n_154),
.B1(n_158),
.B2(n_223),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_577),
.B(n_293),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_464),
.B(n_193),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_L g663 ( 
.A(n_463),
.B(n_253),
.C(n_205),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_467),
.B(n_193),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_562),
.A2(n_273),
.B1(n_274),
.B2(n_288),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_562),
.A2(n_476),
.B1(n_528),
.B2(n_547),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_493),
.B(n_430),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_547),
.B(n_432),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_590),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_460),
.B(n_408),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_495),
.B(n_432),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_468),
.B(n_411),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_497),
.B(n_167),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_493),
.B(n_433),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_549),
.A2(n_442),
.B(n_439),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_468),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_470),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_484),
.B(n_154),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_484),
.B(n_158),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_470),
.B(n_411),
.Y(n_680)
);

NAND2x1p5_ASAP7_75t_L g681 ( 
.A(n_528),
.B(n_195),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_518),
.B(n_223),
.Y(n_682)
);

O2A1O1Ixp33_ASAP7_75t_L g683 ( 
.A1(n_525),
.A2(n_444),
.B(n_433),
.C(n_436),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_518),
.B(n_247),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_482),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_475),
.A2(n_220),
.B1(n_297),
.B2(n_296),
.Y(n_686)
);

BUFx12f_ASAP7_75t_SL g687 ( 
.A(n_512),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_547),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_483),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_533),
.A2(n_220),
.B1(n_297),
.B2(n_296),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_483),
.B(n_411),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_533),
.A2(n_271),
.B1(n_217),
.B2(n_227),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_491),
.Y(n_693)
);

AND2x6_ASAP7_75t_SL g694 ( 
.A(n_512),
.B(n_233),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_571),
.B(n_436),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_494),
.B(n_411),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_494),
.A2(n_247),
.B(n_201),
.C(n_269),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_514),
.A2(n_217),
.B(n_227),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_518),
.B(n_243),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_508),
.B(n_411),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVxp67_ASAP7_75t_SL g702 ( 
.A(n_471),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_469),
.A2(n_269),
.B1(n_245),
.B2(n_250),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_549),
.B(n_411),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_518),
.B(n_243),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_514),
.A2(n_271),
.B1(n_250),
.B2(n_252),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_521),
.A2(n_245),
.B1(n_252),
.B2(n_260),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_533),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_518),
.B(n_260),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_549),
.B(n_411),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_521),
.A2(n_267),
.B(n_444),
.C(n_437),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_471),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_458),
.B(n_586),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_456),
.B(n_437),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_588),
.B(n_169),
.Y(n_715)
);

AND2x4_ASAP7_75t_SL g716 ( 
.A(n_486),
.B(n_249),
.Y(n_716)
);

AOI221xp5_ASAP7_75t_L g717 ( 
.A1(n_594),
.A2(n_254),
.B1(n_283),
.B2(n_302),
.C(n_274),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_512),
.B(n_172),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_549),
.B(n_412),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_565),
.B(n_412),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_485),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_571),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_565),
.B(n_567),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_479),
.B(n_412),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_485),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_562),
.A2(n_292),
.B1(n_298),
.B2(n_294),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_448),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_567),
.B(n_412),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_530),
.B(n_412),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_486),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_448),
.Y(n_732)
);

O2A1O1Ixp33_ASAP7_75t_L g733 ( 
.A1(n_525),
.A2(n_292),
.B(n_298),
.C(n_300),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_535),
.B(n_412),
.Y(n_734)
);

BUFx6f_ASAP7_75t_SL g735 ( 
.A(n_486),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_548),
.B(n_425),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_536),
.B(n_412),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_548),
.B(n_425),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_526),
.B(n_413),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_462),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_462),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_583),
.B(n_413),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_472),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_479),
.B(n_413),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_506),
.B(n_249),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_472),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_479),
.B(n_542),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_542),
.B(n_413),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_489),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_489),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_507),
.B(n_179),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_519),
.B(n_181),
.Y(n_752)
);

NOR2xp67_ASAP7_75t_L g753 ( 
.A(n_591),
.B(n_425),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_520),
.B(n_186),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_542),
.B(n_413),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_559),
.B(n_450),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_559),
.B(n_450),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_450),
.A2(n_300),
.B1(n_442),
.B2(n_439),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_500),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_496),
.B(n_244),
.C(n_197),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_537),
.B(n_442),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_543),
.B(n_439),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_559),
.B(n_413),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_620),
.B(n_546),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_753),
.A2(n_566),
.B(n_544),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_676),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_603),
.A2(n_502),
.B1(n_560),
.B2(n_563),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_SL g768 ( 
.A(n_735),
.B(n_492),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_603),
.A2(n_599),
.B1(n_688),
.B2(n_666),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_634),
.A2(n_510),
.B1(n_450),
.B2(n_520),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_450),
.Y(n_771)
);

INVxp67_ASAP7_75t_SL g772 ( 
.A(n_624),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_635),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_598),
.B(n_546),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_623),
.B(n_492),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_747),
.A2(n_546),
.B(n_471),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_624),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_756),
.A2(n_546),
.B(n_471),
.Y(n_778)
);

NAND3xp33_ASAP7_75t_SL g779 ( 
.A(n_600),
.B(n_266),
.C(n_203),
.Y(n_779)
);

BUFx4f_ASAP7_75t_L g780 ( 
.A(n_726),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_757),
.A2(n_546),
.B(n_561),
.Y(n_781)
);

OAI21xp33_ASAP7_75t_L g782 ( 
.A1(n_613),
.A2(n_275),
.B(n_218),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_627),
.A2(n_561),
.B(n_499),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_715),
.B(n_450),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_L g785 ( 
.A1(n_688),
.A2(n_502),
.B1(n_541),
.B2(n_531),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_624),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_598),
.B(n_515),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_676),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_666),
.A2(n_502),
.B1(n_558),
.B2(n_541),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_598),
.B(n_545),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_677),
.Y(n_791)
);

BUFx12f_ASAP7_75t_L g792 ( 
.A(n_614),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_640),
.B(n_523),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_713),
.A2(n_544),
.B(n_524),
.C(n_527),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_601),
.B(n_524),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_677),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_715),
.B(n_450),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_SL g798 ( 
.A1(n_612),
.A2(n_550),
.B(n_527),
.C(n_529),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_693),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_744),
.A2(n_561),
.B(n_499),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_624),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_748),
.A2(n_561),
.B(n_499),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_714),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_631),
.A2(n_551),
.B(n_529),
.Y(n_804)
);

BUFx4f_ASAP7_75t_L g805 ( 
.A(n_671),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_641),
.B(n_510),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_609),
.B(n_510),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_718),
.A2(n_502),
.B1(n_572),
.B2(n_550),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_596),
.B(n_545),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_755),
.A2(n_561),
.B(n_499),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_644),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_717),
.B(n_238),
.C(n_194),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_615),
.B(n_510),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_693),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_713),
.A2(n_510),
.B1(n_539),
.B2(n_552),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_626),
.B(n_531),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_632),
.A2(n_575),
.B(n_538),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_644),
.Y(n_818)
);

OAI21x1_ASAP7_75t_L g819 ( 
.A1(n_725),
.A2(n_555),
.B(n_490),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_659),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_656),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_716),
.Y(n_822)
);

AO22x1_ASAP7_75t_L g823 ( 
.A1(n_751),
.A2(n_752),
.B1(n_673),
.B2(n_745),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_615),
.B(n_510),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_685),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_602),
.B(n_523),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_598),
.B(n_555),
.Y(n_827)
);

AOI22x1_ASAP7_75t_L g828 ( 
.A1(n_651),
.A2(n_551),
.B1(n_538),
.B2(n_539),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_595),
.Y(n_829)
);

O2A1O1Ixp33_ASAP7_75t_SL g830 ( 
.A1(n_711),
.A2(n_575),
.B(n_558),
.C(n_552),
.Y(n_830)
);

BUFx12f_ASAP7_75t_L g831 ( 
.A(n_694),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_597),
.B(n_566),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_645),
.B(n_219),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_644),
.B(n_499),
.Y(n_834)
);

AOI21x1_ASAP7_75t_L g835 ( 
.A1(n_725),
.A2(n_572),
.B(n_581),
.Y(n_835)
);

O2A1O1Ixp5_ASAP7_75t_L g836 ( 
.A1(n_698),
.A2(n_500),
.B(n_504),
.C(n_581),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_722),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_704),
.A2(n_516),
.B(n_574),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_598),
.B(n_574),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_723),
.A2(n_576),
.B1(n_593),
.B2(n_591),
.Y(n_840)
);

OAI21xp33_ASAP7_75t_SL g841 ( 
.A1(n_689),
.A2(n_576),
.B(n_593),
.Y(n_841)
);

NOR2x1_ASAP7_75t_L g842 ( 
.A(n_618),
.B(n_457),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_701),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_658),
.B(n_589),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_604),
.B(n_589),
.Y(n_845)
);

O2A1O1Ixp5_ASAP7_75t_L g846 ( 
.A1(n_660),
.A2(n_504),
.B(n_487),
.C(n_480),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_724),
.A2(n_580),
.B1(n_457),
.B2(n_465),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_607),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_751),
.A2(n_480),
.B(n_490),
.C(n_457),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_610),
.B(n_465),
.Y(n_850)
);

AOI21xp33_ASAP7_75t_L g851 ( 
.A1(n_673),
.A2(n_224),
.B(n_225),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_710),
.A2(n_516),
.B(n_465),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_L g853 ( 
.A(n_637),
.B(n_556),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_629),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_720),
.A2(n_763),
.B(n_729),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_650),
.B(n_580),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_607),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_613),
.B(n_580),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_653),
.B(n_228),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_668),
.B(n_695),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_608),
.Y(n_861)
);

INVx4_ASAP7_75t_L g862 ( 
.A(n_712),
.Y(n_862)
);

NOR3xp33_ASAP7_75t_L g863 ( 
.A(n_625),
.B(n_230),
.C(n_239),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_752),
.A2(n_480),
.B(n_487),
.C(n_490),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_668),
.B(n_516),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_695),
.B(n_487),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_761),
.B(n_503),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_667),
.B(n_241),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_674),
.B(n_257),
.Y(n_869)
);

AND2x4_ASAP7_75t_L g870 ( 
.A(n_708),
.B(n_503),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_739),
.A2(n_569),
.B(n_568),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_732),
.Y(n_872)
);

NAND2x1p5_ASAP7_75t_L g873 ( 
.A(n_616),
.B(n_516),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_762),
.B(n_503),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_754),
.B(n_616),
.Y(n_875)
);

NAND2x1p5_ASAP7_75t_L g876 ( 
.A(n_712),
.B(n_516),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_763),
.A2(n_391),
.B(n_384),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_732),
.Y(n_878)
);

INVxp67_ASAP7_75t_L g879 ( 
.A(n_653),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_721),
.A2(n_569),
.B(n_568),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_754),
.B(n_569),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_703),
.A2(n_404),
.B(n_568),
.C(n_556),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_742),
.A2(n_391),
.B(n_384),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_736),
.B(n_404),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_649),
.B(n_569),
.Y(n_885)
);

OAI21x1_ASAP7_75t_L g886 ( 
.A1(n_675),
.A2(n_404),
.B(n_568),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_651),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_630),
.A2(n_734),
.B(n_730),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_652),
.B(n_261),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_716),
.B(n_265),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_719),
.A2(n_278),
.B(n_286),
.C(n_295),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_740),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_702),
.B(n_569),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_621),
.A2(n_301),
.B1(n_303),
.B2(n_413),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_648),
.B(n_569),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_L g896 ( 
.A(n_719),
.B(n_663),
.C(n_661),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_621),
.A2(n_420),
.B1(n_423),
.B2(n_384),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_636),
.A2(n_420),
.B1(n_423),
.B2(n_393),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_740),
.B(n_568),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_737),
.A2(n_394),
.B(n_391),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_L g901 ( 
.A1(n_738),
.A2(n_568),
.B1(n_556),
.B2(n_423),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_617),
.A2(n_556),
.B(n_75),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_746),
.B(n_556),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_746),
.B(n_556),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_651),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_712),
.B(n_423),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_749),
.B(n_423),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_664),
.B(n_7),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_633),
.A2(n_394),
.B(n_393),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_760),
.B(n_420),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_759),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_420),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_611),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_662),
.B(n_420),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_639),
.A2(n_394),
.B(n_393),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_622),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_657),
.B(n_65),
.Y(n_917)
);

AOI21x1_ASAP7_75t_L g918 ( 
.A1(n_619),
.A2(n_394),
.B(n_393),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_643),
.A2(n_394),
.B(n_393),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_642),
.A2(n_394),
.B(n_393),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_712),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_686),
.A2(n_683),
.B(n_647),
.C(n_672),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_622),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_646),
.B(n_420),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_646),
.B(n_420),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_655),
.A2(n_394),
.B(n_393),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_654),
.B(n_391),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_670),
.A2(n_391),
.B(n_384),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_681),
.A2(n_7),
.B(n_8),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_637),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_680),
.A2(n_384),
.B(n_391),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_691),
.A2(n_391),
.B(n_63),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_654),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_669),
.B(n_8),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_690),
.B(n_115),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_696),
.A2(n_700),
.B(n_684),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_682),
.A2(n_151),
.B(n_147),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_637),
.Y(n_938)
);

AO21x1_ASAP7_75t_L g939 ( 
.A1(n_681),
.A2(n_10),
.B(n_12),
.Y(n_939)
);

BUFx2_ASAP7_75t_SL g940 ( 
.A(n_735),
.Y(n_940)
);

AO21x1_ASAP7_75t_L g941 ( 
.A1(n_706),
.A2(n_12),
.B(n_13),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_669),
.B(n_17),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_728),
.B(n_18),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_823),
.A2(n_707),
.B(n_750),
.C(n_743),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_805),
.B(n_769),
.Y(n_945)
);

INVx5_ASAP7_75t_L g946 ( 
.A(n_777),
.Y(n_946)
);

NOR2xp67_ASAP7_75t_SL g947 ( 
.A(n_940),
.B(n_709),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_889),
.A2(n_692),
.B(n_727),
.C(n_665),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_777),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_805),
.A2(n_665),
.B1(n_727),
.B2(n_758),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_SL g951 ( 
.A1(n_772),
.A2(n_684),
.B(n_682),
.Y(n_951)
);

BUFx4f_ASAP7_75t_L g952 ( 
.A(n_792),
.Y(n_952)
);

INVx5_ASAP7_75t_L g953 ( 
.A(n_777),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_875),
.A2(n_758),
.B1(n_741),
.B2(n_709),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_889),
.A2(n_637),
.B1(n_705),
.B2(n_699),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_795),
.B(n_705),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_879),
.B(n_687),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_766),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_795),
.A2(n_733),
.B(n_678),
.C(n_679),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_777),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_879),
.B(n_699),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_941),
.A2(n_638),
.B1(n_628),
.B2(n_606),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_780),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_811),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_764),
.A2(n_638),
.B(n_628),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_811),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_803),
.B(n_697),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_788),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_811),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_811),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_803),
.B(n_605),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_796),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_773),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_859),
.B(n_19),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_908),
.A2(n_19),
.B(n_22),
.C(n_25),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_791),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_935),
.B(n_78),
.Y(n_978)
);

AOI22xp33_ASAP7_75t_L g979 ( 
.A1(n_935),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_771),
.A2(n_86),
.B1(n_145),
.B2(n_136),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_829),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_833),
.B(n_33),
.Y(n_982)
);

NOR2x1_ASAP7_75t_R g983 ( 
.A(n_831),
.B(n_42),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_821),
.B(n_45),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_774),
.A2(n_95),
.B(n_125),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_825),
.B(n_46),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_774),
.A2(n_96),
.B(n_122),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_843),
.B(n_47),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_854),
.B(n_50),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_855),
.A2(n_82),
.B(n_118),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_772),
.A2(n_64),
.B1(n_117),
.B2(n_111),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_780),
.B(n_146),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_896),
.A2(n_106),
.B1(n_110),
.B2(n_52),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_851),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_773),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_824),
.A2(n_56),
.B1(n_57),
.B2(n_784),
.Y(n_997)
);

OAI21x1_ASAP7_75t_L g998 ( 
.A1(n_819),
.A2(n_765),
.B(n_918),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_814),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_764),
.A2(n_888),
.B(n_817),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_854),
.B(n_816),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_816),
.B(n_832),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_820),
.B(n_860),
.Y(n_1003)
);

OAI321xp33_ASAP7_75t_L g1004 ( 
.A1(n_812),
.A2(n_908),
.A3(n_779),
.B1(n_782),
.B2(n_869),
.C(n_868),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_826),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_804),
.A2(n_874),
.B(n_867),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_832),
.B(n_858),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_L g1008 ( 
.A1(n_868),
.A2(n_869),
.B(n_775),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_848),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_826),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_787),
.A2(n_827),
.B(n_790),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_844),
.B(n_809),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_809),
.B(n_896),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_863),
.A2(n_891),
.B(n_797),
.C(n_767),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_787),
.A2(n_827),
.B(n_790),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_860),
.B(n_884),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_837),
.B(n_890),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_839),
.A2(n_776),
.B(n_800),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_872),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_898),
.B(n_786),
.Y(n_1020)
);

NOR2xp33_ASAP7_75t_L g1021 ( 
.A(n_887),
.B(n_905),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_839),
.A2(n_810),
.B(n_802),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_878),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_892),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_786),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_911),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_898),
.B(n_801),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_884),
.B(n_818),
.Y(n_1028)
);

AO21x1_ASAP7_75t_L g1029 ( 
.A1(n_932),
.A2(n_881),
.B(n_942),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_801),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_793),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_870),
.B(n_818),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_822),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_916),
.Y(n_1034)
);

NAND2x1p5_ASAP7_75t_L g1035 ( 
.A(n_862),
.B(n_930),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_793),
.Y(n_1036)
);

OAI22xp5_ASAP7_75t_L g1037 ( 
.A1(n_815),
.A2(n_789),
.B1(n_905),
.B2(n_887),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_865),
.A2(n_866),
.B1(n_922),
.B2(n_807),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_857),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_779),
.B(n_863),
.C(n_910),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_793),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_845),
.B(n_850),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_861),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_930),
.B(n_938),
.Y(n_1044)
);

O2A1O1Ixp5_ASAP7_75t_SL g1045 ( 
.A1(n_943),
.A2(n_934),
.B(n_906),
.C(n_847),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_870),
.B(n_914),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_SL g1047 ( 
.A(n_768),
.B(n_939),
.C(n_929),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_862),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_865),
.A2(n_770),
.B1(n_806),
.B2(n_856),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_913),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_894),
.B(n_923),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_917),
.A2(n_794),
.B(n_841),
.C(n_936),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_842),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_846),
.A2(n_895),
.B(n_836),
.C(n_864),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_933),
.Y(n_1055)
);

NOR3xp33_ASAP7_75t_L g1056 ( 
.A(n_808),
.B(n_785),
.C(n_840),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_930),
.B(n_938),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_921),
.B(n_828),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_921),
.B(n_783),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_834),
.B(n_873),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_930),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_846),
.A2(n_836),
.B(n_849),
.C(n_882),
.Y(n_1062)
);

INVx3_ASAP7_75t_SL g1063 ( 
.A(n_938),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_938),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_927),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_885),
.A2(n_893),
.B1(n_876),
.B2(n_919),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_876),
.A2(n_880),
.B1(n_904),
.B2(n_903),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_906),
.B(n_897),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_SL g1069 ( 
.A1(n_871),
.A2(n_838),
.B(n_852),
.C(n_901),
.Y(n_1069)
);

NOR3xp33_ASAP7_75t_SL g1070 ( 
.A(n_937),
.B(n_899),
.C(n_907),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_835),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_912),
.B(n_924),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_778),
.A2(n_781),
.B(n_853),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_900),
.A2(n_883),
.B(n_920),
.C(n_915),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_909),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_926),
.A2(n_931),
.B(n_928),
.C(n_925),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_830),
.Y(n_1077)
);

INVx1_ASAP7_75t_SL g1078 ( 
.A(n_877),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_798),
.B(n_886),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_902),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_889),
.A2(n_603),
.B(n_634),
.C(n_455),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_823),
.B(n_620),
.Y(n_1082)
);

CKINVDCx14_ASAP7_75t_R g1083 ( 
.A(n_826),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_796),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_823),
.B(n_620),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_803),
.B(n_623),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_805),
.B(n_620),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_941),
.A2(n_603),
.B1(n_665),
.B2(n_621),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1000),
.A2(n_1081),
.B(n_1006),
.Y(n_1089)
);

AO32x2_ASAP7_75t_L g1090 ( 
.A1(n_1037),
.A2(n_997),
.A3(n_995),
.B1(n_1038),
.B2(n_1049),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1019),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_1004),
.A2(n_1008),
.B(n_975),
.C(n_1085),
.Y(n_1092)
);

AO21x2_ASAP7_75t_L g1093 ( 
.A1(n_1029),
.A2(n_1062),
.B(n_1054),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1073),
.A2(n_1052),
.B(n_1018),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1086),
.B(n_1017),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_1079),
.A2(n_1014),
.A3(n_1077),
.B(n_1066),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_1088),
.A2(n_979),
.B1(n_948),
.B2(n_950),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1023),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1020),
.A2(n_1027),
.B(n_1022),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1024),
.Y(n_1100)
);

BUFx4_ASAP7_75t_SL g1101 ( 
.A(n_963),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1082),
.B(n_996),
.Y(n_1102)
);

AO31x2_ASAP7_75t_L g1103 ( 
.A1(n_1079),
.A2(n_1067),
.A3(n_959),
.B(n_1058),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_1087),
.B(n_1001),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1026),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_944),
.A2(n_998),
.B(n_1076),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1020),
.A2(n_1027),
.B(n_1087),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_1040),
.A2(n_1088),
.B(n_978),
.C(n_961),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1069),
.A2(n_956),
.B(n_1059),
.Y(n_1109)
);

OAI21x1_ASAP7_75t_L g1110 ( 
.A1(n_1011),
.A2(n_1015),
.B(n_1074),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1074),
.A2(n_1076),
.B(n_965),
.Y(n_1111)
);

INVx1_ASAP7_75t_SL g1112 ( 
.A(n_973),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_1047),
.A2(n_945),
.B(n_978),
.C(n_994),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1040),
.A2(n_961),
.B(n_945),
.C(n_1013),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_952),
.Y(n_1115)
);

OA22x2_ASAP7_75t_L g1116 ( 
.A1(n_993),
.A2(n_1041),
.B1(n_974),
.B2(n_1031),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_1021),
.A2(n_1003),
.B1(n_1053),
.B2(n_982),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1046),
.B(n_957),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_957),
.B(n_1021),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1002),
.B(n_1007),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1069),
.A2(n_1042),
.B(n_1072),
.Y(n_1121)
);

AO21x2_ASAP7_75t_L g1122 ( 
.A1(n_1056),
.A2(n_1070),
.B(n_990),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1042),
.B(n_1016),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_954),
.A2(n_1078),
.B(n_1012),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_1033),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1075),
.A2(n_951),
.B(n_1044),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_1045),
.A2(n_1060),
.B(n_944),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1034),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_964),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_1005),
.B(n_1010),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_1044),
.A2(n_1056),
.B(n_1051),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_1083),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_SL g1133 ( 
.A(n_952),
.B(n_1030),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_1036),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_971),
.B(n_1065),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_980),
.A2(n_971),
.A3(n_986),
.B(n_984),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_958),
.B(n_968),
.Y(n_1137)
);

INVx4_ASAP7_75t_SL g1138 ( 
.A(n_1063),
.Y(n_1138)
);

INVx3_ASAP7_75t_SL g1139 ( 
.A(n_1063),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1068),
.A2(n_946),
.B(n_953),
.Y(n_1140)
);

BUFx4_ASAP7_75t_SL g1141 ( 
.A(n_1057),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_SL g1142 ( 
.A1(n_992),
.A2(n_967),
.B(n_988),
.C(n_989),
.Y(n_1142)
);

AO31x2_ASAP7_75t_L g1143 ( 
.A1(n_977),
.A2(n_999),
.A3(n_991),
.B(n_987),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1035),
.A2(n_985),
.B(n_1028),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1032),
.B(n_979),
.Y(n_1145)
);

HB1xp67_ASAP7_75t_L g1146 ( 
.A(n_1032),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_964),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_947),
.A2(n_955),
.B1(n_972),
.B2(n_976),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1070),
.A2(n_962),
.B(n_1043),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_946),
.A2(n_953),
.B(n_1057),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1055),
.Y(n_1151)
);

OAI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1084),
.A2(n_1009),
.B1(n_1050),
.B2(n_1039),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1061),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_966),
.B(n_970),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_969),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_946),
.A2(n_953),
.B(n_1057),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_964),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1030),
.B(n_946),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1071),
.A2(n_953),
.B(n_1080),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1048),
.B(n_1064),
.Y(n_1160)
);

AO32x2_ASAP7_75t_L g1161 ( 
.A1(n_949),
.A2(n_960),
.A3(n_962),
.B1(n_1071),
.B2(n_1061),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1071),
.A2(n_1025),
.B(n_1048),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1025),
.A2(n_1061),
.B(n_1064),
.C(n_949),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_960),
.B(n_1061),
.Y(n_1164)
);

INVx2_ASAP7_75t_SL g1165 ( 
.A(n_1064),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1064),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_983),
.A2(n_549),
.B(n_542),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1081),
.B(n_603),
.Y(n_1168)
);

INVxp67_ASAP7_75t_L g1169 ( 
.A(n_973),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1029),
.A2(n_1062),
.A3(n_1079),
.B(n_1054),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_996),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1081),
.A2(n_1014),
.B(n_1006),
.Y(n_1175)
);

OAI22x1_ASAP7_75t_L g1176 ( 
.A1(n_978),
.A2(n_603),
.B1(n_993),
.B2(n_905),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_981),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1019),
.Y(n_1178)
);

OR2x6_ASAP7_75t_L g1179 ( 
.A(n_1057),
.B(n_940),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_1005),
.B(n_731),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1019),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1081),
.B(n_477),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1081),
.B(n_477),
.Y(n_1184)
);

NAND3xp33_ASAP7_75t_L g1185 ( 
.A(n_1081),
.B(n_603),
.C(n_634),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1054),
.A2(n_1062),
.B(n_1000),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1061),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1081),
.B(n_603),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1019),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_981),
.Y(n_1191)
);

INVx3_ASAP7_75t_L g1192 ( 
.A(n_1061),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_1081),
.A2(n_948),
.B(n_978),
.C(n_1014),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1081),
.B(n_477),
.Y(n_1195)
);

AOI21x1_ASAP7_75t_SL g1196 ( 
.A1(n_1082),
.A2(n_1085),
.B(n_601),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1019),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_SL g1198 ( 
.A(n_950),
.B(n_522),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1081),
.A2(n_1014),
.B(n_1006),
.Y(n_1200)
);

AO31x2_ASAP7_75t_L g1201 ( 
.A1(n_1029),
.A2(n_1062),
.A3(n_1079),
.B(n_1054),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_1081),
.B(n_603),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1204)
);

AO32x2_ASAP7_75t_L g1205 ( 
.A1(n_1037),
.A2(n_997),
.A3(n_660),
.B1(n_995),
.B2(n_1038),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1207)
);

AO21x2_ASAP7_75t_L g1208 ( 
.A1(n_1000),
.A2(n_1029),
.B(n_1081),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1086),
.B(n_623),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1081),
.B(n_477),
.Y(n_1210)
);

NOR2xp33_ASAP7_75t_L g1211 ( 
.A(n_1081),
.B(n_603),
.Y(n_1211)
);

AOI221x1_ASAP7_75t_L g1212 ( 
.A1(n_1081),
.A2(n_1040),
.B1(n_1047),
.B2(n_997),
.C(n_603),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1081),
.A2(n_1014),
.B(n_1006),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1019),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1218)
);

OAI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1081),
.A2(n_1014),
.B(n_1006),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_973),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1000),
.A2(n_549),
.B(n_542),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_998),
.A2(n_1073),
.B(n_1018),
.Y(n_1223)
);

BUFx2_ASAP7_75t_R g1224 ( 
.A(n_1005),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1081),
.A2(n_1014),
.B(n_1006),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_1083),
.Y(n_1226)
);

AND2x2_ASAP7_75t_SL g1227 ( 
.A(n_979),
.B(n_1088),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_973),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1019),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1081),
.B(n_477),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1081),
.B(n_477),
.Y(n_1231)
);

OAI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1168),
.A2(n_1211),
.B1(n_1202),
.B2(n_1189),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1137),
.Y(n_1233)
);

HB1xp67_ASAP7_75t_L g1234 ( 
.A(n_1112),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1132),
.Y(n_1235)
);

CKINVDCx20_ASAP7_75t_R g1236 ( 
.A(n_1226),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1227),
.A2(n_1185),
.B1(n_1097),
.B2(n_1198),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1097),
.A2(n_1108),
.B1(n_1230),
.B2(n_1195),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1198),
.A2(n_1231),
.B1(n_1230),
.B2(n_1183),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1095),
.B(n_1209),
.Y(n_1240)
);

BUFx8_ASAP7_75t_SL g1241 ( 
.A(n_1173),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1091),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1098),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1183),
.A2(n_1231),
.B1(n_1195),
.B2(n_1184),
.Y(n_1244)
);

BUFx2_ASAP7_75t_L g1245 ( 
.A(n_1125),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1116),
.A2(n_1145),
.B1(n_1184),
.B2(n_1210),
.Y(n_1246)
);

INVx6_ASAP7_75t_L g1247 ( 
.A(n_1138),
.Y(n_1247)
);

BUFx12f_ASAP7_75t_L g1248 ( 
.A(n_1115),
.Y(n_1248)
);

BUFx10_ASAP7_75t_L g1249 ( 
.A(n_1130),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1210),
.A2(n_1116),
.B1(n_1176),
.B2(n_1219),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1100),
.Y(n_1251)
);

AO22x1_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1139),
.B1(n_1119),
.B2(n_1134),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1112),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1220),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1147),
.Y(n_1255)
);

INVx2_ASAP7_75t_SL g1256 ( 
.A(n_1101),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1120),
.B(n_1228),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1224),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1175),
.A2(n_1214),
.B1(n_1225),
.B2(n_1219),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1105),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1118),
.B(n_1146),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1175),
.A2(n_1214),
.B1(n_1200),
.B2(n_1225),
.Y(n_1262)
);

BUFx2_ASAP7_75t_L g1263 ( 
.A(n_1169),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1128),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1102),
.B1(n_1120),
.B2(n_1133),
.Y(n_1265)
);

BUFx6f_ASAP7_75t_L g1266 ( 
.A(n_1129),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1129),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1178),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1181),
.Y(n_1269)
);

INVx3_ASAP7_75t_SL g1270 ( 
.A(n_1138),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1200),
.A2(n_1186),
.B1(n_1093),
.B2(n_1149),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1159),
.B(n_1148),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1138),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1135),
.A2(n_1123),
.B1(n_1114),
.B2(n_1217),
.Y(n_1274)
);

BUFx2_ASAP7_75t_SL g1275 ( 
.A(n_1180),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1190),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1133),
.A2(n_1194),
.B1(n_1123),
.B2(n_1179),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1129),
.Y(n_1278)
);

BUFx10_ASAP7_75t_L g1279 ( 
.A(n_1179),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1179),
.A2(n_1135),
.B1(n_1142),
.B2(n_1122),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1197),
.Y(n_1281)
);

BUFx4_ASAP7_75t_SL g1282 ( 
.A(n_1166),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1147),
.Y(n_1283)
);

BUFx10_ASAP7_75t_L g1284 ( 
.A(n_1164),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1157),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1141),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1122),
.A2(n_1126),
.B1(n_1131),
.B2(n_1151),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1177),
.B(n_1191),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1157),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_1224),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1107),
.A2(n_1099),
.B1(n_1208),
.B2(n_1093),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1153),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1229),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1208),
.A2(n_1149),
.B1(n_1186),
.B2(n_1124),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1188),
.Y(n_1295)
);

OAI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1212),
.A2(n_1158),
.B1(n_1121),
.B2(n_1089),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_1188),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1159),
.B(n_1192),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1154),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1155),
.Y(n_1300)
);

INVx5_ASAP7_75t_L g1301 ( 
.A(n_1192),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1158),
.A2(n_1089),
.B1(n_1094),
.B2(n_1109),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1152),
.A2(n_1090),
.B1(n_1092),
.B2(n_1205),
.Y(n_1303)
);

INVx8_ASAP7_75t_L g1304 ( 
.A(n_1163),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1154),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1165),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1160),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1160),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1162),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1143),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1140),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1167),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1170),
.A2(n_1222),
.B(n_1216),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1143),
.Y(n_1314)
);

BUFx12f_ASAP7_75t_L g1315 ( 
.A(n_1196),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1113),
.A2(n_1150),
.B1(n_1156),
.B2(n_1090),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1144),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1103),
.B(n_1171),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1161),
.Y(n_1319)
);

AOI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1127),
.A2(n_1110),
.B1(n_1106),
.B2(n_1218),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1161),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1090),
.A2(n_1205),
.B1(n_1161),
.B2(n_1106),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1205),
.A2(n_1111),
.B1(n_1223),
.B2(n_1199),
.Y(n_1323)
);

INVx6_ASAP7_75t_L g1324 ( 
.A(n_1136),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1172),
.A2(n_1221),
.B1(n_1204),
.B2(n_1207),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1171),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1187),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1096),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1201),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1174),
.A2(n_1182),
.B1(n_1136),
.B2(n_1193),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1203),
.B(n_1206),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1201),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1213),
.A2(n_1215),
.B1(n_1103),
.B2(n_1096),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1096),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1103),
.A2(n_603),
.B1(n_1189),
.B2(n_1168),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1137),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1227),
.A2(n_1097),
.B1(n_603),
.B2(n_1211),
.Y(n_1337)
);

CKINVDCx11_ASAP7_75t_R g1338 ( 
.A(n_1132),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1137),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1137),
.Y(n_1341)
);

INVx4_ASAP7_75t_L g1342 ( 
.A(n_1138),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1138),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1129),
.Y(n_1344)
);

INVx6_ASAP7_75t_L g1345 ( 
.A(n_1138),
.Y(n_1345)
);

CKINVDCx11_ASAP7_75t_R g1346 ( 
.A(n_1132),
.Y(n_1346)
);

INVx6_ASAP7_75t_L g1347 ( 
.A(n_1138),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1168),
.A2(n_603),
.B(n_1081),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1168),
.A2(n_1189),
.B1(n_1211),
.B2(n_1202),
.Y(n_1349)
);

OR2x2_ASAP7_75t_L g1350 ( 
.A(n_1318),
.B(n_1326),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1334),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1349),
.B(n_1262),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1329),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1332),
.Y(n_1354)
);

INVxp67_ASAP7_75t_L g1355 ( 
.A(n_1245),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1235),
.Y(n_1356)
);

OR2x6_ASAP7_75t_L g1357 ( 
.A(n_1272),
.B(n_1324),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1318),
.B(n_1319),
.Y(n_1358)
);

OAI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1337),
.A2(n_1259),
.B1(n_1262),
.B2(n_1349),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1232),
.A2(n_1238),
.B1(n_1337),
.B2(n_1274),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1310),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1314),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1328),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_L g1364 ( 
.A(n_1240),
.B(n_1299),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_1234),
.Y(n_1365)
);

AO21x2_ASAP7_75t_L g1366 ( 
.A1(n_1296),
.A2(n_1333),
.B(n_1313),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1317),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1238),
.A2(n_1274),
.B1(n_1316),
.B2(n_1322),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1234),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1321),
.B(n_1259),
.Y(n_1370)
);

NOR2x1_ASAP7_75t_L g1371 ( 
.A(n_1348),
.B(n_1311),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1322),
.Y(n_1372)
);

BUFx6f_ASAP7_75t_L g1373 ( 
.A(n_1298),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1287),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1257),
.B(n_1250),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1279),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1320),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1242),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1243),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1305),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1331),
.A2(n_1330),
.B(n_1325),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1251),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1260),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1264),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1250),
.B(n_1237),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1268),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1237),
.B(n_1307),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1296),
.A2(n_1333),
.B(n_1302),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1269),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1276),
.Y(n_1390)
);

BUFx3_ASAP7_75t_L g1391 ( 
.A(n_1279),
.Y(n_1391)
);

NAND2x1p5_ASAP7_75t_L g1392 ( 
.A(n_1280),
.B(n_1309),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1253),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1302),
.A2(n_1335),
.B(n_1277),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1272),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1308),
.B(n_1271),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1261),
.B(n_1241),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1281),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1239),
.B(n_1244),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1293),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1331),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1233),
.Y(n_1402)
);

CKINVDCx14_ASAP7_75t_R g1403 ( 
.A(n_1338),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1294),
.A2(n_1291),
.B(n_1323),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1330),
.A2(n_1325),
.B(n_1323),
.Y(n_1405)
);

CKINVDCx8_ASAP7_75t_R g1406 ( 
.A(n_1275),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1346),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1315),
.Y(n_1408)
);

INVx3_ASAP7_75t_SL g1409 ( 
.A(n_1270),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1291),
.A2(n_1294),
.B(n_1244),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1284),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1239),
.A2(n_1303),
.B(n_1265),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1336),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1246),
.B(n_1303),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1339),
.A2(n_1340),
.B(n_1341),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1327),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1273),
.B(n_1342),
.Y(n_1417)
);

INVx1_ASAP7_75t_SL g1418 ( 
.A(n_1254),
.Y(n_1418)
);

INVx5_ASAP7_75t_L g1419 ( 
.A(n_1304),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1246),
.B(n_1288),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1304),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1301),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1295),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1292),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1312),
.A2(n_1300),
.B1(n_1263),
.B2(n_1286),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1273),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1255),
.A2(n_1252),
.B(n_1282),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1297),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1342),
.A2(n_1266),
.B(n_1344),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1365),
.B(n_1284),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1369),
.B(n_1256),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1396),
.B(n_1267),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1396),
.B(n_1267),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1405),
.A2(n_1290),
.B(n_1258),
.Y(n_1434)
);

INVx4_ASAP7_75t_L g1435 ( 
.A(n_1419),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1372),
.B(n_1266),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1409),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1375),
.B(n_1306),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1372),
.B(n_1267),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1357),
.B(n_1347),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1370),
.B(n_1266),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1378),
.Y(n_1442)
);

A2O1A1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1360),
.A2(n_1270),
.B(n_1247),
.C(n_1345),
.Y(n_1443)
);

NOR2xp33_ASAP7_75t_L g1444 ( 
.A(n_1416),
.B(n_1249),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1420),
.B(n_1423),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1370),
.B(n_1388),
.Y(n_1446)
);

AOI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1388),
.A2(n_1289),
.B(n_1278),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1378),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1388),
.B(n_1249),
.Y(n_1449)
);

OAI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1360),
.A2(n_1283),
.B(n_1236),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1388),
.B(n_1285),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1358),
.B(n_1285),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1359),
.B(n_1289),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_SL g1454 ( 
.A1(n_1359),
.A2(n_1247),
.B(n_1343),
.Y(n_1454)
);

AOI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1352),
.A2(n_1248),
.B1(n_1343),
.B2(n_1345),
.Y(n_1455)
);

NAND4xp25_ASAP7_75t_L g1456 ( 
.A(n_1368),
.B(n_1343),
.C(n_1345),
.D(n_1347),
.Y(n_1456)
);

AOI221xp5_ASAP7_75t_L g1457 ( 
.A1(n_1352),
.A2(n_1374),
.B1(n_1368),
.B2(n_1414),
.C(n_1385),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1390),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1379),
.B(n_1382),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1416),
.A2(n_1385),
.B1(n_1406),
.B2(n_1425),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1416),
.A2(n_1406),
.B1(n_1418),
.B2(n_1371),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1367),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1371),
.A2(n_1412),
.B(n_1399),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1390),
.Y(n_1464)
);

NAND2xp33_ASAP7_75t_R g1465 ( 
.A(n_1416),
.B(n_1426),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1382),
.B(n_1383),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

AO32x1_ASAP7_75t_L g1468 ( 
.A1(n_1353),
.A2(n_1354),
.A3(n_1351),
.B1(n_1362),
.B2(n_1361),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1412),
.A2(n_1399),
.B(n_1414),
.C(n_1410),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1398),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1364),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_L g1473 ( 
.A1(n_1374),
.A2(n_1392),
.B(n_1355),
.C(n_1418),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1383),
.B(n_1384),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1366),
.A2(n_1357),
.B(n_1394),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1412),
.A2(n_1392),
.B(n_1410),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1387),
.B(n_1400),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1387),
.B(n_1400),
.Y(n_1478)
);

AOI21xp33_ASAP7_75t_L g1479 ( 
.A1(n_1394),
.A2(n_1395),
.B(n_1392),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1405),
.A2(n_1410),
.B(n_1381),
.Y(n_1480)
);

O2A1O1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1395),
.A2(n_1409),
.B(n_1394),
.C(n_1428),
.Y(n_1481)
);

NOR2x1_ASAP7_75t_SL g1482 ( 
.A(n_1357),
.B(n_1415),
.Y(n_1482)
);

OA21x2_ASAP7_75t_L g1483 ( 
.A1(n_1381),
.A2(n_1377),
.B(n_1361),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1427),
.B(n_1373),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1427),
.A2(n_1429),
.B(n_1401),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1386),
.B(n_1389),
.Y(n_1486)
);

AO21x1_ASAP7_75t_L g1487 ( 
.A1(n_1421),
.A2(n_1428),
.B(n_1413),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1457),
.A2(n_1394),
.B1(n_1420),
.B2(n_1408),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1442),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1448),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1445),
.B(n_1377),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1432),
.B(n_1404),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1464),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1470),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1477),
.B(n_1415),
.Y(n_1497)
);

NAND2x1p5_ASAP7_75t_SL g1498 ( 
.A(n_1449),
.B(n_1401),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1446),
.B(n_1366),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1432),
.B(n_1404),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1446),
.B(n_1366),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1437),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1459),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1459),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1466),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1462),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1466),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1441),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1366),
.Y(n_1509)
);

NOR2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1456),
.B(n_1437),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1440),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_L g1512 ( 
.A(n_1449),
.B(n_1415),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1471),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1433),
.B(n_1404),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1454),
.A2(n_1408),
.B1(n_1373),
.B2(n_1411),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1474),
.B(n_1380),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1469),
.B(n_1350),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1433),
.B(n_1404),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1451),
.B(n_1404),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1451),
.B(n_1363),
.Y(n_1520)
);

OAI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1443),
.A2(n_1406),
.B1(n_1403),
.B2(n_1413),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1486),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1469),
.B(n_1476),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1468),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1443),
.A2(n_1419),
.B1(n_1380),
.B2(n_1409),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1463),
.B(n_1402),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_L g1527 ( 
.A1(n_1488),
.A2(n_1473),
.B1(n_1481),
.B2(n_1467),
.C(n_1475),
.Y(n_1527)
);

AOI221xp5_ASAP7_75t_L g1528 ( 
.A1(n_1523),
.A2(n_1450),
.B1(n_1479),
.B2(n_1460),
.C(n_1461),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1523),
.B(n_1485),
.C(n_1453),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1526),
.B(n_1441),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1494),
.B(n_1484),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1526),
.B(n_1430),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1508),
.B(n_1452),
.Y(n_1533)
);

NAND2xp67_ASAP7_75t_L g1534 ( 
.A(n_1519),
.B(n_1424),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1489),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1436),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1490),
.Y(n_1537)
);

NAND3xp33_ASAP7_75t_L g1538 ( 
.A(n_1512),
.B(n_1453),
.C(n_1447),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1517),
.B(n_1483),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1516),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1517),
.B(n_1434),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1542)
);

INVxp67_ASAP7_75t_SL g1543 ( 
.A(n_1512),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_SL g1544 ( 
.A1(n_1521),
.A2(n_1525),
.B1(n_1444),
.B2(n_1511),
.Y(n_1544)
);

NOR2xp67_ASAP7_75t_L g1545 ( 
.A(n_1497),
.B(n_1435),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1434),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1489),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1514),
.B(n_1434),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1493),
.B(n_1436),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1522),
.B(n_1439),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1435),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1491),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1521),
.A2(n_1472),
.B1(n_1440),
.B2(n_1438),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1509),
.B(n_1480),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1516),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1499),
.B(n_1480),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1520),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1511),
.B(n_1502),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1511),
.B(n_1440),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1506),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1525),
.A2(n_1440),
.B(n_1482),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1491),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1502),
.B(n_1435),
.Y(n_1565)
);

HB1xp67_ASAP7_75t_L g1566 ( 
.A(n_1520),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1549),
.B(n_1519),
.Y(n_1567)
);

AND2x4_ASAP7_75t_L g1568 ( 
.A(n_1552),
.B(n_1506),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1549),
.B(n_1514),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1531),
.B(n_1518),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1531),
.B(n_1518),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1539),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1552),
.B(n_1506),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1538),
.B(n_1499),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1535),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1497),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1542),
.B(n_1503),
.Y(n_1577)
);

NOR2xp33_ASAP7_75t_L g1578 ( 
.A(n_1532),
.B(n_1431),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1579)
);

INVxp67_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1546),
.B(n_1504),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1539),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1535),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1548),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1530),
.B(n_1504),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1546),
.B(n_1505),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1543),
.B(n_1505),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1544),
.Y(n_1588)
);

INVx2_ASAP7_75t_SL g1589 ( 
.A(n_1561),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1548),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1555),
.B(n_1498),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1555),
.B(n_1498),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1541),
.B(n_1507),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1553),
.Y(n_1594)
);

INVx3_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

NOR2xp67_ASAP7_75t_L g1596 ( 
.A(n_1541),
.B(n_1501),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1537),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1563),
.Y(n_1598)
);

OAI33xp33_ASAP7_75t_L g1599 ( 
.A1(n_1547),
.A2(n_1524),
.A3(n_1501),
.B1(n_1496),
.B2(n_1495),
.B3(n_1492),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1580),
.B(n_1527),
.Y(n_1600)
);

NAND4xp25_ASAP7_75t_L g1601 ( 
.A(n_1580),
.B(n_1528),
.C(n_1544),
.D(n_1554),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1568),
.B(n_1559),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1585),
.B(n_1533),
.Y(n_1604)
);

OR2x6_ASAP7_75t_L g1605 ( 
.A(n_1574),
.B(n_1562),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1568),
.B(n_1573),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1574),
.Y(n_1607)
);

NAND2x1_ASAP7_75t_L g1608 ( 
.A(n_1568),
.B(n_1559),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1534),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1568),
.B(n_1559),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1565),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1585),
.B(n_1536),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1573),
.B(n_1565),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1576),
.B(n_1550),
.Y(n_1614)
);

INVx1_ASAP7_75t_SL g1615 ( 
.A(n_1588),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1573),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

OR2x2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.B(n_1547),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1575),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_SL g1620 ( 
.A1(n_1588),
.A2(n_1534),
.B1(n_1564),
.B2(n_1557),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1551),
.Y(n_1621)
);

AOI32xp33_ASAP7_75t_L g1622 ( 
.A1(n_1570),
.A2(n_1565),
.A3(n_1552),
.B1(n_1515),
.B2(n_1524),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1545),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1597),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1575),
.Y(n_1626)
);

INVxp67_ASAP7_75t_SL g1627 ( 
.A(n_1596),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1573),
.B(n_1561),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1579),
.B(n_1545),
.Y(n_1629)
);

INVxp67_ASAP7_75t_L g1630 ( 
.A(n_1587),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1590),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1590),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1572),
.B(n_1557),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1570),
.B(n_1566),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1572),
.B(n_1498),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1590),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1570),
.B(n_1571),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1572),
.B(n_1563),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1571),
.B(n_1558),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1577),
.B(n_1513),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1615),
.B(n_1407),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1606),
.B(n_1571),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1614),
.B(n_1572),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1600),
.B(n_1356),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1619),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1647)
);

INVx1_ASAP7_75t_SL g1648 ( 
.A(n_1602),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1630),
.B(n_1582),
.Y(n_1649)
);

NAND2xp33_ASAP7_75t_L g1650 ( 
.A(n_1622),
.B(n_1510),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1601),
.B(n_1577),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1617),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1621),
.B(n_1581),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1629),
.B(n_1581),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1638),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1623),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1625),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1606),
.B(n_1569),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1612),
.B(n_1582),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1625),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1662)
);

NOR2xp67_ASAP7_75t_L g1663 ( 
.A(n_1616),
.B(n_1591),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1626),
.Y(n_1664)
);

OAI32xp33_ASAP7_75t_L g1665 ( 
.A1(n_1636),
.A2(n_1591),
.A3(n_1592),
.B1(n_1582),
.B2(n_1465),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1603),
.B(n_1569),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1605),
.A2(n_1620),
.B(n_1627),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1631),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1608),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1634),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1604),
.B(n_1586),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_SL g1672 ( 
.A(n_1605),
.B(n_1408),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1618),
.B(n_1582),
.Y(n_1673)
);

NOR2xp67_ASAP7_75t_SL g1674 ( 
.A(n_1616),
.B(n_1408),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1633),
.B(n_1591),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1635),
.B(n_1586),
.Y(n_1676)
);

OAI322xp33_ASAP7_75t_L g1677 ( 
.A1(n_1651),
.A2(n_1636),
.A3(n_1592),
.B1(n_1633),
.B2(n_1637),
.C1(n_1632),
.C2(n_1639),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1642),
.B(n_1610),
.Y(n_1678)
);

XOR2xp5_ASAP7_75t_L g1679 ( 
.A(n_1667),
.B(n_1455),
.Y(n_1679)
);

NAND2xp33_ASAP7_75t_L g1680 ( 
.A(n_1669),
.B(n_1510),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1610),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1646),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1650),
.A2(n_1605),
.B1(n_1624),
.B2(n_1611),
.Y(n_1683)
);

XOR2x2_ASAP7_75t_L g1684 ( 
.A(n_1645),
.B(n_1397),
.Y(n_1684)
);

AOI32xp33_ASAP7_75t_L g1685 ( 
.A1(n_1672),
.A2(n_1648),
.A3(n_1656),
.B1(n_1643),
.B2(n_1669),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1646),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1648),
.B(n_1635),
.Y(n_1687)
);

INVx1_ASAP7_75t_SL g1688 ( 
.A(n_1653),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1665),
.A2(n_1656),
.B1(n_1672),
.B2(n_1652),
.C(n_1647),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1657),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1665),
.A2(n_1605),
.B(n_1599),
.Y(n_1691)
);

AOI21xp33_ASAP7_75t_L g1692 ( 
.A1(n_1657),
.A2(n_1592),
.B(n_1639),
.Y(n_1692)
);

OR2x6_ASAP7_75t_L g1693 ( 
.A(n_1663),
.B(n_1408),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1663),
.A2(n_1599),
.B(n_1624),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1640),
.Y(n_1695)
);

OAI31xp33_ASAP7_75t_L g1696 ( 
.A1(n_1655),
.A2(n_1624),
.A3(n_1611),
.B(n_1613),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1662),
.Y(n_1697)
);

AOI22xp33_ASAP7_75t_L g1698 ( 
.A1(n_1671),
.A2(n_1613),
.B1(n_1560),
.B2(n_1628),
.Y(n_1698)
);

INVx2_ASAP7_75t_SL g1699 ( 
.A(n_1666),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1674),
.A2(n_1596),
.B(n_1640),
.C(n_1628),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1674),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_SL g1702 ( 
.A1(n_1691),
.A2(n_1649),
.B(n_1668),
.C(n_1664),
.Y(n_1702)
);

INVxp67_ASAP7_75t_L g1703 ( 
.A(n_1688),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1688),
.B(n_1666),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1699),
.B(n_1659),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1685),
.A2(n_1689),
.B(n_1683),
.C(n_1696),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1682),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1693),
.Y(n_1708)
);

AOI222xp33_ASAP7_75t_L g1709 ( 
.A1(n_1687),
.A2(n_1664),
.B1(n_1668),
.B2(n_1676),
.C1(n_1659),
.C2(n_1654),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1687),
.B(n_1644),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1693),
.Y(n_1711)
);

NAND2xp33_ASAP7_75t_SL g1712 ( 
.A(n_1678),
.B(n_1675),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1690),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1681),
.B(n_1567),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_SL g1716 ( 
.A1(n_1679),
.A2(n_1675),
.B(n_1644),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1677),
.A2(n_1660),
.B1(n_1649),
.B2(n_1673),
.C(n_1661),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1697),
.B(n_1660),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1695),
.Y(n_1719)
);

INVxp67_ASAP7_75t_L g1720 ( 
.A(n_1693),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1703),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1703),
.B(n_1694),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1704),
.Y(n_1723)
);

XNOR2x1_ASAP7_75t_L g1724 ( 
.A(n_1719),
.B(n_1684),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1716),
.B(n_1701),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1715),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1712),
.Y(n_1727)
);

INVxp67_ASAP7_75t_SL g1728 ( 
.A(n_1720),
.Y(n_1728)
);

INVx1_ASAP7_75t_SL g1729 ( 
.A(n_1712),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1706),
.B(n_1680),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1702),
.A2(n_1700),
.B(n_1698),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1727),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1729),
.B(n_1717),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1728),
.B(n_1709),
.Y(n_1734)
);

OAI321xp33_ASAP7_75t_L g1735 ( 
.A1(n_1731),
.A2(n_1718),
.A3(n_1720),
.B1(n_1710),
.B2(n_1711),
.C(n_1705),
.Y(n_1735)
);

AOI21xp33_ASAP7_75t_SL g1736 ( 
.A1(n_1724),
.A2(n_1708),
.B(n_1713),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_SL g1737 ( 
.A(n_1721),
.B(n_1692),
.Y(n_1737)
);

NAND2x1p5_ASAP7_75t_L g1738 ( 
.A(n_1730),
.B(n_1707),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1726),
.B(n_1714),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_1692),
.C(n_1658),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1728),
.Y(n_1741)
);

OAI21xp33_ASAP7_75t_L g1742 ( 
.A1(n_1725),
.A2(n_1673),
.B(n_1670),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1733),
.B(n_1723),
.C(n_1670),
.D(n_1661),
.Y(n_1743)
);

OAI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1723),
.B(n_1658),
.C(n_1411),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1735),
.A2(n_1634),
.B1(n_1587),
.B2(n_1589),
.C(n_1594),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1737),
.A2(n_1589),
.B(n_1597),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1741),
.Y(n_1747)
);

OAI211xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1742),
.A2(n_1732),
.B(n_1740),
.C(n_1736),
.Y(n_1748)
);

AOI221xp5_ASAP7_75t_L g1749 ( 
.A1(n_1748),
.A2(n_1738),
.B1(n_1739),
.B2(n_1589),
.C(n_1587),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1743),
.A2(n_1738),
.B1(n_1594),
.B2(n_1411),
.C(n_1595),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1744),
.A2(n_1408),
.B(n_1427),
.C(n_1417),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1747),
.B(n_1376),
.C(n_1391),
.Y(n_1752)
);

AOI211xp5_ASAP7_75t_L g1753 ( 
.A1(n_1746),
.A2(n_1417),
.B(n_1391),
.C(n_1376),
.Y(n_1753)
);

OAI22x1_ASAP7_75t_L g1754 ( 
.A1(n_1745),
.A2(n_1595),
.B1(n_1594),
.B2(n_1597),
.Y(n_1754)
);

NAND4xp75_ASAP7_75t_L g1755 ( 
.A(n_1749),
.B(n_1750),
.C(n_1751),
.D(n_1752),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1753),
.B(n_1595),
.Y(n_1756)
);

XNOR2xp5_ASAP7_75t_L g1757 ( 
.A(n_1754),
.B(n_1376),
.Y(n_1757)
);

NAND4xp75_ASAP7_75t_L g1758 ( 
.A(n_1749),
.B(n_1429),
.C(n_1487),
.D(n_1593),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1754),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1759),
.B(n_1595),
.Y(n_1760)
);

HB1xp67_ASAP7_75t_L g1761 ( 
.A(n_1757),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1755),
.B(n_1595),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1762),
.A2(n_1756),
.B1(n_1758),
.B2(n_1593),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1763),
.Y(n_1764)
);

INVx6_ASAP7_75t_L g1765 ( 
.A(n_1764),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1760),
.B1(n_1761),
.B2(n_1593),
.Y(n_1766)
);

XNOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1766),
.B(n_1417),
.Y(n_1767)
);

OAI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1765),
.A2(n_1598),
.B1(n_1584),
.B2(n_1641),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1767),
.B(n_1567),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

XNOR2xp5_ASAP7_75t_L g1771 ( 
.A(n_1770),
.B(n_1417),
.Y(n_1771)
);

OAI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1769),
.B(n_1567),
.Y(n_1772)
);

INVx6_ASAP7_75t_L g1773 ( 
.A(n_1772),
.Y(n_1773)
);

OAI221xp5_ASAP7_75t_R g1774 ( 
.A1(n_1773),
.A2(n_1465),
.B1(n_1598),
.B2(n_1584),
.C(n_1391),
.Y(n_1774)
);

AOI211xp5_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1421),
.B(n_1426),
.C(n_1422),
.Y(n_1775)
);


endmodule