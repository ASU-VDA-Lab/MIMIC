module real_jpeg_12810_n_17 (n_5, n_4, n_8, n_0, n_12, n_310, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_310;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g82 ( 
.A(n_0),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_3),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_4),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_4),
.B(n_56),
.C(n_60),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_4),
.B(n_45),
.Y(n_131)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_4),
.A2(n_138),
.B(n_141),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_30),
.B(n_44),
.C(n_169),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_123),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_4),
.B(n_25),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_5),
.A2(n_35),
.B1(n_56),
.B2(n_57),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_5),
.A2(n_35),
.B1(n_46),
.B2(n_47),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_9),
.A2(n_56),
.B1(n_57),
.B2(n_135),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_9),
.A2(n_30),
.B1(n_31),
.B2(n_135),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_135),
.Y(n_242)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_11),
.A2(n_56),
.B1(n_57),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_140),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_140),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_140),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_12),
.B(n_31),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_13),
.A2(n_27),
.B1(n_56),
.B2(n_57),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_13),
.A2(n_27),
.B1(n_46),
.B2(n_47),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_13),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_94),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_14),
.A2(n_30),
.B1(n_31),
.B2(n_94),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_15),
.A2(n_40),
.B1(n_46),
.B2(n_47),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_40),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_15),
.A2(n_40),
.B1(n_56),
.B2(n_57),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_16),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_16),
.A2(n_56),
.B1(n_57),
.B2(n_65),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_95),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_20),
.B(n_95),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_68),
.C(n_76),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_21),
.B(n_68),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_36),
.B2(n_67),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_22),
.A2(n_23),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_37),
.C(n_53),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_29),
.B2(n_34),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_24),
.A2(n_29),
.B(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_26),
.A2(n_28),
.B(n_123),
.C(n_214),
.Y(n_213)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_26),
.A2(n_30),
.A3(n_32),
.B1(n_215),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_28),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_28),
.A2(n_29),
.B1(n_34),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_28),
.A2(n_29),
.B1(n_242),
.B2(n_262),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_28),
.A2(n_262),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_33),
.Y(n_28)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_29),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_29),
.B(n_93),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_29),
.A2(n_90),
.B(n_242),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_52),
.B1(n_53),
.B2(n_66),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_37),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_45),
.B2(n_49),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_41),
.B(n_176),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_43),
.A2(n_46),
.B(n_123),
.Y(n_169)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_45),
.B(n_176),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_46),
.A2(n_47),
.B1(n_59),
.B2(n_60),
.Y(n_62)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_47),
.B(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_50),
.A2(n_70),
.B1(n_72),
.B2(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_53),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_61),
.B(n_63),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_61),
.B1(n_87),
.B2(n_88),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_54),
.B(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_54),
.A2(n_61),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_54),
.A2(n_61),
.B1(n_221),
.B2(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_54),
.A2(n_61),
.B1(n_87),
.B2(n_249),
.Y(n_255)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_64),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_134),
.B(n_136),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_55),
.B(n_123),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_55),
.A2(n_136),
.B(n_220),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_57),
.B(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_61),
.B(n_125),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_68),
.A2(n_69),
.B(n_73),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_70),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_70),
.A2(n_72),
.B1(n_189),
.B2(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_70),
.A2(n_175),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_264),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_72),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_72),
.A2(n_190),
.B(n_264),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_74),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_74),
.A2(n_124),
.B(n_202),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_76),
.B(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_80),
.B(n_89),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_77),
.A2(n_78),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_79),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_81),
.A2(n_82),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_81),
.B(n_142),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_81),
.A2(n_82),
.B1(n_232),
.B2(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_82),
.B(n_142),
.Y(n_141)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_84),
.A2(n_138),
.B1(n_155),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_89),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_304),
.B(n_308),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_291),
.B(n_303),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_274),
.B(n_290),
.Y(n_112)
);

OAI321xp33_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_234),
.A3(n_267),
.B1(n_272),
.B2(n_273),
.C(n_310),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_206),
.B(n_233),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_183),
.B(n_205),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_164),
.B(n_182),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_143),
.B(n_163),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_128),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_119),
.B(n_128),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_126),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_121),
.B1(n_126),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_133),
.C(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_138),
.A2(n_155),
.B1(n_171),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_138),
.A2(n_155),
.B1(n_197),
.B2(n_231),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_151),
.B(n_162),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_145),
.B(n_149),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_157),
.B(n_161),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_154),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_155),
.A2(n_156),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_165),
.B(n_166),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_177),
.C(n_181),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_170),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_177),
.B1(n_180),
.B2(n_181),
.Y(n_172)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_173),
.Y(n_181)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_179),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_198),
.B2(n_199),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_201),
.C(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_192),
.C(n_196),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_196),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_201),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_208),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_223),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_209),
.B(n_224),
.C(n_225),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_216),
.B2(n_222),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_217),
.C(n_219),
.Y(n_250)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_230),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_251),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_251),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.C(n_250),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_237),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_244),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_250),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_248),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_266),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_259),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_259),
.C(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_257),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_263),
.C(n_265),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_268),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_289),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_275),
.B(n_289),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_280),
.B2(n_281),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_287),
.B2(n_288),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_285),
.C(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_293),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_302),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_296),
.B(n_297),
.C(n_302),
.Y(n_307)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_305),
.B(n_307),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_307),
.Y(n_308)
);


endmodule