module fake_jpeg_28330_n_204 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

CKINVDCx6p67_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_56),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_47),
.B(n_35),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_23),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_21),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_53),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_34),
.Y(n_53)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_55),
.B(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_20),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_64),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_33),
.B1(n_27),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_29),
.B1(n_27),
.B2(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_87),
.Y(n_104)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_33),
.B1(n_40),
.B2(n_43),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_33),
.B1(n_43),
.B2(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_79),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_43),
.B(n_35),
.C(n_36),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_71),
.A2(n_84),
.B(n_38),
.C(n_32),
.Y(n_119)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_37),
.B1(n_44),
.B2(n_28),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_44),
.B1(n_20),
.B2(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_31),
.B1(n_27),
.B2(n_29),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_83),
.Y(n_97)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_28),
.B1(n_18),
.B2(n_22),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_80),
.Y(n_106)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_54),
.A2(n_28),
.B1(n_22),
.B2(n_19),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_30),
.B1(n_20),
.B2(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_86),
.B(n_90),
.Y(n_117)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_95),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_89),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

CKINVDCx12_ASAP7_75t_R g95 ( 
.A(n_54),
.Y(n_95)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_75),
.B(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_81),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_55),
.B1(n_57),
.B2(n_60),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_103),
.A2(n_105),
.B1(n_119),
.B2(n_88),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_50),
.C(n_51),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_38),
.C(n_88),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_29),
.A3(n_30),
.B1(n_19),
.B2(n_20),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

AO22x1_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_57),
.B1(n_60),
.B2(n_20),
.Y(n_110)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_94),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_83),
.B1(n_67),
.B2(n_25),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_30),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_74),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_93),
.B(n_80),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_134),
.B(n_108),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_121),
.B(n_125),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_68),
.B1(n_86),
.B2(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_132),
.B1(n_143),
.B2(n_100),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_75),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_123),
.B(n_126),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_69),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_136),
.C(n_103),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_117),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_140),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_102),
.A2(n_73),
.B1(n_92),
.B2(n_82),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_91),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_90),
.B(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_16),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_116),
.B1(n_106),
.B2(n_119),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_138),
.Y(n_156)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_139),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_113),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_114),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_67),
.B1(n_25),
.B2(n_77),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_144),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_146),
.A2(n_162),
.B1(n_156),
.B2(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_154),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_97),
.B(n_111),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_155),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_157),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_111),
.B(n_109),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_143),
.B(n_128),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_124),
.C(n_136),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_167),
.C(n_169),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_166),
.B(n_155),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_161),
.A2(n_120),
.B(n_125),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_142),
.C(n_130),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_120),
.B(n_123),
.C(n_131),
.D(n_127),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_159),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_132),
.C(n_137),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_177),
.B1(n_162),
.B2(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_96),
.C(n_115),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_96),
.C(n_115),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_105),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_172),
.A2(n_149),
.B(n_146),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_172),
.C(n_165),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_145),
.C(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_183),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_182),
.B(n_184),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_170),
.A2(n_152),
.B1(n_14),
.B2(n_13),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_152),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_186),
.A2(n_152),
.B(n_169),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_187),
.A2(n_192),
.B(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_174),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_191),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_194),
.A3(n_197),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_200)
);

O2A1O1Ixp5_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_180),
.B(n_178),
.C(n_175),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_0),
.B(n_2),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_190),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_78),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_199),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_193),
.C(n_196),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_202),
.A2(n_198),
.B1(n_8),
.B2(n_9),
.Y(n_203)
);

AOI321xp33_ASAP7_75t_L g204 ( 
.A1(n_203),
.A2(n_11),
.A3(n_12),
.B1(n_201),
.B2(n_196),
.C(n_194),
.Y(n_204)
);


endmodule