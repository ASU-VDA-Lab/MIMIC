module real_jpeg_27711_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_0),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_56),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_0),
.A2(n_33),
.B1(n_35),
.B2(n_56),
.Y(n_133)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_1),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_65),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_65),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_2),
.A2(n_33),
.B1(n_35),
.B2(n_65),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_3),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_171),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_171),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_3),
.A2(n_33),
.B1(n_35),
.B2(n_171),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_53),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_33),
.B1(n_35),
.B2(n_53),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_6),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_6),
.B(n_59),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_46),
.Y(n_229)
);

AOI21xp33_ASAP7_75t_L g233 ( 
.A1(n_6),
.A2(n_46),
.B(n_229),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_190),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_6),
.A2(n_30),
.B(n_33),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_6),
.B(n_138),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_6),
.A2(n_86),
.B1(n_89),
.B2(n_277),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_8),
.A2(n_63),
.B1(n_64),
.B2(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_8),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_142),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_142),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_8),
.A2(n_33),
.B1(n_35),
.B2(n_142),
.Y(n_264)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_10),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_10),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_113)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_12),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_12),
.A2(n_46),
.B1(n_47),
.B2(n_192),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_192),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_12),
.A2(n_33),
.B1(n_35),
.B2(n_192),
.Y(n_277)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_15),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_102),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_83),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_21),
.A2(n_22),
.B1(n_73),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_57),
.B1(n_71),
.B2(n_72),
.Y(n_22)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_39),
.B2(n_40),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_24),
.A2(n_25),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_40),
.C(n_57),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_36),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_26),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_26),
.A2(n_32),
.B1(n_97),
.B2(n_136),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_26),
.A2(n_36),
.B(n_98),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_26),
.A2(n_32),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_26),
.A2(n_78),
.B(n_237),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_26),
.A2(n_32),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_26),
.A2(n_32),
.B1(n_236),
.B2(n_254),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_32),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_29),
.B1(n_44),
.B2(n_49),
.Y(n_50)
);

AOI32xp33_ASAP7_75t_L g227 ( 
.A1(n_28),
.A2(n_47),
.A3(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_29),
.B(n_44),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_29),
.A2(n_31),
.B(n_190),
.C(n_256),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_32),
.A2(n_80),
.B(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_32),
.B(n_190),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_33),
.Y(n_35)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_35),
.B(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_37),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_51),
.B(n_54),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_41),
.A2(n_54),
.B(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_41),
.A2(n_112),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_50),
.B1(n_52),
.B2(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_42),
.B(n_55),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_42),
.A2(n_50),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_42),
.A2(n_50),
.B1(n_186),
.B2(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_42),
.A2(n_50),
.B1(n_215),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_43)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_44),
.Y(n_228)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_46),
.A2(n_47),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_46),
.B(n_60),
.Y(n_203)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_47),
.A2(n_68),
.B1(n_189),
.B2(n_203),
.Y(n_202)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_50),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_50),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_72),
.B1(n_104),
.B2(n_116),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B(n_66),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_58),
.B(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_62),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_58),
.A2(n_106),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_58),
.A2(n_106),
.B1(n_170),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_60),
.B(n_64),
.C(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_59),
.B(n_100),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_59),
.A2(n_67),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_64),
.Y(n_68)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g189 ( 
.A(n_64),
.B(n_190),
.CON(n_189),
.SN(n_189)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_73),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_114),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_83),
.A2(n_84),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_95),
.B(n_99),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_99),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_85),
.A2(n_96),
.B1(n_125),
.B2(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_90),
.B(n_93),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_86),
.A2(n_160),
.B(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_86),
.A2(n_160),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_86),
.A2(n_134),
.B(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_86),
.A2(n_89),
.B1(n_269),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_132),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_87),
.A2(n_94),
.B(n_162),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_87),
.A2(n_91),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_89),
.B(n_190),
.Y(n_281)
);

INVx5_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_94),
.Y(n_134)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_91),
.Y(n_206)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_96),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_117),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_115),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_141),
.B(n_143),
.Y(n_140)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_113),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_148),
.B(n_321),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_144),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_121),
.B(n_144),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_127),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_126),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_127),
.A2(n_128),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_137),
.C(n_139),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_135),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_130),
.B(n_135),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_131),
.A2(n_205),
.B(n_206),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_139),
.B1(n_140),
.B2(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_137),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_175),
.B(n_320),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_172),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_150),
.B(n_172),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_157),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_155),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_157),
.B(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_166),
.C(n_168),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_158),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_165),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_165),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_166),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_314),
.B(n_319),
.Y(n_175)
);

O2A1O1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_219),
.B(n_300),
.C(n_313),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_207),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_178),
.B(n_207),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_193),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_180),
.B(n_181),
.C(n_193),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_188),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_188),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_201),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_195),
.B(n_199),
.C(n_201),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_213),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_208),
.A2(n_209),
.B1(n_295),
.B2(n_297),
.Y(n_294)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.C(n_218),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_218),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_299),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_292),
.B(n_298),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_247),
.B(n_291),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_238),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_223),
.B(n_238),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_231),
.C(n_234),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_224),
.A2(n_225),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_227),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_243),
.B2(n_244),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_245),
.C(n_246),
.Y(n_293)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_285),
.B(n_290),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_265),
.B(n_284),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_250),
.B(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_255),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_255),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_263),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_262),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_273),
.B(n_283),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_271),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_267),
.B(n_271),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_278),
.B(n_282),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_293),
.B(n_294),
.Y(n_298)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_295),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_311),
.B2(n_312),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_308),
.C(n_312),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_316),
.Y(n_319)
);


endmodule