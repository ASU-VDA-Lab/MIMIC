module fake_netlist_5_843_n_5624 (n_82, n_10, n_24, n_86, n_83, n_61, n_75, n_65, n_78, n_74, n_57, n_37, n_31, n_13, n_66, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_38, n_80, n_4, n_35, n_73, n_17, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_62, n_71, n_85, n_59, n_26, n_55, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_27, n_64, n_77, n_81, n_28, n_70, n_68, n_72, n_32, n_41, n_56, n_51, n_63, n_11, n_7, n_15, n_48, n_50, n_52, n_5624);

input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_37;
input n_31;
input n_13;
input n_66;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_62;
input n_71;
input n_85;
input n_59;
input n_26;
input n_55;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_70;
input n_68;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;

output n_5624;

wire n_924;
wire n_977;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_4706;
wire n_5567;
wire n_2380;
wire n_3241;
wire n_3006;
wire n_532;
wire n_5287;
wire n_2327;
wire n_1488;
wire n_2899;
wire n_790;
wire n_5484;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2395;
wire n_5161;
wire n_5512;
wire n_5207;
wire n_2347;
wire n_4963;
wire n_4240;
wire n_4508;
wire n_2021;
wire n_2391;
wire n_5035;
wire n_5282;
wire n_1960;
wire n_2843;
wire n_551;
wire n_3615;
wire n_2059;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_3202;
wire n_4977;
wire n_3813;
wire n_671;
wire n_3341;
wire n_3587;
wire n_4128;
wire n_3445;
wire n_2001;
wire n_4145;
wire n_3785;
wire n_5033;
wire n_1462;
wire n_4211;
wire n_3448;
wire n_3019;
wire n_2096;
wire n_877;
wire n_3776;
wire n_2530;
wire n_4517;
wire n_1696;
wire n_2483;
wire n_4425;
wire n_4950;
wire n_4988;
wire n_1285;
wire n_1860;
wire n_4615;
wire n_87;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_5480;
wire n_668;
wire n_301;
wire n_2147;
wire n_3010;
wire n_2770;
wire n_4131;
wire n_5402;
wire n_2584;
wire n_171;
wire n_3188;
wire n_5509;
wire n_3403;
wire n_3624;
wire n_3461;
wire n_3082;
wire n_2189;
wire n_3796;
wire n_5154;
wire n_1242;
wire n_3283;
wire n_519;
wire n_5469;
wire n_2323;
wire n_2597;
wire n_3340;
wire n_3277;
wire n_5453;
wire n_281;
wire n_2052;
wire n_4499;
wire n_4927;
wire n_731;
wire n_5202;
wire n_1314;
wire n_1512;
wire n_1490;
wire n_317;
wire n_569;
wire n_3214;
wire n_1517;
wire n_2091;
wire n_4311;
wire n_3631;
wire n_3806;
wire n_4691;
wire n_1449;
wire n_4678;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2587;
wire n_156;
wire n_5406;
wire n_219;
wire n_157;
wire n_3947;
wire n_3490;
wire n_600;
wire n_223;
wire n_1948;
wire n_3868;
wire n_3183;
wire n_3437;
wire n_3353;
wire n_264;
wire n_4203;
wire n_3687;
wire n_5241;
wire n_882;
wire n_2384;
wire n_3156;
wire n_696;
wire n_3376;
wire n_646;
wire n_5037;
wire n_436;
wire n_4468;
wire n_3653;
wire n_5562;
wire n_3702;
wire n_1040;
wire n_4976;
wire n_2202;
wire n_2648;
wire n_5008;
wire n_2159;
wire n_2976;
wire n_3876;
wire n_2353;
wire n_2439;
wire n_4811;
wire n_5398;
wire n_2276;
wire n_2089;
wire n_3420;
wire n_1561;
wire n_1165;
wire n_5144;
wire n_1034;
wire n_3361;
wire n_4758;
wire n_1600;
wire n_521;
wire n_845;
wire n_528;
wire n_4255;
wire n_1796;
wire n_5577;
wire n_395;
wire n_553;
wire n_901;
wire n_4484;
wire n_3668;
wire n_4237;
wire n_2934;
wire n_1672;
wire n_1880;
wire n_3550;
wire n_1626;
wire n_637;
wire n_144;
wire n_2079;
wire n_2238;
wire n_96;
wire n_1151;
wire n_1405;
wire n_1706;
wire n_3418;
wire n_342;
wire n_4901;
wire n_197;
wire n_2859;
wire n_1075;
wire n_3395;
wire n_4917;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_2968;
wire n_1585;
wire n_2684;
wire n_3593;
wire n_5343;
wire n_1599;
wire n_4421;
wire n_4836;
wire n_5062;
wire n_4020;
wire n_2730;
wire n_2251;
wire n_3915;
wire n_1377;
wire n_4469;
wire n_4414;
wire n_190;
wire n_5184;
wire n_4532;
wire n_3339;
wire n_228;
wire n_283;
wire n_3349;
wire n_3735;
wire n_2248;
wire n_3007;
wire n_1000;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_5463;
wire n_2100;
wire n_5236;
wire n_310;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_3983;
wire n_332;
wire n_1053;
wire n_1224;
wire n_4405;
wire n_5433;
wire n_1926;
wire n_1331;
wire n_4195;
wire n_279;
wire n_1014;
wire n_4969;
wire n_1241;
wire n_4504;
wire n_1385;
wire n_440;
wire n_793;
wire n_2776;
wire n_4408;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_4531;
wire n_476;
wire n_2987;
wire n_1527;
wire n_4567;
wire n_4164;
wire n_5315;
wire n_4234;
wire n_345;
wire n_4130;
wire n_3611;
wire n_2862;
wire n_5348;
wire n_2175;
wire n_5055;
wire n_2324;
wire n_2606;
wire n_3187;
wire n_2828;
wire n_5397;
wire n_182;
wire n_4471;
wire n_5031;
wire n_407;
wire n_3392;
wire n_3975;
wire n_3430;
wire n_4444;
wire n_3208;
wire n_207;
wire n_3331;
wire n_2379;
wire n_4983;
wire n_2911;
wire n_2154;
wire n_4916;
wire n_3649;
wire n_4302;
wire n_2514;
wire n_5189;
wire n_5381;
wire n_4786;
wire n_3257;
wire n_1027;
wire n_326;
wire n_4160;
wire n_2293;
wire n_5516;
wire n_4051;
wire n_2028;
wire n_558;
wire n_3009;
wire n_1276;
wire n_1412;
wire n_3981;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1841;
wire n_154;
wire n_2581;
wire n_3224;
wire n_4647;
wire n_3752;
wire n_870;
wire n_1711;
wire n_1891;
wire n_5254;
wire n_434;
wire n_3526;
wire n_2546;
wire n_965;
wire n_3790;
wire n_3491;
wire n_935;
wire n_817;
wire n_1175;
wire n_4613;
wire n_4649;
wire n_1888;
wire n_5615;
wire n_1963;
wire n_4795;
wire n_2226;
wire n_2891;
wire n_4028;
wire n_103;
wire n_97;
wire n_5479;
wire n_1690;
wire n_3819;
wire n_2449;
wire n_5083;
wire n_431;
wire n_1194;
wire n_2297;
wire n_4186;
wire n_4731;
wire n_1759;
wire n_2177;
wire n_3747;
wire n_5592;
wire n_2227;
wire n_4618;
wire n_127;
wire n_2190;
wire n_3346;
wire n_4742;
wire n_2876;
wire n_4099;
wire n_452;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_2479;
wire n_1464;
wire n_4295;
wire n_649;
wire n_5303;
wire n_1444;
wire n_4694;
wire n_4533;
wire n_3038;
wire n_5081;
wire n_5124;
wire n_3068;
wire n_2871;
wire n_4244;
wire n_4603;
wire n_2943;
wire n_4254;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_4697;
wire n_2607;
wire n_4190;
wire n_3994;
wire n_4810;
wire n_3317;
wire n_1121;
wire n_433;
wire n_4391;
wire n_949;
wire n_3263;
wire n_2582;
wire n_4157;
wire n_4283;
wire n_4681;
wire n_1001;
wire n_1503;
wire n_4638;
wire n_1468;
wire n_3455;
wire n_5047;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_5346;
wire n_1994;
wire n_5517;
wire n_1195;
wire n_4707;
wire n_2577;
wire n_4527;
wire n_5109;
wire n_2796;
wire n_757;
wire n_2342;
wire n_106;
wire n_4156;
wire n_1851;
wire n_4848;
wire n_2937;
wire n_3095;
wire n_2805;
wire n_1145;
wire n_524;
wire n_394;
wire n_4918;
wire n_1153;
wire n_3856;
wire n_741;
wire n_2914;
wire n_4898;
wire n_1964;
wire n_2869;
wire n_4002;
wire n_1163;
wire n_1207;
wire n_5010;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_2925;
wire n_3773;
wire n_3918;
wire n_2398;
wire n_2857;
wire n_5358;
wire n_4528;
wire n_3932;
wire n_4619;
wire n_4673;
wire n_940;
wire n_3516;
wire n_4822;
wire n_2155;
wire n_2516;
wire n_3797;
wire n_1596;
wire n_2947;
wire n_123;
wire n_978;
wire n_5580;
wire n_4299;
wire n_4801;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_3515;
wire n_2886;
wire n_267;
wire n_2093;
wire n_2473;
wire n_1208;
wire n_3287;
wire n_3378;
wire n_5435;
wire n_1431;
wire n_4279;
wire n_4769;
wire n_4632;
wire n_5373;
wire n_660;
wire n_4294;
wire n_1732;
wire n_5279;
wire n_4232;
wire n_4125;
wire n_4949;
wire n_374;
wire n_2941;
wire n_2457;
wire n_5493;
wire n_4790;
wire n_459;
wire n_962;
wire n_723;
wire n_2536;
wire n_1336;
wire n_1758;
wire n_2952;
wire n_4847;
wire n_5321;
wire n_3058;
wire n_5096;
wire n_4365;
wire n_1878;
wire n_3505;
wire n_4610;
wire n_88;
wire n_3730;
wire n_4489;
wire n_168;
wire n_974;
wire n_727;
wire n_5210;
wire n_4967;
wire n_957;
wire n_4992;
wire n_3001;
wire n_303;
wire n_3945;
wire n_4542;
wire n_2261;
wire n_2729;
wire n_3597;
wire n_1612;
wire n_2897;
wire n_2077;
wire n_4198;
wire n_2909;
wire n_4534;
wire n_4500;
wire n_5014;
wire n_3185;
wire n_1300;
wire n_1127;
wire n_3523;
wire n_1785;
wire n_2829;
wire n_4597;
wire n_4329;
wire n_1006;
wire n_4087;
wire n_3811;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_2231;
wire n_2017;
wire n_2604;
wire n_4257;
wire n_3453;
wire n_322;
wire n_2390;
wire n_3213;
wire n_1041;
wire n_3077;
wire n_1562;
wire n_383;
wire n_3474;
wire n_3984;
wire n_239;
wire n_630;
wire n_2151;
wire n_2106;
wire n_2716;
wire n_4665;
wire n_1913;
wire n_1823;
wire n_3679;
wire n_3422;
wire n_3888;
wire n_4189;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_3707;
wire n_1846;
wire n_5584;
wire n_3429;
wire n_1903;
wire n_3849;
wire n_3946;
wire n_860;
wire n_3229;
wire n_4463;
wire n_1805;
wire n_429;
wire n_4687;
wire n_948;
wire n_4670;
wire n_4084;
wire n_4703;
wire n_4037;
wire n_2922;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2727;
wire n_560;
wire n_340;
wire n_3421;
wire n_2240;
wire n_2436;
wire n_1552;
wire n_3618;
wire n_574;
wire n_2593;
wire n_5262;
wire n_3683;
wire n_3642;
wire n_3286;
wire n_3808;
wire n_824;
wire n_359;
wire n_1327;
wire n_4763;
wire n_1684;
wire n_3590;
wire n_5310;
wire n_366;
wire n_815;
wire n_4594;
wire n_3424;
wire n_1381;
wire n_1037;
wire n_2301;
wire n_3583;
wire n_3560;
wire n_4076;
wire n_4714;
wire n_2419;
wire n_3215;
wire n_5146;
wire n_589;
wire n_4776;
wire n_2122;
wire n_2512;
wire n_4102;
wire n_2786;
wire n_3171;
wire n_1437;
wire n_645;
wire n_238;
wire n_5213;
wire n_3020;
wire n_3677;
wire n_3462;
wire n_5441;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_222;
wire n_1123;
wire n_1467;
wire n_2163;
wire n_634;
wire n_2254;
wire n_1382;
wire n_925;
wire n_3546;
wire n_424;
wire n_2647;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_4443;
wire n_5461;
wire n_4507;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_4575;
wire n_380;
wire n_419;
wire n_3244;
wire n_389;
wire n_3130;
wire n_3822;
wire n_3569;
wire n_912;
wire n_136;
wire n_968;
wire n_4452;
wire n_4348;
wire n_5430;
wire n_619;
wire n_5362;
wire n_376;
wire n_4355;
wire n_3494;
wire n_515;
wire n_351;
wire n_5050;
wire n_885;
wire n_5063;
wire n_5229;
wire n_2125;
wire n_3771;
wire n_5199;
wire n_683;
wire n_3110;
wire n_1057;
wire n_1051;
wire n_721;
wire n_1157;
wire n_3073;
wire n_4572;
wire n_5527;
wire n_802;
wire n_5609;
wire n_5416;
wire n_4026;
wire n_2265;
wire n_4104;
wire n_1608;
wire n_4512;
wire n_3554;
wire n_4377;
wire n_280;
wire n_1305;
wire n_5266;
wire n_3178;
wire n_873;
wire n_5355;
wire n_2334;
wire n_690;
wire n_4521;
wire n_583;
wire n_4488;
wire n_2289;
wire n_3051;
wire n_302;
wire n_1343;
wire n_2783;
wire n_2263;
wire n_3750;
wire n_2341;
wire n_3632;
wire n_4588;
wire n_2733;
wire n_1288;
wire n_212;
wire n_2785;
wire n_2415;
wire n_3299;
wire n_4519;
wire n_5551;
wire n_3715;
wire n_972;
wire n_3040;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_3568;
wire n_5475;
wire n_3737;
wire n_1185;
wire n_991;
wire n_1967;
wire n_576;
wire n_1329;
wire n_3255;
wire n_4856;
wire n_2997;
wire n_4400;
wire n_5168;
wire n_943;
wire n_3326;
wire n_3734;
wire n_650;
wire n_4778;
wire n_286;
wire n_2429;
wire n_883;
wire n_470;
wire n_325;
wire n_132;
wire n_5322;
wire n_856;
wire n_1793;
wire n_4352;
wire n_4441;
wire n_918;
wire n_4761;
wire n_942;
wire n_1804;
wire n_189;
wire n_4347;
wire n_4095;
wire n_3196;
wire n_4593;
wire n_2364;
wire n_2533;
wire n_3492;
wire n_2780;
wire n_4727;
wire n_4568;
wire n_5371;
wire n_195;
wire n_2291;
wire n_4043;
wire n_1636;
wire n_3601;
wire n_5418;
wire n_1350;
wire n_1865;
wire n_2973;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_2393;
wire n_1697;
wire n_5316;
wire n_3831;
wire n_3801;
wire n_225;
wire n_2043;
wire n_2751;
wire n_192;
wire n_4893;
wire n_5032;
wire n_1549;
wire n_1934;
wire n_4948;
wire n_4000;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1446;
wire n_4406;
wire n_2758;
wire n_1458;
wire n_472;
wire n_1807;
wire n_387;
wire n_2618;
wire n_398;
wire n_5112;
wire n_5386;
wire n_2559;
wire n_763;
wire n_4748;
wire n_2295;
wire n_3931;
wire n_1219;
wire n_4010;
wire n_2840;
wire n_5017;
wire n_1814;
wire n_2822;
wire n_4710;
wire n_287;
wire n_555;
wire n_4607;
wire n_5123;
wire n_4117;
wire n_3636;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_4487;
wire n_5001;
wire n_2795;
wire n_2981;
wire n_2282;
wire n_2800;
wire n_4817;
wire n_311;
wire n_3380;
wire n_2098;
wire n_1296;
wire n_3460;
wire n_3409;
wire n_3538;
wire n_2068;
wire n_4849;
wire n_4867;
wire n_5424;
wire n_445;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_4728;
wire n_588;
wire n_789;
wire n_4247;
wire n_4933;
wire n_107;
wire n_4018;
wire n_3900;
wire n_1105;
wire n_4902;
wire n_4518;
wire n_4409;
wire n_4411;
wire n_3872;
wire n_4336;
wire n_149;
wire n_2270;
wire n_4777;
wire n_2653;
wire n_836;
wire n_2496;
wire n_1908;
wire n_2259;
wire n_3877;
wire n_458;
wire n_2995;
wire n_5496;
wire n_2494;
wire n_3547;
wire n_3977;
wire n_1102;
wire n_4052;
wire n_3459;
wire n_1499;
wire n_4398;
wire n_3155;
wire n_2633;
wire n_4954;
wire n_2435;
wire n_1392;
wire n_1164;
wire n_2097;
wire n_5460;
wire n_4304;
wire n_3911;
wire n_5333;
wire n_1303;
wire n_4431;
wire n_4192;
wire n_5570;
wire n_3736;
wire n_4805;
wire n_118;
wire n_601;
wire n_4885;
wire n_253;
wire n_1661;
wire n_3565;
wire n_172;
wire n_4701;
wire n_2575;
wire n_5040;
wire n_861;
wire n_1658;
wire n_1904;
wire n_1345;
wire n_176;
wire n_1899;
wire n_1003;
wire n_2067;
wire n_2219;
wire n_3533;
wire n_2877;
wire n_2148;
wire n_393;
wire n_4631;
wire n_1726;
wire n_3035;
wire n_421;
wire n_5194;
wire n_5464;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_3639;
wire n_708;
wire n_735;
wire n_2501;
wire n_3079;
wire n_4965;
wire n_1915;
wire n_5610;
wire n_1109;
wire n_5239;
wire n_1310;
wire n_2605;
wire n_4747;
wire n_5197;
wire n_1399;
wire n_1979;
wire n_193;
wire n_2924;
wire n_4111;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_4587;
wire n_3731;
wire n_2946;
wire n_5305;
wire n_4538;
wire n_435;
wire n_766;
wire n_541;
wire n_1117;
wire n_2754;
wire n_687;
wire n_1742;
wire n_5376;
wire n_2489;
wire n_536;
wire n_5204;
wire n_2012;
wire n_1291;
wire n_4094;
wire n_3503;
wire n_2866;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_2917;
wire n_2425;
wire n_3536;
wire n_3661;
wire n_4150;
wire n_827;
wire n_4878;
wire n_1703;
wire n_1650;
wire n_1137;
wire n_3934;
wire n_4985;
wire n_3922;
wire n_3846;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_2498;
wire n_2697;
wire n_850;
wire n_3074;
wire n_1999;
wire n_2372;
wire n_3673;
wire n_3768;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_3943;
wire n_353;
wire n_2430;
wire n_493;
wire n_2433;
wire n_3293;
wire n_5508;
wire n_5582;
wire n_4022;
wire n_1531;
wire n_840;
wire n_1334;
wire n_4852;
wire n_2528;
wire n_4869;
wire n_4700;
wire n_4035;
wire n_2316;
wire n_1898;
wire n_3294;
wire n_4426;
wire n_554;
wire n_3415;
wire n_2284;
wire n_2817;
wire n_3139;
wire n_5292;
wire n_2598;
wire n_4601;
wire n_2687;
wire n_1120;
wire n_198;
wire n_1890;
wire n_714;
wire n_4220;
wire n_1944;
wire n_909;
wire n_1497;
wire n_3431;
wire n_3169;
wire n_3151;
wire n_2078;
wire n_3284;
wire n_3070;
wire n_4066;
wire n_119;
wire n_2884;
wire n_4515;
wire n_4351;
wire n_5264;
wire n_3126;
wire n_4403;
wire n_1981;
wire n_1663;
wire n_1718;
wire n_4509;
wire n_4858;
wire n_3700;
wire n_5504;
wire n_509;
wire n_147;
wire n_1518;
wire n_4223;
wire n_1281;
wire n_1889;
wire n_209;
wire n_1489;
wire n_5025;
wire n_2966;
wire n_1376;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_186;
wire n_756;
wire n_1429;
wire n_4644;
wire n_4456;
wire n_5060;
wire n_399;
wire n_5334;
wire n_2448;
wire n_4346;
wire n_3170;
wire n_2748;
wire n_3311;
wire n_3272;
wire n_2898;
wire n_2717;
wire n_1861;
wire n_760;
wire n_5581;
wire n_3691;
wire n_3628;
wire n_220;
wire n_4235;
wire n_1867;
wire n_1945;
wire n_3018;
wire n_481;
wire n_2573;
wire n_4435;
wire n_2939;
wire n_3807;
wire n_271;
wire n_2447;
wire n_4764;
wire n_886;
wire n_1221;
wire n_5394;
wire n_167;
wire n_2774;
wire n_1707;
wire n_853;
wire n_4655;
wire n_3161;
wire n_377;
wire n_4581;
wire n_751;
wire n_4827;
wire n_2488;
wire n_392;
wire n_3477;
wire n_5421;
wire n_2476;
wire n_704;
wire n_4399;
wire n_2781;
wire n_5309;
wire n_2778;
wire n_771;
wire n_4782;
wire n_1520;
wire n_4363;
wire n_2887;
wire n_1287;
wire n_4864;
wire n_1262;
wire n_2691;
wire n_1411;
wire n_3054;
wire n_4335;
wire n_2526;
wire n_2703;
wire n_2167;
wire n_5428;
wire n_3391;
wire n_4259;
wire n_5541;
wire n_2709;
wire n_5543;
wire n_816;
wire n_1536;
wire n_4865;
wire n_4056;
wire n_1344;
wire n_4564;
wire n_1246;
wire n_3840;
wire n_1339;
wire n_5085;
wire n_3518;
wire n_2956;
wire n_3733;
wire n_328;
wire n_2173;
wire n_1842;
wire n_871;
wire n_3738;
wire n_685;
wire n_5116;
wire n_3464;
wire n_2018;
wire n_4526;
wire n_1555;
wire n_3245;
wire n_4417;
wire n_499;
wire n_98;
wire n_402;
wire n_4899;
wire n_796;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1012;
wire n_5411;
wire n_2453;
wire n_4798;
wire n_1525;
wire n_740;
wire n_3509;
wire n_3352;
wire n_3076;
wire n_3535;
wire n_2182;
wire n_277;
wire n_1061;
wire n_3251;
wire n_92;
wire n_2931;
wire n_5185;
wire n_1193;
wire n_3118;
wire n_3511;
wire n_1226;
wire n_3443;
wire n_2146;
wire n_1487;
wire n_3644;
wire n_5076;
wire n_3336;
wire n_3935;
wire n_781;
wire n_542;
wire n_3521;
wire n_5379;
wire n_3562;
wire n_3948;
wire n_4750;
wire n_1515;
wire n_2918;
wire n_3232;
wire n_1673;
wire n_2112;
wire n_1739;
wire n_2958;
wire n_3114;
wire n_3125;
wire n_4981;
wire n_2394;
wire n_3612;
wire n_2954;
wire n_4835;
wire n_4430;
wire n_5565;
wire n_4081;
wire n_1103;
wire n_3132;
wire n_4407;
wire n_648;
wire n_312;
wire n_3951;
wire n_4894;
wire n_3238;
wire n_3210;
wire n_2036;
wire n_3267;
wire n_4995;
wire n_480;
wire n_425;
wire n_695;
wire n_5524;
wire n_3964;
wire n_3772;
wire n_229;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_4446;
wire n_3884;
wire n_3726;
wire n_805;
wire n_2525;
wire n_2892;
wire n_113;
wire n_2907;
wire n_3577;
wire n_2820;
wire n_269;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1741;
wire n_1160;
wire n_4057;
wire n_4332;
wire n_1258;
wire n_4314;
wire n_1074;
wire n_3347;
wire n_3216;
wire n_1621;
wire n_3809;
wire n_2113;
wire n_1448;
wire n_4288;
wire n_3567;
wire n_5066;
wire n_1634;
wire n_3939;
wire n_5401;
wire n_4241;
wire n_3321;
wire n_3212;
wire n_666;
wire n_1433;
wire n_2256;
wire n_3152;
wire n_5106;
wire n_319;
wire n_5468;
wire n_2920;
wire n_4265;
wire n_1186;
wire n_5319;
wire n_1018;
wire n_2247;
wire n_713;
wire n_1622;
wire n_166;
wire n_1180;
wire n_3705;
wire n_2802;
wire n_4705;
wire n_3159;
wire n_5455;
wire n_2268;
wire n_3778;
wire n_5337;
wire n_3304;
wire n_1378;
wire n_3912;
wire n_1729;
wire n_2739;
wire n_469;
wire n_2771;
wire n_4604;
wire n_549;
wire n_5223;
wire n_3795;
wire n_5020;
wire n_4419;
wire n_4477;
wire n_3179;
wire n_3256;
wire n_667;
wire n_2386;
wire n_1501;
wire n_3086;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_4217;
wire n_4395;
wire n_2821;
wire n_5074;
wire n_1099;
wire n_2568;
wire n_5364;
wire n_564;
wire n_1738;
wire n_3728;
wire n_3064;
wire n_3088;
wire n_1021;
wire n_4639;
wire n_3713;
wire n_3663;
wire n_5046;
wire n_5166;
wire n_3246;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_819;
wire n_5088;
wire n_2302;
wire n_5457;
wire n_951;
wire n_5532;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_2069;
wire n_417;
wire n_3434;
wire n_1806;
wire n_933;
wire n_1563;
wire n_4227;
wire n_4033;
wire n_4289;
wire n_2024;
wire n_4780;
wire n_755;
wire n_4243;
wire n_4982;
wire n_530;
wire n_4330;
wire n_3695;
wire n_556;
wire n_2482;
wire n_2677;
wire n_5544;
wire n_3832;
wire n_3987;
wire n_902;
wire n_5352;
wire n_4991;
wire n_5538;
wire n_579;
wire n_1698;
wire n_2329;
wire n_1098;
wire n_2142;
wire n_320;
wire n_5410;
wire n_3332;
wire n_1135;
wire n_3048;
wire n_3937;
wire n_2203;
wire n_4525;
wire n_1243;
wire n_101;
wire n_3782;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_4208;
wire n_3786;
wire n_371;
wire n_2888;
wire n_3638;
wire n_5503;
wire n_1236;
wire n_1633;
wire n_4177;
wire n_3763;
wire n_2669;
wire n_1778;
wire n_2306;
wire n_3022;
wire n_4264;
wire n_335;
wire n_3087;
wire n_3489;
wire n_2566;
wire n_343;
wire n_308;
wire n_5129;
wire n_2149;
wire n_1078;
wire n_5500;
wire n_3060;
wire n_4276;
wire n_5219;
wire n_5605;
wire n_3013;
wire n_1984;
wire n_5170;
wire n_2408;
wire n_5320;
wire n_1877;
wire n_3049;
wire n_1723;
wire n_5107;
wire n_339;
wire n_4485;
wire n_183;
wire n_4626;
wire n_1036;
wire n_1097;
wire n_347;
wire n_798;
wire n_2659;
wire n_1414;
wire n_290;
wire n_4975;
wire n_1852;
wire n_578;
wire n_344;
wire n_5602;
wire n_3089;
wire n_422;
wire n_2470;
wire n_5405;
wire n_3985;
wire n_5253;
wire n_496;
wire n_1391;
wire n_670;
wire n_4760;
wire n_4652;
wire n_4624;
wire n_663;
wire n_2551;
wire n_1587;
wire n_2682;
wire n_813;
wire n_1284;
wire n_3440;
wire n_1748;
wire n_4569;
wire n_2699;
wire n_4897;
wire n_888;
wire n_2769;
wire n_3542;
wire n_3436;
wire n_5491;
wire n_2615;
wire n_3940;
wire n_446;
wire n_1064;
wire n_858;
wire n_2985;
wire n_691;
wire n_5065;
wire n_2753;
wire n_363;
wire n_1582;
wire n_3637;
wire n_2842;
wire n_4523;
wire n_1836;
wire n_2868;
wire n_5492;
wire n_3141;
wire n_5084;
wire n_3164;
wire n_3570;
wire n_5260;
wire n_4919;
wire n_4025;
wire n_461;
wire n_2712;
wire n_5328;
wire n_3936;
wire n_4503;
wire n_3507;
wire n_3821;
wire n_2700;
wire n_1211;
wire n_3367;
wire n_4464;
wire n_907;
wire n_3096;
wire n_3496;
wire n_4114;
wire n_989;
wire n_2544;
wire n_2356;
wire n_488;
wire n_892;
wire n_4556;
wire n_5454;
wire n_2620;
wire n_1581;
wire n_4089;
wire n_5621;
wire n_586;
wire n_2919;
wire n_4327;
wire n_230;
wire n_953;
wire n_4218;
wire n_2150;
wire n_3146;
wire n_5165;
wire n_2241;
wire n_2757;
wire n_963;
wire n_1052;
wire n_954;
wire n_5573;
wire n_478;
wire n_4353;
wire n_2042;
wire n_534;
wire n_884;
wire n_1754;
wire n_1623;
wire n_2921;
wire n_2720;
wire n_1854;
wire n_4990;
wire n_5529;
wire n_1856;
wire n_143;
wire n_4959;
wire n_4161;
wire n_237;
wire n_832;
wire n_1319;
wire n_3992;
wire n_2616;
wire n_1906;
wire n_4103;
wire n_1387;
wire n_4466;
wire n_2262;
wire n_2462;
wire n_1532;
wire n_3625;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_686;
wire n_2837;
wire n_847;
wire n_4844;
wire n_2979;
wire n_5257;
wire n_3655;
wire n_4688;
wire n_4765;
wire n_702;
wire n_2548;
wire n_822;
wire n_5180;
wire n_2108;
wire n_3640;
wire n_4388;
wire n_4206;
wire n_1538;
wire n_1779;
wire n_4738;
wire n_1369;
wire n_3909;
wire n_3207;
wire n_3944;
wire n_809;
wire n_4434;
wire n_4837;
wire n_3042;
wire n_1942;
wire n_2510;
wire n_4219;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_411;
wire n_414;
wire n_5012;
wire n_1293;
wire n_1876;
wire n_4620;
wire n_1810;
wire n_2813;
wire n_4438;
wire n_2009;
wire n_2222;
wire n_3510;
wire n_3218;
wire n_2667;
wire n_3150;
wire n_747;
wire n_4325;
wire n_1733;
wire n_2413;
wire n_615;
wire n_851;
wire n_843;
wire n_705;
wire n_4133;
wire n_3775;
wire n_678;
wire n_4184;
wire n_5203;
wire n_2518;
wire n_2629;
wire n_367;
wire n_4481;
wire n_3416;
wire n_4379;
wire n_2181;
wire n_1829;
wire n_547;
wire n_4030;
wire n_116;
wire n_4490;
wire n_3138;
wire n_4397;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_4820;
wire n_590;
wire n_3770;
wire n_1308;
wire n_5094;
wire n_4938;
wire n_4179;
wire n_3469;
wire n_5336;
wire n_372;
wire n_677;
wire n_2723;
wire n_368;
wire n_314;
wire n_3220;
wire n_4641;
wire n_2539;
wire n_5548;
wire n_5601;
wire n_100;
wire n_3855;
wire n_1008;
wire n_2054;
wire n_5339;
wire n_1559;
wire n_4931;
wire n_1765;
wire n_3158;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_295;
wire n_133;
wire n_3113;
wire n_2718;
wire n_3760;
wire n_4078;
wire n_1760;
wire n_568;
wire n_2856;
wire n_1832;
wire n_4146;
wire n_4360;
wire n_3666;
wire n_3828;
wire n_93;
wire n_3288;
wire n_5514;
wire n_4404;
wire n_5091;
wire n_1509;
wire n_1874;
wire n_4787;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_3667;
wire n_878;
wire n_5486;
wire n_1306;
wire n_3703;
wire n_4903;
wire n_3558;
wire n_2545;
wire n_2787;
wire n_5599;
wire n_906;
wire n_919;
wire n_4356;
wire n_658;
wire n_2061;
wire n_4432;
wire n_5251;
wire n_2378;
wire n_1740;
wire n_1586;
wire n_4291;
wire n_535;
wire n_5403;
wire n_4386;
wire n_4149;
wire n_1492;
wire n_592;
wire n_1692;
wire n_2982;
wire n_2481;
wire n_3545;
wire n_2507;
wire n_4019;
wire n_2900;
wire n_1095;
wire n_1614;
wire n_2339;
wire n_457;
wire n_4637;
wire n_603;
wire n_4935;
wire n_4785;
wire n_3426;
wire n_3820;
wire n_3454;
wire n_5608;
wire n_3741;
wire n_3410;
wire n_2029;
wire n_995;
wire n_1609;
wire n_5298;
wire n_5596;
wire n_396;
wire n_1887;
wire n_4413;
wire n_1073;
wire n_2346;
wire n_662;
wire n_3990;
wire n_4493;
wire n_218;
wire n_3475;
wire n_1215;
wire n_1592;
wire n_2882;
wire n_1721;
wire n_2338;
wire n_3672;
wire n_5290;
wire n_3197;
wire n_3109;
wire n_2721;
wire n_1043;
wire n_5095;
wire n_486;
wire n_3002;
wire n_337;
wire n_5324;
wire n_3897;
wire n_1159;
wire n_3845;
wire n_2081;
wire n_299;
wire n_4570;
wire n_2156;
wire n_5101;
wire n_4296;
wire n_1820;
wire n_5019;
wire n_2418;
wire n_5589;
wire n_2179;
wire n_1416;
wire n_1724;
wire n_2521;
wire n_3458;
wire n_1420;
wire n_1132;
wire n_3330;
wire n_4606;
wire n_4774;
wire n_2477;
wire n_3887;
wire n_4093;
wire n_1486;
wire n_4672;
wire n_3519;
wire n_4174;
wire n_3374;
wire n_3045;
wire n_1870;
wire n_309;
wire n_2367;
wire n_4766;
wire n_2896;
wire n_652;
wire n_1365;
wire n_4074;
wire n_4600;
wire n_1927;
wire n_5583;
wire n_1349;
wire n_4460;
wire n_288;
wire n_1031;
wire n_3645;
wire n_3223;
wire n_3929;
wire n_834;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1965;
wire n_1902;
wire n_1941;
wire n_5501;
wire n_3938;
wire n_5377;
wire n_2878;
wire n_504;
wire n_874;
wire n_3498;
wire n_2015;
wire n_1982;
wire n_4110;
wire n_3189;
wire n_2066;
wire n_993;
wire n_3154;
wire n_1551;
wire n_545;
wire n_450;
wire n_2905;
wire n_3965;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_4349;
wire n_628;
wire n_3788;
wire n_2410;
wire n_4313;
wire n_1084;
wire n_970;
wire n_1935;
wire n_3366;
wire n_1534;
wire n_1351;
wire n_2696;
wire n_4863;
wire n_1205;
wire n_3242;
wire n_495;
wire n_3525;
wire n_3486;
wire n_2405;
wire n_3995;
wire n_2088;
wire n_2953;
wire n_4036;
wire n_921;
wire n_5100;
wire n_1795;
wire n_2578;
wire n_3483;
wire n_128;
wire n_1821;
wire n_3894;
wire n_3478;
wire n_4015;
wire n_3890;
wire n_2740;
wire n_5367;
wire n_2656;
wire n_1080;
wire n_1274;
wire n_3524;
wire n_5616;
wire n_5034;
wire n_1708;
wire n_426;
wire n_562;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2092;
wire n_2075;
wire n_3658;
wire n_1776;
wire n_4807;
wire n_2281;
wire n_2131;
wire n_3026;
wire n_1757;
wire n_890;
wire n_1919;
wire n_960;
wire n_4230;
wire n_3419;
wire n_1290;
wire n_1047;
wire n_2053;
wire n_1958;
wire n_1252;
wire n_348;
wire n_3784;
wire n_2969;
wire n_3941;
wire n_2864;
wire n_3195;
wire n_3190;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_3456;
wire n_444;
wire n_1808;
wire n_316;
wire n_2266;
wire n_2650;
wire n_4428;
wire n_146;
wire n_5003;
wire n_5252;
wire n_408;
wire n_967;
wire n_2731;
wire n_5614;
wire n_5134;
wire n_3953;
wire n_3166;
wire n_4122;
wire n_3976;
wire n_1357;
wire n_3979;
wire n_4582;
wire n_2998;
wire n_4684;
wire n_4840;
wire n_3162;
wire n_983;
wire n_2760;
wire n_3377;
wire n_3749;
wire n_3962;
wire n_1826;
wire n_2304;
wire n_762;
wire n_1283;
wire n_5325;
wire n_2637;
wire n_5375;
wire n_4384;
wire n_4423;
wire n_4096;
wire n_2881;
wire n_1203;
wire n_3282;
wire n_821;
wire n_1763;
wire n_3231;
wire n_1966;
wire n_321;
wire n_4996;
wire n_621;
wire n_2475;
wire n_4598;
wire n_5064;
wire n_4478;
wire n_507;
wire n_2646;
wire n_5536;
wire n_1605;
wire n_5173;
wire n_1228;
wire n_3920;
wire n_4890;
wire n_5027;
wire n_3203;
wire n_3866;
wire n_2903;
wire n_3921;
wire n_828;
wire n_779;
wire n_4106;
wire n_3717;
wire n_2743;
wire n_2675;
wire n_1439;
wire n_3052;
wire n_5215;
wire n_945;
wire n_3743;
wire n_1932;
wire n_4721;
wire n_5597;
wire n_984;
wire n_694;
wire n_1983;
wire n_4029;
wire n_1594;
wire n_900;
wire n_3870;
wire n_4496;
wire n_3529;
wire n_1147;
wire n_1977;
wire n_2153;
wire n_4338;
wire n_3094;
wire n_2310;
wire n_3952;
wire n_2287;
wire n_2860;
wire n_2056;
wire n_1470;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2502;
wire n_2504;
wire n_4762;
wire n_4495;
wire n_2974;
wire n_2901;
wire n_1940;
wire n_2793;
wire n_3442;
wire n_1201;
wire n_1114;
wire n_3998;
wire n_2285;
wire n_3147;
wire n_4141;
wire n_669;
wire n_1176;
wire n_1149;
wire n_1020;
wire n_211;
wire n_5121;
wire n_1824;
wire n_1917;
wire n_3386;
wire n_4107;
wire n_4667;
wire n_2325;
wire n_178;
wire n_5555;
wire n_2446;
wire n_3488;
wire n_1035;
wire n_4547;
wire n_2893;
wire n_2588;
wire n_2962;
wire n_4004;
wire n_661;
wire n_5576;
wire n_4668;
wire n_4953;
wire n_5466;
wire n_3898;
wire n_849;
wire n_584;
wire n_1786;
wire n_430;
wire n_5284;
wire n_4997;
wire n_5308;
wire n_4274;
wire n_2627;
wire n_4759;
wire n_1413;
wire n_801;
wire n_4467;
wire n_2080;
wire n_2377;
wire n_2340;
wire n_3552;
wire n_875;
wire n_357;
wire n_3684;
wire n_4735;
wire n_3137;
wire n_165;
wire n_5578;
wire n_2361;
wire n_1173;
wire n_1603;
wire n_969;
wire n_1401;
wire n_4113;
wire n_1019;
wire n_1998;
wire n_4686;
wire n_5530;
wire n_304;
wire n_3759;
wire n_4321;
wire n_4342;
wire n_2034;
wire n_3933;
wire n_3206;
wire n_5506;
wire n_3966;
wire n_5243;
wire n_5449;
wire n_1702;
wire n_5221;
wire n_4183;
wire n_778;
wire n_1122;
wire n_4068;
wire n_4872;
wire n_4233;
wire n_3192;
wire n_3764;
wire n_4709;
wire n_5038;
wire n_5311;
wire n_2649;
wire n_1187;
wire n_1929;
wire n_5575;
wire n_2807;
wire n_2542;
wire n_2313;
wire n_489;
wire n_1174;
wire n_3324;
wire n_3914;
wire n_4625;
wire n_2558;
wire n_2063;
wire n_3803;
wire n_3742;
wire n_2252;
wire n_4819;
wire n_1685;
wire n_917;
wire n_1714;
wire n_1541;
wire n_2576;
wire n_4900;
wire n_3390;
wire n_1573;
wire n_3746;
wire n_2373;
wire n_1713;
wire n_3817;
wire n_2745;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_2493;
wire n_4930;
wire n_5276;
wire n_1059;
wire n_1133;
wire n_5078;
wire n_4537;
wire n_2885;
wire n_5011;
wire n_3318;
wire n_4070;
wire n_4282;
wire n_3485;
wire n_4180;
wire n_665;
wire n_3839;
wire n_1440;
wire n_5205;
wire n_3333;
wire n_2845;
wire n_4143;
wire n_4659;
wire n_2602;
wire n_205;
wire n_4579;
wire n_4616;
wire n_1496;
wire n_1125;
wire n_3014;
wire n_2547;
wire n_5023;
wire n_1812;
wire n_4105;
wire n_232;
wire n_2532;
wire n_3791;
wire n_2665;
wire n_5351;
wire n_3905;
wire n_427;
wire n_3368;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_2401;
wire n_3135;
wire n_5476;
wire n_2003;
wire n_1457;
wire n_5446;
wire n_4895;
wire n_3573;
wire n_3148;
wire n_2264;
wire n_3534;
wire n_1482;
wire n_4275;
wire n_1266;
wire n_3970;
wire n_3438;
wire n_4098;
wire n_872;
wire n_594;
wire n_200;
wire n_1297;
wire n_4789;
wire n_1972;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_5312;
wire n_985;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_5111;
wire n_4055;
wire n_2926;
wire n_626;
wire n_3540;
wire n_3973;
wire n_3670;
wire n_2023;
wire n_3249;
wire n_2351;
wire n_676;
wire n_5113;
wire n_4442;
wire n_4698;
wire n_642;
wire n_1602;
wire n_194;
wire n_1178;
wire n_4779;
wire n_2286;
wire n_4966;
wire n_503;
wire n_2065;
wire n_4017;
wire n_3397;
wire n_3740;
wire n_620;
wire n_1081;
wire n_4418;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_703;
wire n_1318;
wire n_780;
wire n_2977;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_3600;
wire n_245;
wire n_4134;
wire n_1388;
wire n_2836;
wire n_672;
wire n_581;
wire n_1625;
wire n_2130;
wire n_5167;
wire n_898;
wire n_3239;
wire n_5117;
wire n_2773;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_4913;
wire n_1452;
wire n_5612;
wire n_265;
wire n_443;
wire n_1791;
wire n_2850;
wire n_1747;
wire n_4251;
wire n_1817;
wire n_3982;
wire n_2654;
wire n_4621;
wire n_1326;
wire n_3176;
wire n_4559;
wire n_2186;
wire n_4368;
wire n_4740;
wire n_5301;
wire n_5007;
wire n_3581;
wire n_2562;
wire n_4077;
wire n_4642;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_3576;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_4049;
wire n_941;
wire n_3862;
wire n_5214;
wire n_5487;
wire n_5563;
wire n_3495;
wire n_3879;
wire n_2348;
wire n_5497;
wire n_4724;
wire n_1238;
wire n_1772;
wire n_282;
wire n_752;
wire n_1476;
wire n_1108;
wire n_5526;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_2129;
wire n_3345;
wire n_1395;
wire n_4546;
wire n_862;
wire n_3584;
wire n_3756;
wire n_381;
wire n_2889;
wire n_390;
wire n_5593;
wire n_5021;
wire n_2772;
wire n_5444;
wire n_1675;
wire n_1924;
wire n_4382;
wire n_1554;
wire n_3999;
wire n_2844;
wire n_2138;
wire n_5211;
wire n_5230;
wire n_2260;
wire n_5389;
wire n_1813;
wire n_4833;
wire n_3056;
wire n_2345;
wire n_1172;
wire n_5110;
wire n_379;
wire n_428;
wire n_1341;
wire n_3295;
wire n_2382;
wire n_4719;
wire n_4178;
wire n_3062;
wire n_2317;
wire n_5425;
wire n_3289;
wire n_1973;
wire n_786;
wire n_1142;
wire n_2579;
wire n_1770;
wire n_138;
wire n_4228;
wire n_4401;
wire n_1756;
wire n_1716;
wire n_2788;
wire n_2984;
wire n_3364;
wire n_5560;
wire n_1873;
wire n_3201;
wire n_221;
wire n_622;
wire n_1087;
wire n_3472;
wire n_2874;
wire n_5179;
wire n_4605;
wire n_4877;
wire n_3235;
wire n_4968;
wire n_1272;
wire n_104;
wire n_5030;
wire n_3949;
wire n_3543;
wire n_1247;
wire n_591;
wire n_3050;
wire n_313;
wire n_1478;
wire n_3903;
wire n_4834;
wire n_1210;
wire n_1364;
wire n_5272;
wire n_2183;
wire n_2742;
wire n_3314;
wire n_4158;
wire n_2360;
wire n_3254;
wire n_5361;
wire n_369;
wire n_4171;
wire n_4045;
wire n_598;
wire n_1367;
wire n_4562;
wire n_5068;
wire n_3634;
wire n_1460;
wire n_2834;
wire n_2531;
wire n_517;
wire n_413;
wire n_5015;
wire n_2702;
wire n_2030;
wire n_903;
wire n_3115;
wire n_4749;
wire n_203;
wire n_4390;
wire n_5302;
wire n_4979;
wire n_1404;
wire n_1794;
wire n_2234;
wire n_4804;
wire n_5545;
wire n_2209;
wire n_4270;
wire n_2797;
wire n_1255;
wire n_5152;
wire n_2321;
wire n_722;
wire n_3680;
wire n_844;
wire n_201;
wire n_3497;
wire n_1601;
wire n_5409;
wire n_2940;
wire n_2612;
wire n_1495;
wire n_5128;
wire n_4566;
wire n_979;
wire n_2841;
wire n_3322;
wire n_4576;
wire n_846;
wire n_2427;
wire n_2505;
wire n_4061;
wire n_2070;
wire n_3250;
wire n_585;
wire n_270;
wire n_2594;
wire n_1914;
wire n_2335;
wire n_2904;
wire n_5307;
wire n_4767;
wire n_4328;
wire n_3004;
wire n_3112;
wire n_2349;
wire n_1379;
wire n_3874;
wire n_5415;
wire n_4676;
wire n_4544;
wire n_2170;
wire n_1091;
wire n_641;
wire n_3175;
wire n_3522;
wire n_4429;
wire n_575;
wire n_4591;
wire n_3266;
wire n_4646;
wire n_1130;
wire n_4725;
wire n_4563;
wire n_2210;
wire n_4169;
wire n_5331;
wire n_3247;
wire n_3091;
wire n_3066;
wire n_246;
wire n_2426;
wire n_657;
wire n_4320;
wire n_5341;
wire n_4881;
wire n_491;
wire n_160;
wire n_566;
wire n_565;
wire n_5271;
wire n_5089;
wire n_5263;
wire n_3613;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_4012;
wire n_5518;
wire n_651;
wire n_4636;
wire n_4584;
wire n_5622;
wire n_807;
wire n_3910;
wire n_4711;
wire n_835;
wire n_3319;
wire n_5240;
wire n_3335;
wire n_99;
wire n_3413;
wire n_5495;
wire n_1969;
wire n_4680;
wire n_2044;
wire n_1138;
wire n_5546;
wire n_927;
wire n_2689;
wire n_3259;
wire n_5482;
wire n_4191;
wire n_5224;
wire n_4293;
wire n_2010;
wire n_3688;
wire n_3016;
wire n_1693;
wire n_5393;
wire n_2599;
wire n_904;
wire n_3338;
wire n_3414;
wire n_1827;
wire n_4671;
wire n_4209;
wire n_1271;
wire n_1542;
wire n_5041;
wire n_1423;
wire n_1166;
wire n_1751;
wire n_5431;
wire n_1508;
wire n_785;
wire n_2200;
wire n_3261;
wire n_5026;
wire n_1161;
wire n_3863;
wire n_3027;
wire n_2746;
wire n_1150;
wire n_5059;
wire n_5505;
wire n_3127;
wire n_226;
wire n_1780;
wire n_3732;
wire n_4250;
wire n_5329;
wire n_1055;
wire n_3596;
wire n_4699;
wire n_111;
wire n_3906;
wire n_4127;
wire n_880;
wire n_3297;
wire n_544;
wire n_155;
wire n_2683;
wire n_1370;
wire n_1360;
wire n_2388;
wire n_4292;
wire n_3641;
wire n_4577;
wire n_4854;
wire n_105;
wire n_4202;
wire n_5212;
wire n_5000;
wire n_2853;
wire n_1323;
wire n_688;
wire n_3766;
wire n_1353;
wire n_800;
wire n_2880;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_4165;
wire n_4866;
wire n_4038;
wire n_4109;
wire n_5297;
wire n_915;
wire n_864;
wire n_5420;
wire n_1264;
wire n_447;
wire n_4412;
wire n_3407;
wire n_3599;
wire n_3621;
wire n_1580;
wire n_5234;
wire n_2244;
wire n_3815;
wire n_2257;
wire n_497;
wire n_1607;
wire n_2538;
wire n_2105;
wire n_5259;
wire n_3163;
wire n_5440;
wire n_1118;
wire n_1686;
wire n_947;
wire n_373;
wire n_3710;
wire n_307;
wire n_4155;
wire n_1359;
wire n_2031;
wire n_3891;
wire n_1230;
wire n_4144;
wire n_375;
wire n_2165;
wire n_929;
wire n_3379;
wire n_4374;
wire n_3532;
wire n_1124;
wire n_5131;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1257;
wire n_1182;
wire n_3531;
wire n_2963;
wire n_3834;
wire n_4548;
wire n_3258;
wire n_4989;
wire n_4622;
wire n_1016;
wire n_4315;
wire n_2959;
wire n_2047;
wire n_1845;
wire n_240;
wire n_2193;
wire n_2478;
wire n_5140;
wire n_4816;
wire n_231;
wire n_1483;
wire n_2983;
wire n_227;
wire n_3810;
wire n_1289;
wire n_94;
wire n_2715;
wire n_5598;
wire n_2085;
wire n_1669;
wire n_370;
wire n_5306;
wire n_4483;
wire n_5342;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_2651;
wire n_4358;
wire n_5147;
wire n_3656;
wire n_2071;
wire n_2561;
wire n_2643;
wire n_1374;
wire n_4793;
wire n_4168;
wire n_3446;
wire n_955;
wire n_5511;
wire n_3028;
wire n_4806;
wire n_1146;
wire n_4350;
wire n_5533;
wire n_550;
wire n_897;
wire n_5280;
wire n_1428;
wire n_1216;
wire n_5235;
wire n_3836;
wire n_3963;
wire n_1872;
wire n_3389;
wire n_1931;
wire n_4187;
wire n_1070;
wire n_4166;
wire n_5206;
wire n_1030;
wire n_3222;
wire n_1071;
wire n_1267;
wire n_1801;
wire n_5419;
wire n_1513;
wire n_2970;
wire n_2235;
wire n_673;
wire n_837;
wire n_4937;
wire n_3980;
wire n_2791;
wire n_5103;
wire n_680;
wire n_1473;
wire n_3755;
wire n_4258;
wire n_4498;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_5285;
wire n_3563;
wire n_2506;
wire n_675;
wire n_4064;
wire n_4936;
wire n_5387;
wire n_1556;
wire n_184;
wire n_1863;
wire n_3841;
wire n_114;
wire n_2118;
wire n_4770;
wire n_2944;
wire n_881;
wire n_2407;
wire n_4907;
wire n_468;
wire n_5058;
wire n_129;
wire n_3262;
wire n_1450;
wire n_5018;
wire n_4006;
wire n_4861;
wire n_1322;
wire n_3690;
wire n_889;
wire n_2358;
wire n_973;
wire n_5192;
wire n_5141;
wire n_3716;
wire n_5133;
wire n_1700;
wire n_2833;
wire n_4712;
wire n_477;
wire n_3191;
wire n_3837;
wire n_3193;
wire n_1971;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_3544;
wire n_4310;
wire n_1523;
wire n_1950;
wire n_1447;
wire n_2370;
wire n_5159;
wire n_3954;
wire n_3025;
wire n_4674;
wire n_4908;
wire n_736;
wire n_5097;
wire n_2750;
wire n_3899;
wire n_1278;
wire n_4159;
wire n_3714;
wire n_3071;
wire n_3739;
wire n_593;
wire n_4069;
wire n_2784;
wire n_3718;
wire n_3470;
wire n_3092;
wire n_4862;
wire n_2557;
wire n_5300;
wire n_1248;
wire n_289;
wire n_4850;
wire n_3781;
wire n_4813;
wire n_4912;
wire n_2590;
wire n_2330;
wire n_2942;
wire n_5525;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_944;
wire n_3889;
wire n_4256;
wire n_4224;
wire n_3508;
wire n_4024;
wire n_2218;
wire n_2267;
wire n_857;
wire n_2636;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_5400;
wire n_2759;
wire n_4415;
wire n_5552;
wire n_4702;
wire n_4252;
wire n_4457;
wire n_971;
wire n_117;
wire n_404;
wire n_5139;
wire n_1393;
wire n_2319;
wire n_596;
wire n_3481;
wire n_5481;
wire n_2808;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_4491;
wire n_266;
wire n_2930;
wire n_1838;
wire n_3514;
wire n_2777;
wire n_2434;
wire n_4132;
wire n_2660;
wire n_2611;
wire n_4261;
wire n_1660;
wire n_4886;
wire n_4090;
wire n_2529;
wire n_2698;
wire n_5043;
wire n_1662;
wire n_1481;
wire n_4001;
wire n_3047;
wire n_868;
wire n_2454;
wire n_4371;
wire n_914;
wire n_5281;
wire n_4473;
wire n_3120;
wire n_4007;
wire n_1743;
wire n_4268;
wire n_5048;
wire n_5521;
wire n_5028;
wire n_1479;
wire n_4480;
wire n_2350;
wire n_3895;
wire n_4194;
wire n_759;
wire n_5585;
wire n_4824;
wire n_1892;
wire n_4120;
wire n_4427;
wire n_3745;
wire n_806;
wire n_2990;
wire n_1766;
wire n_324;
wire n_1571;
wire n_3119;
wire n_4142;
wire n_1189;
wire n_4082;
wire n_5561;
wire n_3479;
wire n_4085;
wire n_4073;
wire n_4260;
wire n_1649;
wire n_4163;
wire n_4439;
wire n_2064;
wire n_3867;
wire n_4372;
wire n_3500;
wire n_3279;
wire n_2621;
wire n_5073;
wire n_5024;
wire n_523;
wire n_1537;
wire n_4262;
wire n_2671;
wire n_1798;
wire n_1790;
wire n_4720;
wire n_525;
wire n_1647;
wire n_4685;
wire n_2563;
wire n_2387;
wire n_4334;
wire n_1674;
wire n_1830;
wire n_2073;
wire n_4511;
wire n_5515;
wire n_139;
wire n_4014;
wire n_5250;
wire n_3144;
wire n_4757;
wire n_2913;
wire n_2336;
wire n_254;
wire n_1233;
wire n_5607;
wire n_1615;
wire n_4175;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_244;
wire n_4648;
wire n_1333;
wire n_5006;
wire n_1443;
wire n_946;
wire n_1539;
wire n_4892;
wire n_3823;
wire n_1866;
wire n_4173;
wire n_689;
wire n_738;
wire n_1624;
wire n_4970;
wire n_640;
wire n_3816;
wire n_1279;
wire n_5404;
wire n_4108;
wire n_4486;
wire n_610;
wire n_2960;
wire n_1090;
wire n_5438;
wire n_633;
wire n_439;
wire n_4627;
wire n_758;
wire n_2290;
wire n_2045;
wire n_3369;
wire n_3783;
wire n_2040;
wire n_3199;
wire n_3843;
wire n_1049;
wire n_2145;
wire n_1639;
wire n_1068;
wire n_3030;
wire n_2580;
wire n_3685;
wire n_4249;
wire n_122;
wire n_331;
wire n_5163;
wire n_2039;
wire n_4961;
wire n_90;
wire n_3753;
wire n_2035;
wire n_4718;
wire n_3555;
wire n_3579;
wire n_5190;
wire n_2509;
wire n_3236;
wire n_4317;
wire n_1362;
wire n_4855;
wire n_3969;
wire n_2459;
wire n_4154;
wire n_152;
wire n_3396;
wire n_1445;
wire n_4023;
wire n_4420;
wire n_1923;
wire n_5138;
wire n_1017;
wire n_5374;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1828;
wire n_2320;
wire n_1045;
wire n_5349;
wire n_2038;
wire n_2137;
wire n_4973;
wire n_4640;
wire n_2583;
wire n_484;
wire n_1033;
wire n_4396;
wire n_5127;
wire n_636;
wire n_4367;
wire n_2087;
wire n_5485;
wire n_5216;
wire n_1009;
wire n_109;
wire n_454;
wire n_1989;
wire n_3818;
wire n_2523;
wire n_255;
wire n_4387;
wire n_4951;
wire n_4453;
wire n_4170;
wire n_1578;
wire n_3719;
wire n_1959;
wire n_3681;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_4308;
wire n_2812;
wire n_473;
wire n_2355;
wire n_2133;
wire n_1426;
wire n_3830;
wire n_2585;
wire n_2725;
wire n_614;
wire n_5175;
wire n_3883;
wire n_1355;
wire n_2565;
wire n_4152;
wire n_773;
wire n_208;
wire n_142;
wire n_743;
wire n_4392;
wire n_4660;
wire n_3149;
wire n_5611;
wire n_296;
wire n_3268;
wire n_4281;
wire n_4661;
wire n_4200;
wire n_3614;
wire n_2111;
wire n_3301;
wire n_3466;
wire n_4962;
wire n_1237;
wire n_2595;
wire n_761;
wire n_3411;
wire n_4958;
wire n_329;
wire n_4271;
wire n_5171;
wire n_3586;
wire n_1390;
wire n_5554;
wire n_4071;
wire n_4921;
wire n_130;
wire n_1980;
wire n_5427;
wire n_3065;
wire n_4361;
wire n_1093;
wire n_5417;
wire n_263;
wire n_4614;
wire n_1265;
wire n_224;
wire n_2681;
wire n_3103;
wire n_765;
wire n_4945;
wire n_2424;
wire n_4922;
wire n_4732;
wire n_1015;
wire n_1651;
wire n_2775;
wire n_4693;
wire n_5488;
wire n_511;
wire n_358;
wire n_1101;
wire n_1106;
wire n_4326;
wire n_3557;
wire n_2230;
wire n_5447;
wire n_5383;
wire n_4744;
wire n_2851;
wire n_4305;
wire n_174;
wire n_1455;
wire n_767;
wire n_2490;
wire n_1407;
wire n_441;
wire n_4213;
wire n_2849;
wire n_3692;
wire n_2204;
wire n_365;
wire n_4929;
wire n_729;
wire n_1961;
wire n_4964;
wire n_911;
wire n_1430;
wire n_4802;
wire n_513;
wire n_1354;
wire n_4139;
wire n_1044;
wire n_3029;
wire n_2508;
wire n_4031;
wire n_2416;
wire n_5437;
wire n_623;
wire n_3881;
wire n_2461;
wire n_490;
wire n_2243;
wire n_4583;
wire n_233;
wire n_572;
wire n_4210;
wire n_5245;
wire n_4666;
wire n_2929;
wire n_3751;
wire n_2555;
wire n_2662;
wire n_1611;
wire n_2368;
wire n_2890;
wire n_2554;
wire n_3927;
wire n_3698;
wire n_1082;
wire n_1840;
wire n_4540;
wire n_3961;
wire n_716;
wire n_1630;
wire n_4891;
wire n_391;
wire n_701;
wire n_1023;
wire n_5603;
wire n_539;
wire n_803;
wire n_1092;
wire n_3559;
wire n_2661;
wire n_2572;
wire n_3993;
wire n_4940;
wire n_5208;
wire n_1056;
wire n_3588;
wire n_2308;
wire n_4590;
wire n_5606;
wire n_4830;
wire n_5231;
wire n_5237;
wire n_4664;
wire n_3860;
wire n_1029;
wire n_1206;
wire n_5456;
wire n_3160;
wire n_2191;
wire n_5093;
wire n_2428;
wire n_3847;
wire n_4946;
wire n_1346;
wire n_4906;
wire n_2158;
wire n_3290;
wire n_4663;
wire n_5390;
wire n_1060;
wire n_5347;
wire n_2824;
wire n_3033;
wire n_3298;
wire n_248;
wire n_2440;
wire n_4883;
wire n_1386;
wire n_2923;
wire n_1442;
wire n_4162;
wire n_3665;
wire n_5115;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_483;
wire n_4297;
wire n_1632;
wire n_1085;
wire n_1066;
wire n_3800;
wire n_2403;
wire n_5407;
wire n_4608;
wire n_5232;
wire n_2792;
wire n_2870;
wire n_3991;
wire n_378;
wire n_1112;
wire n_3134;
wire n_4172;
wire n_4791;
wire n_4536;
wire n_5149;
wire n_2463;
wire n_5151;
wire n_4773;
wire n_5345;
wire n_5357;
wire n_4497;
wire n_2472;
wire n_4611;
wire n_4755;
wire n_1768;
wire n_2294;
wire n_4960;
wire n_455;
wire n_2993;
wire n_1719;
wire n_3864;
wire n_385;
wire n_4658;
wire n_5135;
wire n_2732;
wire n_2309;
wire n_2948;
wire n_1560;
wire n_5494;
wire n_4362;
wire n_4306;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_4422;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_3482;
wire n_2233;
wire n_1312;
wire n_804;
wire n_537;
wire n_4555;
wire n_2827;
wire n_5136;
wire n_5228;
wire n_153;
wire n_1504;
wire n_3956;
wire n_5323;
wire n_3572;
wire n_250;
wire n_992;
wire n_4215;
wire n_4280;
wire n_3375;
wire n_4047;
wire n_260;
wire n_5471;
wire n_842;
wire n_5434;
wire n_2082;
wire n_1643;
wire n_3167;
wire n_5558;
wire n_5350;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_5338;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3854;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3078;
wire n_540;
wire n_323;
wire n_894;
wire n_3253;
wire n_4027;
wire n_831;
wire n_2280;
wire n_4599;
wire n_3363;
wire n_4812;
wire n_1511;
wire n_234;
wire n_3689;
wire n_2020;
wire n_4628;
wire n_1881;
wire n_988;
wire n_2749;
wire n_3451;
wire n_4873;
wire n_5588;
wire n_4657;
wire n_2971;
wire n_2311;
wire n_3950;
wire n_4458;
wire n_4121;
wire n_1616;
wire n_5090;
wire n_4476;
wire n_5613;
wire n_2298;
wire n_4756;
wire n_3869;
wire n_4307;
wire n_5104;
wire n_5042;
wire n_4860;
wire n_4359;
wire n_635;
wire n_2303;
wire n_2810;
wire n_2747;
wire n_1848;
wire n_5571;
wire n_2126;
wire n_4573;
wire n_5289;
wire n_4118;
wire n_5513;
wire n_4803;
wire n_4079;
wire n_4091;
wire n_681;
wire n_1638;
wire n_2002;
wire n_5145;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_5132;
wire n_830;
wire n_5191;
wire n_3085;
wire n_1655;
wire n_749;
wire n_5359;
wire n_2574;
wire n_1134;
wire n_5293;
wire n_1358;
wire n_717;
wire n_4316;
wire n_939;
wire n_3697;
wire n_482;
wire n_1232;
wire n_734;
wire n_2638;
wire n_4044;
wire n_4062;
wire n_4524;
wire n_4843;
wire n_3971;
wire n_1338;
wire n_5510;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_2711;
wire n_5363;
wire n_5200;
wire n_338;
wire n_1653;
wire n_1506;
wire n_5618;
wire n_990;
wire n_2867;
wire n_1894;
wire n_975;
wire n_2794;
wire n_567;
wire n_3145;
wire n_3124;
wire n_4253;
wire n_5356;
wire n_151;
wire n_5369;
wire n_2608;
wire n_5258;
wire n_2657;
wire n_770;
wire n_5255;
wire n_2852;
wire n_2392;
wire n_711;
wire n_3517;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_1834;
wire n_3758;
wire n_3356;
wire n_2835;
wire n_617;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_5080;
wire n_1516;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_2409;
wire n_3402;
wire n_5295;
wire n_217;
wire n_4679;
wire n_4115;
wire n_726;
wire n_4998;
wire n_2988;
wire n_1731;
wire n_818;
wire n_1970;
wire n_2766;
wire n_2201;
wire n_2117;
wire n_4167;
wire n_1993;
wire n_5155;
wire n_3835;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_3967;
wire n_5016;
wire n_1912;
wire n_3401;
wire n_3226;
wire n_1410;
wire n_707;
wire n_3902;
wire n_4730;
wire n_937;
wire n_2779;
wire n_1584;
wire n_487;
wire n_3654;
wire n_2164;
wire n_2115;
wire n_2232;
wire n_5327;
wire n_1302;
wire n_1774;
wire n_4713;
wire n_5137;
wire n_2811;
wire n_3348;
wire n_179;
wire n_410;
wire n_895;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_4204;
wire n_5098;
wire n_1543;
wire n_1991;
wire n_2224;
wire n_732;
wire n_4743;
wire n_500;
wire n_1067;
wire n_3805;
wire n_3825;
wire n_148;
wire n_3657;
wire n_4924;
wire n_3928;
wire n_4859;
wire n_2692;
wire n_538;
wire n_2008;
wire n_4654;
wire n_5423;
wire n_799;
wire n_1213;
wire n_4733;
wire n_3792;
wire n_4272;
wire n_3974;
wire n_3871;
wire n_1753;
wire n_2283;
wire n_3278;
wire n_89;
wire n_1689;
wire n_4269;
wire n_4695;
wire n_1855;
wire n_869;
wire n_401;
wire n_3312;
wire n_1352;
wire n_2197;
wire n_2199;
wire n_5069;
wire n_3285;
wire n_137;
wire n_294;
wire n_3968;
wire n_5099;
wire n_2228;
wire n_4704;
wire n_4551;
wire n_5052;
wire n_684;
wire n_124;
wire n_268;
wire n_2421;
wire n_2902;
wire n_4957;
wire n_664;
wire n_2480;
wire n_235;
wire n_2363;
wire n_643;
wire n_4072;
wire n_916;
wire n_5579;
wire n_1115;
wire n_4781;
wire n_3606;
wire n_5004;
wire n_2550;
wire n_467;
wire n_4424;
wire n_823;
wire n_725;
wire n_3055;
wire n_3711;
wire n_3315;
wire n_3172;
wire n_3292;
wire n_4436;
wire n_3878;
wire n_4450;
wire n_3553;
wire n_719;
wire n_4746;
wire n_1683;
wire n_1530;
wire n_997;
wire n_932;
wire n_3131;
wire n_5118;
wire n_5105;
wire n_1409;
wire n_3850;
wire n_788;
wire n_4459;
wire n_1268;
wire n_2996;
wire n_559;
wire n_5591;
wire n_508;
wire n_1320;
wire n_4050;
wire n_986;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_2102;
wire n_5623;
wire n_1063;
wire n_4853;
wire n_981;
wire n_867;
wire n_2422;
wire n_134;
wire n_2239;
wire n_5256;
wire n_587;
wire n_2950;
wire n_5220;
wire n_3852;
wire n_548;
wire n_5178;
wire n_812;
wire n_4520;
wire n_518;
wire n_2057;
wire n_4008;
wire n_5507;
wire n_905;
wire n_5077;
wire n_782;
wire n_3858;
wire n_1901;
wire n_4502;
wire n_3032;
wire n_4851;
wire n_1330;
wire n_3072;
wire n_3313;
wire n_3081;
wire n_2710;
wire n_1745;
wire n_3924;
wire n_769;
wire n_4571;
wire n_2006;
wire n_934;
wire n_5314;
wire n_1618;
wire n_826;
wire n_2343;
wire n_3439;
wire n_5049;
wire n_654;
wire n_2535;
wire n_4205;
wire n_2726;
wire n_570;
wire n_5277;
wire n_4723;
wire n_5176;
wire n_2799;
wire n_4454;
wire n_4229;
wire n_1083;
wire n_4739;
wire n_2376;
wire n_5483;
wire n_3017;
wire n_787;
wire n_2456;
wire n_3904;
wire n_5150;
wire n_2678;
wire n_95;
wire n_4838;
wire n_2872;
wire n_2451;
wire n_5075;
wire n_522;
wire n_4879;
wire n_5051;
wire n_930;
wire n_181;
wire n_3926;
wire n_1962;
wire n_3996;
wire n_4221;
wire n_1577;
wire n_2854;
wire n_386;
wire n_1701;
wire n_4181;
wire n_1550;
wire n_2764;
wire n_1498;
wire n_4225;
wire n_682;
wire n_141;
wire n_2567;
wire n_5142;
wire n_3102;
wire n_922;
wire n_1648;
wire n_4153;
wire n_5156;
wire n_3627;
wire n_4300;
wire n_3551;
wire n_432;
wire n_1769;
wire n_4783;
wire n_839;
wire n_2964;
wire n_3769;
wire n_2673;
wire n_4530;
wire n_4267;
wire n_140;
wire n_2292;
wire n_3865;
wire n_3859;
wire n_3722;
wire n_2442;
wire n_928;
wire n_1943;
wire n_3117;
wire n_3428;
wire n_2961;
wire n_3351;
wire n_3527;
wire n_236;
wire n_1396;
wire n_1348;
wire n_2883;
wire n_1752;
wire n_4182;
wire n_2912;
wire n_1315;
wire n_4825;
wire n_4440;
wire n_4549;
wire n_1910;
wire n_3955;
wire n_462;
wire n_5120;
wire n_5470;
wire n_4565;
wire n_4039;
wire n_3227;
wire n_3300;
wire n_4303;
wire n_4574;
wire n_471;
wire n_4839;
wire n_5222;
wire n_1028;
wire n_4016;
wire n_474;
wire n_3435;
wire n_3575;
wire n_1546;
wire n_595;
wire n_632;
wire n_4231;
wire n_3165;
wire n_4923;
wire n_3652;
wire n_4097;
wire n_170;
wire n_161;
wire n_4083;
wire n_1937;
wire n_4461;
wire n_3234;
wire n_5392;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3916;
wire n_2569;
wire n_3556;
wire n_4101;
wire n_2196;
wire n_3591;
wire n_4273;
wire n_3024;
wire n_5443;
wire n_3512;
wire n_5600;
wire n_4939;
wire n_5169;
wire n_4389;
wire n_3930;
wire n_4448;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_2503;
wire n_1540;
wire n_1936;
wire n_5502;
wire n_2027;
wire n_5568;
wire n_453;
wire n_403;
wire n_2642;
wire n_720;
wire n_2500;
wire n_1918;
wire n_863;
wire n_4831;
wire n_2513;
wire n_2695;
wire n_3480;
wire n_3057;
wire n_3194;
wire n_2414;
wire n_1402;
wire n_3662;
wire n_4319;
wire n_5474;
wire n_644;
wire n_2229;
wire n_1397;
wire n_4596;
wire n_5413;
wire n_2004;
wire n_5412;
wire n_251;
wire n_3694;
wire n_2586;
wire n_4726;
wire n_1398;
wire n_1879;
wire n_4751;
wire n_4222;
wire n_1196;
wire n_2274;
wire n_2972;
wire n_3225;
wire n_811;
wire n_334;
wire n_175;
wire n_4119;
wire n_3799;
wire n_4298;
wire n_5201;
wire n_4474;
wire n_1089;
wire n_5217;
wire n_1004;
wire n_242;
wire n_2511;
wire n_1681;
wire n_3383;
wire n_3585;
wire n_2975;
wire n_5490;
wire n_438;
wire n_5029;
wire n_2704;
wire n_4214;
wire n_5158;
wire n_4884;
wire n_533;
wire n_4366;
wire n_1251;
wire n_4009;
wire n_278;
wire n_4580;
wire n_1263;
wire n_611;
wire n_1126;
wire n_4129;
wire n_4871;
wire n_2617;
wire n_4999;
wire n_1859;
wire n_1677;
wire n_5557;
wire n_5472;
wire n_2955;
wire n_4112;
wire n_4337;
wire n_4138;
wire n_5396;
wire n_552;
wire n_1528;
wire n_5335;
wire n_1292;
wire n_2520;
wire n_1198;
wire n_956;
wire n_423;
wire n_2134;
wire n_4236;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_5002;
wire n_3595;
wire n_1347;
wire n_5143;
wire n_4238;
wire n_1451;
wire n_1022;
wire n_1545;
wire n_2374;
wire n_173;
wire n_859;
wire n_1947;
wire n_2114;
wire n_3571;
wire n_854;
wire n_1799;
wire n_2396;
wire n_4734;
wire n_674;
wire n_1939;
wire n_2486;
wire n_516;
wire n_4635;
wire n_1152;
wire n_3501;
wire n_1869;
wire n_4013;
wire n_606;
wire n_3039;
wire n_275;
wire n_2011;
wire n_4242;
wire n_4984;
wire n_3851;
wire n_2543;
wire n_150;
wire n_3036;
wire n_1896;
wire n_3180;
wire n_5283;
wire n_5268;
wire n_191;
wire n_1705;
wire n_659;
wire n_4561;
wire n_2639;
wire n_3325;
wire n_3107;
wire n_4021;
wire n_3880;
wire n_5122;
wire n_1261;
wire n_938;
wire n_3186;
wire n_4955;
wire n_1154;
wire n_5556;
wire n_5462;
wire n_4501;
wire n_3696;
wire n_406;
wire n_546;
wire n_1280;
wire n_3650;
wire n_291;
wire n_2761;
wire n_257;
wire n_3157;
wire n_709;
wire n_2537;
wire n_2144;
wire n_920;
wire n_2515;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_5330;
wire n_4197;
wire n_4829;
wire n_976;
wire n_1949;
wire n_1946;
wire n_2936;
wire n_775;
wire n_1484;
wire n_1328;
wire n_4715;
wire n_5039;
wire n_2141;
wire n_4369;
wire n_5378;
wire n_4543;
wire n_2099;
wire n_4941;
wire n_5542;
wire n_1831;
wire n_1598;
wire n_4394;
wire n_1850;
wire n_163;
wire n_243;
wire n_5519;
wire n_1749;
wire n_3101;
wire n_3669;
wire n_215;
wire n_350;
wire n_196;
wire n_5278;
wire n_2663;
wire n_1394;
wire n_5586;
wire n_580;
wire n_2693;
wire n_4065;
wire n_3798;
wire n_5187;
wire n_4944;
wire n_926;
wire n_2249;
wire n_2180;
wire n_4135;
wire n_1218;
wire n_2632;
wire n_475;
wire n_1547;
wire n_777;
wire n_1755;
wire n_415;
wire n_485;
wire n_958;
wire n_2908;
wire n_3744;
wire n_4263;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_3291;
wire n_4716;
wire n_4942;
wire n_164;
wire n_2432;
wire n_1521;
wire n_3405;
wire n_214;
wire n_4745;
wire n_2337;
wire n_1167;
wire n_1384;
wire n_3907;
wire n_5344;
wire n_923;
wire n_4629;
wire n_213;
wire n_2932;
wire n_2980;
wire n_464;
wire n_5225;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_4857;
wire n_3136;
wire n_4080;
wire n_4226;
wire n_4741;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_4752;
wire n_5265;
wire n_1750;
wire n_1459;
wire n_460;
wire n_3986;
wire n_4376;
wire n_4753;
wire n_571;
wire n_4552;
wire n_3885;
wire n_2713;
wire n_5196;
wire n_5181;
wire n_2644;
wire n_1197;
wire n_2951;
wire n_3008;
wire n_3709;
wire n_5574;
wire n_5126;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_3427;
wire n_4067;
wire n_1403;
wire n_5553;
wire n_4176;
wire n_4042;
wire n_4385;
wire n_3320;
wire n_5009;
wire n_2688;
wire n_5368;
wire n_1202;
wire n_1463;
wire n_3651;
wire n_4333;
wire n_3359;
wire n_2865;
wire n_349;
wire n_2706;
wire n_5499;
wire n_3676;
wire n_4375;
wire n_4788;
wire n_4717;
wire n_4986;
wire n_5604;
wire n_3789;
wire n_2152;
wire n_3598;
wire n_627;
wire n_4815;
wire n_4246;
wire n_3580;
wire n_2139;
wire n_4609;
wire n_5291;
wire n_5114;
wire n_91;
wire n_2674;
wire n_1565;
wire n_4088;
wire n_3682;
wire n_4357;
wire n_3371;
wire n_1809;
wire n_4462;
wire n_4472;
wire n_647;
wire n_3433;
wire n_1072;
wire n_5288;
wire n_2305;
wire n_5540;
wire n_2450;
wire n_561;
wire n_3447;
wire n_3305;
wire n_4151;
wire n_4148;
wire n_1712;
wire n_3528;
wire n_4373;
wire n_4934;
wire n_5218;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_4630;
wire n_5408;
wire n_4643;
wire n_4331;
wire n_3989;
wire n_4475;
wire n_4846;
wire n_3804;
wire n_4344;
wire n_1775;
wire n_3296;
wire n_1368;
wire n_2762;
wire n_4683;
wire n_5366;
wire n_728;
wire n_1162;
wire n_272;
wire n_1847;
wire n_2767;
wire n_2603;
wire n_3116;
wire n_1884;
wire n_3602;
wire n_2967;
wire n_409;
wire n_887;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_2195;
wire n_5477;
wire n_300;
wire n_5451;
wire n_3923;
wire n_931;
wire n_599;
wire n_4696;
wire n_2626;
wire n_3441;
wire n_1978;
wire n_1544;
wire n_639;
wire n_5086;
wire n_1629;
wire n_2801;
wire n_4011;
wire n_4905;
wire n_121;
wire n_2763;
wire n_360;
wire n_2825;
wire n_3643;
wire n_4876;
wire n_1997;
wire n_3748;
wire n_1477;
wire n_3142;
wire n_4278;
wire n_1635;
wire n_4623;
wire n_187;
wire n_4910;
wire n_2690;
wire n_4410;
wire n_3370;
wire n_2215;
wire n_5053;
wire n_1259;
wire n_4553;
wire n_706;
wire n_746;
wire n_784;
wire n_3978;
wire n_110;
wire n_4809;
wire n_5226;
wire n_1244;
wire n_1925;
wire n_3660;
wire n_1815;
wire n_1788;
wire n_2491;
wire n_5079;
wire n_5590;
wire n_913;
wire n_3833;
wire n_865;
wire n_697;
wire n_1222;
wire n_1679;
wire n_4841;
wire n_776;
wire n_2022;
wire n_3814;
wire n_1415;
wire n_2592;
wire n_2838;
wire n_4842;
wire n_4911;
wire n_4340;
wire n_3513;
wire n_3133;
wire n_4645;
wire n_1191;
wire n_2992;
wire n_3725;
wire n_1833;
wire n_4920;
wire n_4972;
wire n_2517;
wire n_284;
wire n_3128;
wire n_5426;
wire n_744;
wire n_629;
wire n_2631;
wire n_2178;
wire n_1767;
wire n_1529;
wire n_2469;
wire n_3355;
wire n_604;
wire n_2007;
wire n_3917;
wire n_3942;
wire n_2736;
wire n_3765;
wire n_498;
wire n_5531;
wire n_3000;
wire n_252;
wire n_624;
wire n_5429;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_3108;
wire n_3111;
wire n_1839;
wire n_1837;
wire n_4557;
wire n_5248;
wire n_4451;
wire n_2875;
wire n_936;
wire n_1500;
wire n_3844;
wire n_3280;
wire n_4054;
wire n_5448;
wire n_3471;
wire n_5432;
wire n_259;
wire n_448;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_5160;
wire n_2741;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_1656;
wire n_3564;
wire n_1158;
wire n_3988;
wire n_563;
wire n_3457;
wire n_204;
wire n_1678;
wire n_4324;
wire n_4821;
wire n_1871;
wire n_5445;
wire n_3630;
wire n_3271;
wire n_4771;
wire n_908;
wire n_4086;
wire n_2412;
wire n_4814;
wire n_724;
wire n_2084;
wire n_1781;
wire n_3648;
wire n_3075;
wire n_3173;
wire n_5332;
wire n_5108;
wire n_4692;
wire n_456;
wire n_959;
wire n_3031;
wire n_3701;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_2666;
wire n_3385;
wire n_2171;
wire n_4708;
wire n_2768;
wire n_2314;
wire n_4826;
wire n_2420;
wire n_3343;
wire n_514;
wire n_1079;
wire n_5489;
wire n_1593;
wire n_3767;
wire n_442;
wire n_2299;
wire n_131;
wire n_2540;
wire n_2873;
wire n_4589;
wire n_5057;
wire n_4578;
wire n_1640;
wire n_2162;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_3221;
wire n_742;
wire n_750;
wire n_5436;
wire n_2168;
wire n_2790;
wire n_5072;
wire n_3629;
wire n_3021;
wire n_185;
wire n_2359;
wire n_3674;
wire n_5286;
wire n_3502;
wire n_3098;
wire n_1383;
wire n_5013;
wire n_2312;
wire n_3015;
wire n_1171;
wire n_1920;
wire n_1065;
wire n_5569;
wire n_5439;
wire n_5619;
wire n_4147;
wire n_2048;
wire n_3607;
wire n_4925;
wire n_1921;
wire n_1309;
wire n_4974;
wire n_355;
wire n_1800;
wire n_1548;
wire n_4932;
wire n_1421;
wire n_4510;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_3787;
wire n_5119;
wire n_2124;
wire n_613;
wire n_1119;
wire n_1240;
wire n_3827;
wire n_829;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_4447;
wire n_4285;
wire n_4651;
wire n_361;
wire n_700;
wire n_573;
wire n_4818;
wire n_4514;
wire n_388;
wire n_1366;
wire n_4800;
wire n_3960;
wire n_3248;
wire n_2277;
wire n_1568;
wire n_2110;
wire n_274;
wire n_582;
wire n_1332;
wire n_4433;
wire n_2879;
wire n_2474;
wire n_2090;
wire n_3153;
wire n_512;
wire n_1591;
wire n_2033;
wire n_4341;
wire n_1682;
wire n_4312;
wire n_2628;
wire n_3399;
wire n_1249;
wire n_1111;
wire n_2132;
wire n_2400;
wire n_4633;
wire n_609;
wire n_3838;
wire n_1909;
wire n_4277;
wire n_112;
wire n_4140;
wire n_3675;
wire n_5092;
wire n_1140;
wire n_891;
wire n_3387;
wire n_5186;
wire n_4662;
wire n_3779;
wire n_2464;
wire n_2831;
wire n_102;
wire n_1456;
wire n_4882;
wire n_4993;
wire n_2365;
wire n_4832;
wire n_4207;
wire n_987;
wire n_4545;
wire n_3037;
wire n_261;
wire n_4868;
wire n_1885;
wire n_2452;
wire n_3925;
wire n_2176;
wire n_1816;
wire n_5238;
wire n_4059;
wire n_2455;
wire n_4595;
wire n_1849;
wire n_1131;
wire n_5054;
wire n_2467;
wire n_1094;
wire n_2288;
wire n_4063;
wire n_5399;
wire n_346;
wire n_1209;
wire n_3592;
wire n_4650;
wire n_602;
wire n_4888;
wire n_5326;
wire n_1435;
wire n_879;
wire n_3394;
wire n_4874;
wire n_3793;
wire n_4669;
wire n_405;
wire n_4339;
wire n_1645;
wire n_4041;
wire n_5459;
wire n_2858;
wire n_4060;
wire n_996;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_2128;
wire n_5528;
wire n_3097;
wire n_5391;
wire n_120;
wire n_327;
wire n_135;
wire n_4541;
wire n_5422;
wire n_3824;
wire n_3388;
wire n_5267;
wire n_4494;
wire n_3059;
wire n_5523;
wire n_3465;
wire n_1316;
wire n_4796;
wire n_1438;
wire n_3589;
wire n_952;
wire n_2534;
wire n_1229;
wire n_4799;
wire n_5153;
wire n_3449;
wire n_2694;
wire n_2198;
wire n_2610;
wire n_2989;
wire n_2789;
wire n_4775;
wire n_2216;
wire n_531;
wire n_5044;
wire n_1897;
wire n_764;
wire n_1424;
wire n_162;
wire n_5365;
wire n_2933;
wire n_5045;
wire n_4381;
wire n_4266;
wire n_3886;
wire n_5354;
wire n_4455;
wire n_2328;
wire n_199;
wire n_4248;
wire n_5452;
wire n_4754;
wire n_4554;
wire n_5595;
wire n_4845;
wire n_3053;
wire n_1299;
wire n_3893;
wire n_1141;
wire n_2465;
wire n_3548;
wire n_4585;
wire n_418;
wire n_315;
wire n_451;
wire n_1699;
wire n_3334;
wire n_2541;
wire n_4383;
wire n_1139;
wire n_397;
wire n_5535;
wire n_1432;
wire n_3875;
wire n_5370;
wire n_4003;
wire n_5372;
wire n_5299;
wire n_2402;
wire n_5594;
wire n_4301;
wire n_1050;
wire n_841;
wire n_4586;
wire n_1954;
wire n_4048;
wire n_1844;
wire n_3777;
wire n_4784;
wire n_2999;
wire n_1644;
wire n_5550;
wire n_5082;
wire n_4046;
wire n_1974;
wire n_2086;
wire n_5209;
wire n_3537;
wire n_3080;
wire n_4199;
wire n_2701;
wire n_3362;
wire n_1631;
wire n_5559;
wire n_3105;
wire n_5478;
wire n_1179;
wire n_753;
wire n_1048;
wire n_4286;
wire n_5102;
wire n_2556;
wire n_2269;
wire n_3274;
wire n_3041;
wire n_4470;
wire n_2236;
wire n_330;
wire n_2816;
wire n_692;
wire n_820;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_4058;
wire n_3664;
wire n_4188;
wire n_1668;
wire n_3913;
wire n_3417;
wire n_1143;
wire n_1579;
wire n_4034;
wire n_1688;
wire n_492;
wire n_3327;
wire n_5275;
wire n_4689;
wire n_341;
wire n_5071;
wire n_3067;
wire n_2755;
wire n_543;
wire n_3237;
wire n_1992;
wire n_4402;
wire n_4239;
wire n_3400;
wire n_449;
wire n_4550;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3382;
wire n_3574;
wire n_5227;
wire n_2169;
wire n_1557;
wire n_4201;
wire n_618;
wire n_896;
wire n_3316;
wire n_5242;
wire n_356;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1730;
wire n_3603;
wire n_4123;
wire n_2192;
wire n_5520;
wire n_964;
wire n_3633;
wire n_4479;
wire n_1373;
wire n_2670;
wire n_1646;
wire n_1307;
wire n_4416;
wire n_3372;
wire n_4539;
wire n_814;
wire n_2707;
wire n_2471;
wire n_1472;
wire n_1671;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_4682;
wire n_5353;
wire n_3708;
wire n_5294;
wire n_1204;
wire n_3729;
wire n_4978;
wire n_4690;
wire n_4437;
wire n_5458;
wire n_3861;
wire n_5617;
wire n_4736;
wire n_3780;
wire n_783;
wire n_1928;
wire n_5244;
wire n_5382;
wire n_1188;
wire n_3957;
wire n_5274;
wire n_3848;
wire n_4284;
wire n_2600;
wire n_3919;
wire n_336;
wire n_5384;
wire n_3608;
wire n_510;
wire n_216;
wire n_4513;
wire n_3233;
wire n_3829;
wire n_3177;
wire n_4053;
wire n_2352;
wire n_5125;
wire n_4040;
wire n_2207;
wire n_5587;
wire n_2619;
wire n_2444;
wire n_241;
wire n_1110;
wire n_3123;
wire n_5056;
wire n_1088;
wire n_5249;
wire n_3393;
wire n_638;
wire n_866;
wire n_5198;
wire n_5360;
wire n_5233;
wire n_4887;
wire n_4617;
wire n_5269;
wire n_3520;
wire n_2492;
wire n_249;
wire n_577;
wire n_4005;
wire n_1687;
wire n_1637;
wire n_4904;
wire n_1419;
wire n_693;
wire n_4792;
wire n_3578;
wire n_3812;
wire n_1886;
wire n_1389;
wire n_1256;
wire n_4980;
wire n_1465;
wire n_4290;
wire n_5247;
wire n_306;
wire n_1375;
wire n_3727;
wire n_5317;
wire n_3774;
wire n_3093;
wire n_1843;
wire n_3061;
wire n_1597;
wire n_1659;
wire n_2431;
wire n_1371;
wire n_4956;
wire n_5380;
wire n_2206;
wire n_3182;
wire n_2564;
wire n_4947;
wire n_876;
wire n_4656;
wire n_1190;
wire n_3896;
wire n_3958;
wire n_3450;
wire n_966;
wire n_4729;
wire n_4987;
wire n_5182;
wire n_4971;
wire n_1116;
wire n_2000;
wire n_1212;
wire n_2074;
wire n_206;
wire n_3174;
wire n_982;
wire n_1453;
wire n_2217;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_3408;
wire n_899;
wire n_2722;
wire n_5388;
wire n_2640;
wire n_4823;
wire n_4875;
wire n_1628;
wire n_3432;
wire n_1514;
wire n_1771;
wire n_557;
wire n_1005;
wire n_607;
wire n_679;
wire n_710;
wire n_3090;
wire n_527;
wire n_1168;
wire n_2437;
wire n_3762;
wire n_5564;
wire n_2445;
wire n_1427;
wire n_108;
wire n_1835;
wire n_177;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_4137;
wire n_2634;
wire n_4529;
wire n_910;
wire n_4323;
wire n_3034;
wire n_2212;
wire n_3972;
wire n_125;
wire n_529;
wire n_5539;
wire n_126;
wire n_202;
wire n_3308;
wire n_791;
wire n_1533;
wire n_5036;
wire n_5547;
wire n_4772;
wire n_3467;
wire n_4322;
wire n_1720;
wire n_2830;
wire n_4354;
wire n_159;
wire n_4653;
wire n_2354;
wire n_2246;
wire n_5273;
wire n_4677;
wire n_3901;
wire n_715;
wire n_1480;
wire n_5261;
wire n_3757;
wire n_3381;
wire n_5193;
wire n_1782;
wire n_2245;
wire n_4909;
wire n_1524;
wire n_1485;
wire n_115;
wire n_810;
wire n_2965;
wire n_416;
wire n_3635;
wire n_5022;
wire n_5005;
wire n_1144;
wire n_2814;
wire n_1570;
wire n_3882;
wire n_3046;
wire n_1170;
wire n_305;
wire n_2213;
wire n_3826;
wire n_3211;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_4634;
wire n_3337;
wire n_2527;
wire n_855;
wire n_5534;
wire n_1461;
wire n_3204;
wire n_2136;
wire n_5174;
wire n_1273;
wire n_1822;
wire n_4952;
wire n_5157;
wire n_3005;
wire n_1235;
wire n_4380;
wire n_980;
wire n_698;
wire n_3129;
wire n_4126;
wire n_1282;
wire n_1783;
wire n_2601;
wire n_5087;
wire n_3043;
wire n_998;
wire n_3802;
wire n_2375;
wire n_4506;
wire n_4880;
wire n_1907;
wire n_501;
wire n_2686;
wire n_2344;
wire n_3892;
wire n_4896;
wire n_5620;
wire n_1417;
wire n_1295;
wire n_5061;
wire n_5572;
wire n_1985;
wire n_2107;
wire n_3219;
wire n_2906;
wire n_4943;
wire n_382;
wire n_2187;
wire n_1762;
wire n_1013;
wire n_718;
wire n_3023;
wire n_4193;
wire n_4075;
wire n_3104;
wire n_612;
wire n_4737;
wire n_3647;
wire n_825;
wire n_2819;
wire n_506;
wire n_737;
wire n_5195;
wire n_3609;
wire n_4136;
wire n_1715;
wire n_1952;
wire n_4393;
wire n_3720;
wire n_4535;
wire n_733;
wire n_1922;
wire n_2560;
wire n_4522;
wire n_4794;
wire n_3959;
wire n_792;
wire n_3140;
wire n_5246;
wire n_3724;
wire n_298;
wire n_2104;
wire n_505;
wire n_3011;
wire n_5164;
wire n_4196;
wire n_1425;
wire n_4592;
wire n_4675;
wire n_5340;
wire n_3069;
wire n_5498;
wire n_4370;
wire n_1900;
wire n_1620;
wire n_5183;
wire n_3084;
wire n_1727;
wire n_2735;
wire n_2497;
wire n_3412;
wire n_1995;
wire n_5549;
wire n_2411;
wire n_1046;
wire n_3761;
wire n_4889;
wire n_2014;
wire n_2986;
wire n_5442;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_4828;
wire n_5385;
wire n_4558;
wire n_2172;
wire n_4722;
wire n_1129;
wire n_158;
wire n_4768;
wire n_3626;
wire n_4100;
wire n_961;
wire n_2250;
wire n_276;
wire n_1225;
wire n_169;
wire n_400;
wire n_4092;
wire n_3908;
wire n_2423;
wire n_3671;
wire n_994;
wire n_3344;
wire n_2194;
wire n_848;
wire n_4465;
wire n_3302;
wire n_5537;
wire n_5304;
wire n_1223;
wire n_2680;
wire n_5130;
wire n_1567;
wire n_3122;
wire n_5162;
wire n_4808;
wire n_3842;
wire n_145;
wire n_3265;
wire n_1857;
wire n_4482;
wire n_2041;
wire n_631;
wire n_479;
wire n_1797;
wire n_2957;
wire n_2357;
wire n_1250;
wire n_3309;
wire n_608;
wire n_772;
wire n_3260;
wire n_4926;
wire n_3357;
wire n_1589;
wire n_4116;
wire n_1086;
wire n_2570;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_5473;
wire n_3754;
wire n_4612;
wire n_1469;
wire n_2744;
wire n_4287;
wire n_2397;
wire n_384;
wire n_2208;
wire n_3063;
wire n_5177;
wire n_3617;
wire n_333;
wire n_1298;
wire n_1652;
wire n_4516;
wire n_3794;
wire n_2809;
wire n_2050;
wire n_4505;
wire n_1676;
wire n_258;
wire n_1113;
wire n_1277;
wire n_2591;
wire n_188;
wire n_3384;
wire n_852;
wire n_4602;
wire n_5172;
wire n_4449;
wire n_1864;
wire n_463;
wire n_5070;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_4445;
wire n_699;
wire n_5566;
wire n_5414;
wire n_1627;
wire n_1245;
wire n_4870;
wire n_2438;
wire n_465;
wire n_2832;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_273;
wire n_3181;
wire n_616;
wire n_2278;
wire n_4915;
wire n_5296;
wire n_2135;
wire n_5450;
wire n_3493;
wire n_5313;
wire n_3323;
wire n_2734;
wire n_4914;
wire n_1076;
wire n_2823;
wire n_1408;
wire n_494;
wire n_1761;
wire n_730;
wire n_354;
wire n_5270;
wire n_795;
wire n_4345;
wire n_5188;
wire n_180;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_4318;
wire n_2485;
wire n_2655;
wire n_4185;
wire n_4797;
wire n_2366;
wire n_1526;
wire n_3997;
wire n_1604;
wire n_1275;
wire n_5465;
wire n_4032;
wire n_1764;
wire n_3582;
wire n_712;
wire n_1583;
wire n_2826;
wire n_3539;
wire n_1042;
wire n_285;
wire n_412;
wire n_4343;
wire n_1493;
wire n_4212;
wire n_4124;
wire n_5467;
wire n_5522;
wire n_4492;
wire n_2708;
wire n_5148;
wire n_4994;
wire n_4245;
wire n_4364;
wire n_4928;
wire n_2225;
wire n_1507;
wire n_4378;
wire n_2383;
wire n_1996;
wire n_597;
wire n_3406;
wire n_3604;
wire n_3853;
wire n_4216;
wire n_2019;
wire n_1340;
wire n_1558;
wire n_2166;
wire n_2938;
wire n_4309;
wire n_3594;
wire n_262;
wire n_1704;
wire n_3721;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1234;
wire n_2109;
wire n_364;
wire n_2013;
wire n_1990;
wire n_1032;
wire n_2614;
wire n_2991;
wire n_2242;
wire n_2752;
wire n_2894;
wire n_3473;
wire n_4560;
wire n_5318;
wire n_2839;
wire n_1588;
wire n_5395;
wire n_2237;
wire n_3463;
wire n_3699;
wire n_5067;
wire n_3360;
wire n_2524;
wire n_3873;
wire n_3693;
wire n_2728;
wire n_3857;

CKINVDCx5p33_ASAP7_75t_R g87 ( 
.A(n_60),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_16),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_6),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_40),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_19),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_18),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

CKINVDCx5p33_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_2),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_0),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_63),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_31),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_20),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_44),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_4),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_24),
.Y(n_115)
);

CKINVDCx5p33_ASAP7_75t_R g116 ( 
.A(n_30),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_82),
.Y(n_117)
);

CKINVDCx5p33_ASAP7_75t_R g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_46),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_70),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_27),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_15),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_6),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_79),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_5),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_33),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

BUFx8_ASAP7_75t_SL g128 ( 
.A(n_16),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_7),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_83),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_24),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_54),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_12),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_28),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_32),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_0),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_37),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_78),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_50),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_25),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_25),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_49),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_32),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_19),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_30),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_5),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_48),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_51),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_44),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_3),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_28),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_61),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_37),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_66),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_74),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_64),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_41),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_4),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_66),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_45),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_49),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_29),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_53),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_83),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_63),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_11),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_61),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_39),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_105),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVxp33_ASAP7_75t_SL g184 ( 
.A(n_99),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_105),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_111),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_91),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_123),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_111),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_111),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_136),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_173),
.B(n_169),
.Y(n_199)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_169),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_185),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_123),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

BUFx8_ASAP7_75t_SL g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_195),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_190),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_120),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_195),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_120),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_175),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_169),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_175),
.B(n_169),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_115),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_178),
.Y(n_223)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_180),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_115),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g227 ( 
.A(n_178),
.B(n_120),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_178),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_181),
.B(n_120),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

BUFx8_ASAP7_75t_SL g231 ( 
.A(n_174),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g234 ( 
.A(n_182),
.B(n_115),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_182),
.B(n_94),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_199),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_182),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

BUFx8_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_222),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_208),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_187),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_234),
.B(n_127),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_213),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_127),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_177),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_182),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_213),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_200),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

AND3x2_ASAP7_75t_L g260 ( 
.A(n_204),
.B(n_142),
.C(n_127),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_200),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_226),
.B(n_183),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_213),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_234),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_183),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_221),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_214),
.B(n_183),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_199),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_202),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_202),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_208),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_183),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_216),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_202),
.Y(n_283)
);

AND2x6_ASAP7_75t_L g284 ( 
.A(n_200),
.B(n_188),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_202),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_208),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_201),
.B(n_188),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_223),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

NAND2xp33_ASAP7_75t_SL g290 ( 
.A(n_204),
.B(n_142),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_201),
.B(n_188),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_223),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_201),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_201),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_201),
.B(n_188),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_201),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_205),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_214),
.B(n_192),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g301 ( 
.A(n_225),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_223),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_202),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_219),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_205),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_223),
.Y(n_307)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_229),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_216),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_205),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_193),
.B(n_192),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_219),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_227),
.B(n_196),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_200),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_214),
.B(n_192),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_200),
.B(n_192),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_219),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_205),
.B(n_193),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_219),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_224),
.B(n_177),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_219),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_223),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_222),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_205),
.B(n_193),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_219),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_232),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_223),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_223),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_205),
.B(n_193),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_211),
.B(n_194),
.Y(n_336)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_239),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_239),
.Y(n_339)
);

OAI22xp33_ASAP7_75t_L g340 ( 
.A1(n_252),
.A2(n_196),
.B1(n_191),
.B2(n_150),
.Y(n_340)
);

OR2x6_ASAP7_75t_L g341 ( 
.A(n_308),
.B(n_225),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_239),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_239),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_239),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_246),
.B(n_177),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_270),
.B(n_222),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_251),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_251),
.Y(n_348)
);

AOI21x1_ASAP7_75t_L g349 ( 
.A1(n_237),
.A2(n_226),
.B(n_220),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_251),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_251),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_270),
.B(n_222),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_251),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_255),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_255),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_255),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_255),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_255),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_236),
.B(n_211),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_256),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_270),
.B(n_225),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_256),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_256),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_256),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_236),
.B(n_211),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_256),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_257),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_236),
.B(n_225),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_257),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_308),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_257),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_257),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_257),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_263),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_263),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_263),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_263),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_263),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_248),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_246),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_247),
.B(n_224),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_247),
.B(n_252),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_248),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_248),
.Y(n_386)
);

INVxp33_ASAP7_75t_L g387 ( 
.A(n_244),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_236),
.B(n_240),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_269),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_269),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_332),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_240),
.B(n_259),
.Y(n_394)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_308),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_332),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_247),
.B(n_224),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_294),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_240),
.B(n_211),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_240),
.B(n_211),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_294),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_269),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_269),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_295),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_269),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_295),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_269),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_269),
.Y(n_410)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_313),
.B(n_221),
.C(n_227),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_269),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_300),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_237),
.A2(n_292),
.B(n_287),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_295),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_259),
.B(n_196),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_259),
.B(n_225),
.Y(n_417)
);

CKINVDCx6p67_ASAP7_75t_R g418 ( 
.A(n_247),
.Y(n_418)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_301),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_259),
.B(n_211),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_247),
.A2(n_170),
.B1(n_142),
.B2(n_147),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_264),
.B(n_232),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_300),
.Y(n_423)
);

NAND3xp33_ASAP7_75t_L g424 ( 
.A(n_313),
.B(n_221),
.C(n_227),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_327),
.Y(n_425)
);

OAI22xp33_ASAP7_75t_L g426 ( 
.A1(n_252),
.A2(n_191),
.B1(n_147),
.B2(n_150),
.Y(n_426)
);

AO21x2_ASAP7_75t_L g427 ( 
.A1(n_253),
.A2(n_226),
.B(n_235),
.Y(n_427)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_273),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_247),
.A2(n_224),
.B1(n_216),
.B2(n_184),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_246),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_264),
.B(n_232),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_300),
.Y(n_432)
);

CKINVDCx6p67_ASAP7_75t_R g433 ( 
.A(n_249),
.Y(n_433)
);

AOI21x1_ASAP7_75t_L g434 ( 
.A1(n_237),
.A2(n_226),
.B(n_220),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_238),
.B(n_224),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_264),
.B(n_232),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_300),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_238),
.B(n_224),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_327),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_273),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_308),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_298),
.Y(n_442)
);

AND2x6_ASAP7_75t_L g443 ( 
.A(n_241),
.B(n_214),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_264),
.B(n_232),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_265),
.B(n_232),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_308),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_265),
.B(n_225),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_298),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_298),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_300),
.Y(n_450)
);

OAI21xp33_ASAP7_75t_SL g451 ( 
.A1(n_265),
.A2(n_235),
.B(n_191),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_249),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_299),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_300),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_299),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_300),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_265),
.B(n_225),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_275),
.A2(n_184),
.B1(n_176),
.B2(n_136),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_301),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_273),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_238),
.B(n_224),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_300),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_299),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_275),
.B(n_276),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_275),
.B(n_214),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_306),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_306),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_275),
.B(n_225),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_238),
.B(n_225),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_276),
.A2(n_147),
.B1(n_150),
.B2(n_170),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_306),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_276),
.A2(n_170),
.B1(n_94),
.B2(n_176),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_310),
.Y(n_473)
);

INVx8_ASAP7_75t_L g474 ( 
.A(n_301),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_310),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g476 ( 
.A(n_328),
.B(n_153),
.Y(n_476)
);

INVx6_ASAP7_75t_L g477 ( 
.A(n_308),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_242),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_310),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_243),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_276),
.B(n_214),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_243),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_277),
.B(n_207),
.Y(n_483)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_246),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_277),
.B(n_207),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_243),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_238),
.B(n_200),
.Y(n_487)
);

AO21x2_ASAP7_75t_L g488 ( 
.A1(n_253),
.A2(n_235),
.B(n_220),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_308),
.Y(n_489)
);

OAI22xp33_ASAP7_75t_L g490 ( 
.A1(n_281),
.A2(n_309),
.B1(n_277),
.B2(n_283),
.Y(n_490)
);

INVxp33_ASAP7_75t_L g491 ( 
.A(n_244),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_243),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_243),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_243),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_241),
.B(n_216),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_243),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_243),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_277),
.A2(n_176),
.B1(n_108),
.B2(n_107),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_274),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_274),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_274),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_327),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_274),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_274),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_274),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_238),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_281),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_250),
.B(n_180),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_274),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_238),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_274),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_278),
.B(n_207),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_279),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_279),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_238),
.B(n_200),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_279),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_279),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_279),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_238),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_278),
.B(n_207),
.Y(n_520)
);

AND2x2_ASAP7_75t_SL g521 ( 
.A(n_328),
.B(n_311),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_279),
.Y(n_522)
);

AND3x2_ASAP7_75t_L g523 ( 
.A(n_250),
.B(n_92),
.C(n_90),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_250),
.B(n_179),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_278),
.B(n_157),
.Y(n_525)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_279),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_238),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_278),
.B(n_207),
.Y(n_528)
);

CKINVDCx6p67_ASAP7_75t_R g529 ( 
.A(n_253),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_279),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_286),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_283),
.B(n_285),
.Y(n_532)
);

OAI22xp33_ASAP7_75t_L g533 ( 
.A1(n_281),
.A2(n_157),
.B1(n_166),
.B2(n_167),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_283),
.B(n_216),
.Y(n_534)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_286),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_250),
.B(n_179),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_244),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_283),
.B(n_166),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_421),
.B(n_197),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_309),
.Y(n_541)
);

AND2x2_ASAP7_75t_SL g542 ( 
.A(n_429),
.B(n_328),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_474),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_377),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_452),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_377),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_351),
.B(n_285),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_377),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_377),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_338),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_345),
.B(n_242),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_338),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_390),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_338),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_338),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_421),
.B(n_197),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_425),
.B(n_268),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_339),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_339),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_339),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_339),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_349),
.A2(n_304),
.B(n_285),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_425),
.B(n_268),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_343),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_390),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_343),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_439),
.B(n_502),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_309),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_343),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_474),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_343),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_351),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_340),
.B(n_209),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_534),
.B(n_285),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_452),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_344),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_344),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_351),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_478),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_344),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_344),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_347),
.Y(n_583)
);

OR2x6_ASAP7_75t_L g584 ( 
.A(n_395),
.B(n_244),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_347),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_340),
.B(n_426),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_347),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_347),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_465),
.A2(n_328),
.B(n_305),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_502),
.B(n_268),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_348),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_348),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_348),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_478),
.B(n_268),
.Y(n_594)
);

INVxp67_ASAP7_75t_SL g595 ( 
.A(n_348),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_350),
.Y(n_596)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_345),
.B(n_244),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_346),
.B(n_290),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_346),
.B(n_290),
.Y(n_599)
);

INVxp33_ASAP7_75t_L g600 ( 
.A(n_345),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_350),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_350),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_350),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_354),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_353),
.B(n_304),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_390),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_389),
.B(n_304),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_426),
.B(n_209),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_354),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_354),
.Y(n_610)
);

INVxp33_ASAP7_75t_L g611 ( 
.A(n_508),
.Y(n_611)
);

AND2x6_ASAP7_75t_SL g612 ( 
.A(n_353),
.B(n_90),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_416),
.B(n_304),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_354),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_358),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_358),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_358),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_358),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_359),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_433),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g621 ( 
.A(n_433),
.B(n_209),
.Y(n_621)
);

NAND2x1p5_ASAP7_75t_L g622 ( 
.A(n_351),
.B(n_286),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_359),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_359),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_416),
.B(n_305),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_433),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_508),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_359),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_395),
.B(n_477),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_363),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_363),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_363),
.Y(n_632)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_470),
.B(n_231),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_363),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_364),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_416),
.B(n_305),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_429),
.B(n_241),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_418),
.B(n_241),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_385),
.B(n_305),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_364),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_395),
.B(n_477),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_364),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_364),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_367),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_367),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_367),
.Y(n_646)
);

NAND2x1p5_ASAP7_75t_L g647 ( 
.A(n_351),
.B(n_286),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_367),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_524),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_368),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_368),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_368),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_368),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_370),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_411),
.A2(n_317),
.B(n_312),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_370),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_382),
.B(n_312),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_370),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_370),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_389),
.B(n_394),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_385),
.B(n_312),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_372),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_372),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_SL g664 ( 
.A(n_418),
.B(n_231),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_372),
.Y(n_665)
);

INVxp33_ASAP7_75t_L g666 ( 
.A(n_524),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_372),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_391),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_524),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_373),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_373),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_411),
.A2(n_317),
.B(n_312),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_385),
.B(n_317),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_394),
.B(n_317),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_373),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_351),
.B(n_241),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_385),
.B(n_321),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_373),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_375),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_395),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_536),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_375),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_464),
.B(n_321),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_391),
.B(n_291),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_386),
.B(n_321),
.Y(n_685)
);

XOR2xp5_ASAP7_75t_L g686 ( 
.A(n_470),
.B(n_231),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_375),
.Y(n_687)
);

BUFx6f_ASAP7_75t_L g688 ( 
.A(n_351),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_386),
.B(n_381),
.Y(n_689)
);

INVx4_ASAP7_75t_SL g690 ( 
.A(n_495),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_351),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_375),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_376),
.Y(n_693)
);

XNOR2x2_ASAP7_75t_L g694 ( 
.A(n_384),
.B(n_323),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_376),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_376),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_376),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_378),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_378),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_378),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_378),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_536),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_536),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_458),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_379),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_379),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_379),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_443),
.Y(n_708)
);

CKINVDCx20_ASAP7_75t_R g709 ( 
.A(n_458),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_351),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_386),
.B(n_321),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_379),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_342),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_342),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_342),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_474),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_352),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_386),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_352),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_464),
.B(n_325),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_352),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_391),
.B(n_291),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_424),
.A2(n_331),
.B(n_325),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_355),
.Y(n_724)
);

XNOR2x2_ASAP7_75t_L g725 ( 
.A(n_384),
.B(n_323),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_382),
.B(n_325),
.Y(n_726)
);

INVxp67_ASAP7_75t_SL g727 ( 
.A(n_516),
.Y(n_727)
);

NOR2xp67_ASAP7_75t_L g728 ( 
.A(n_525),
.B(n_323),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_467),
.Y(n_729)
);

XOR2xp5_ASAP7_75t_L g730 ( 
.A(n_533),
.B(n_231),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_467),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_467),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_369),
.B(n_325),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_388),
.Y(n_734)
);

OAI21xp5_ASAP7_75t_L g735 ( 
.A1(n_424),
.A2(n_331),
.B(n_286),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_532),
.B(n_331),
.Y(n_736)
);

INVx4_ASAP7_75t_SL g737 ( 
.A(n_495),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_SL g738 ( 
.A(n_383),
.B(n_241),
.Y(n_738)
);

CKINVDCx20_ASAP7_75t_R g739 ( 
.A(n_382),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_388),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_430),
.B(n_331),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_388),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_474),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_430),
.B(n_260),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_355),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_532),
.B(n_286),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_388),
.Y(n_747)
);

INVxp33_ASAP7_75t_SL g748 ( 
.A(n_440),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_404),
.B(n_291),
.Y(n_749)
);

BUFx6f_ASAP7_75t_SL g750 ( 
.A(n_404),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_430),
.Y(n_751)
);

CKINVDCx16_ASAP7_75t_R g752 ( 
.A(n_476),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_355),
.Y(n_753)
);

AOI21x1_ASAP7_75t_L g754 ( 
.A1(n_349),
.A2(n_315),
.B(n_271),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_392),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_474),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_392),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_392),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_SL g759 ( 
.A(n_383),
.B(n_241),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_392),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_484),
.B(n_260),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_393),
.Y(n_762)
);

XOR2x2_ASAP7_75t_L g763 ( 
.A(n_472),
.B(n_260),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_484),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_393),
.Y(n_765)
);

OAI21xp5_ASAP7_75t_L g766 ( 
.A1(n_465),
.A2(n_286),
.B(n_267),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_525),
.B(n_241),
.Y(n_767)
);

CKINVDCx16_ASAP7_75t_R g768 ( 
.A(n_476),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_381),
.B(n_271),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_356),
.Y(n_770)
);

CKINVDCx20_ASAP7_75t_R g771 ( 
.A(n_484),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_393),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_381),
.B(n_271),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_393),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_538),
.B(n_271),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_396),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_404),
.B(n_291),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_396),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_396),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_396),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_398),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_538),
.B(n_271),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_398),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_575),
.B(n_387),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_586),
.A2(n_418),
.B1(n_397),
.B2(n_387),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_598),
.B(n_599),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_735),
.A2(n_451),
.B(n_417),
.Y(n_787)
);

NOR2x1p5_ASAP7_75t_L g788 ( 
.A(n_626),
.B(n_529),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_586),
.A2(n_397),
.B1(n_537),
.B2(n_491),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_575),
.B(n_541),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_567),
.B(n_551),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_557),
.B(n_440),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_542),
.A2(n_537),
.B1(n_491),
.B2(n_407),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_605),
.B(n_428),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_542),
.A2(n_625),
.B1(n_636),
.B2(n_613),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_570),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_689),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_689),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_716),
.B(n_474),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_660),
.B(n_428),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_629),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_674),
.B(n_460),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_683),
.B(n_460),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_541),
.B(n_507),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_545),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_729),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_563),
.B(n_380),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_637),
.A2(n_451),
.B1(n_356),
.B2(n_361),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_608),
.B(n_380),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_748),
.B(n_533),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_716),
.B(n_474),
.Y(n_811)
);

OR2x6_ASAP7_75t_L g812 ( 
.A(n_629),
.B(n_474),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_720),
.B(n_507),
.Y(n_813)
);

BUFx6f_ASAP7_75t_SL g814 ( 
.A(n_629),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_729),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_731),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_733),
.A2(n_728),
.B1(n_607),
.B2(n_736),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_657),
.B(n_380),
.Y(n_818)
);

OAI221xp5_ASAP7_75t_L g819 ( 
.A1(n_539),
.A2(n_472),
.B1(n_498),
.B2(n_407),
.C(n_410),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_726),
.B(n_380),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_733),
.B(n_356),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_733),
.B(n_357),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_733),
.A2(n_357),
.B1(n_365),
.B2(n_361),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_733),
.B(n_357),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_745),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_745),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_748),
.B(n_498),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_716),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_741),
.B(n_380),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_753),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_733),
.B(n_639),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_611),
.B(n_361),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_775),
.B(n_365),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_SL g834 ( 
.A(n_574),
.B(n_337),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_731),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_775),
.B(n_365),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_732),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_553),
.B(n_380),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_553),
.B(n_565),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_716),
.B(n_743),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_565),
.B(n_402),
.Y(n_841)
);

OR2x6_ASAP7_75t_L g842 ( 
.A(n_629),
.B(n_374),
.Y(n_842)
);

BUFx12f_ASAP7_75t_L g843 ( 
.A(n_626),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_733),
.A2(n_374),
.B1(n_490),
.B2(n_417),
.Y(n_844)
);

INVxp33_ASAP7_75t_L g845 ( 
.A(n_666),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_655),
.A2(n_369),
.B1(n_457),
.B2(n_447),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_732),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_753),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_641),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_770),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_606),
.B(n_402),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_639),
.B(n_374),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_661),
.B(n_481),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_600),
.B(n_481),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_661),
.B(n_490),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_672),
.A2(n_447),
.B1(n_468),
.B2(n_457),
.Y(n_856)
);

BUFx8_ASAP7_75t_SL g857 ( 
.A(n_620),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_606),
.B(n_402),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_668),
.B(n_752),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_764),
.B(n_405),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_590),
.B(n_405),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_668),
.B(n_402),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_547),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_770),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_590),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_769),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_769),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_782),
.B(n_468),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_718),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_568),
.B(n_782),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_718),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_568),
.B(n_405),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_560),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_560),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_746),
.A2(n_526),
.B(n_516),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_673),
.B(n_407),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_673),
.B(n_409),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_544),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_768),
.B(n_402),
.Y(n_879)
);

OAI22x1_ASAP7_75t_L g880 ( 
.A1(n_539),
.A2(n_556),
.B1(n_686),
.B2(n_633),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_677),
.B(n_409),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_540),
.B(n_669),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_677),
.B(n_409),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_685),
.B(n_410),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_739),
.B(n_751),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_544),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_771),
.B(n_410),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_548),
.Y(n_889)
);

NAND2x1_ASAP7_75t_L g890 ( 
.A(n_543),
.B(n_337),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_723),
.A2(n_362),
.B(n_413),
.C(n_412),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_556),
.B(n_412),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_594),
.Y(n_893)
);

OAI22xp5_ASAP7_75t_L g894 ( 
.A1(n_685),
.A2(n_529),
.B1(n_362),
.B2(n_366),
.Y(n_894)
);

INVxp67_ASAP7_75t_L g895 ( 
.A(n_594),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_548),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_580),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_597),
.A2(n_529),
.B1(n_412),
.B2(n_423),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_711),
.B(n_360),
.Y(n_899)
);

NOR2xp67_ASAP7_75t_L g900 ( 
.A(n_680),
.B(n_413),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_R g901 ( 
.A(n_580),
.B(n_349),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_577),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_597),
.B(n_413),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_684),
.B(n_402),
.Y(n_904)
);

INVxp67_ASAP7_75t_L g905 ( 
.A(n_744),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_767),
.A2(n_438),
.B(n_461),
.C(n_435),
.Y(n_906)
);

INVxp33_ASAP7_75t_L g907 ( 
.A(n_633),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_684),
.B(n_441),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_711),
.B(n_360),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_684),
.B(n_441),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_641),
.B(n_423),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_722),
.B(n_441),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_584),
.A2(n_529),
.B1(n_423),
.B2(n_437),
.Y(n_913)
);

AOI22xp5_ASAP7_75t_L g914 ( 
.A1(n_584),
.A2(n_704),
.B1(n_709),
.B2(n_738),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_641),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_595),
.B(n_366),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_722),
.B(n_441),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_576),
.B(n_489),
.C(n_441),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_763),
.A2(n_450),
.B1(n_454),
.B2(n_437),
.C(n_432),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_584),
.A2(n_432),
.B1(n_450),
.B2(n_437),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_584),
.A2(n_759),
.B1(n_763),
.B2(n_547),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_577),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_549),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_722),
.B(n_441),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_596),
.B(n_399),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_773),
.B(n_399),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_749),
.B(n_489),
.Y(n_927)
);

BUFx5_ASAP7_75t_L g928 ( 
.A(n_547),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_749),
.B(n_489),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_581),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_581),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_641),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_773),
.B(n_400),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_609),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_609),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_547),
.A2(n_432),
.B1(n_454),
.B2(n_450),
.Y(n_936)
);

INVx2_ASAP7_75t_SL g937 ( 
.A(n_749),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_547),
.A2(n_454),
.B1(n_462),
.B2(n_456),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_589),
.B(n_400),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_549),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_761),
.B(n_456),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_638),
.A2(n_420),
.B1(n_431),
.B2(n_422),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_643),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_777),
.B(n_489),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_643),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_727),
.B(n_456),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_627),
.B(n_462),
.Y(n_947)
);

AND2x4_ASAP7_75t_SL g948 ( 
.A(n_743),
.B(n_506),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_686),
.B(n_462),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_547),
.A2(n_488),
.B1(n_315),
.B2(n_427),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_658),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_734),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_658),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_550),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_546),
.B(n_506),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_777),
.B(n_489),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_777),
.B(n_521),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_649),
.B(n_523),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_550),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_734),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_766),
.B(n_506),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_740),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_602),
.B(n_506),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_554),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_740),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_681),
.B(n_523),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_554),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_573),
.B(n_489),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_602),
.B(n_506),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_742),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_713),
.B(n_420),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_555),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_573),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_610),
.B(n_506),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_610),
.B(n_510),
.Y(n_975)
);

INVx8_ASAP7_75t_L g976 ( 
.A(n_547),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_680),
.A2(n_477),
.B1(n_395),
.B2(n_487),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_645),
.B(n_646),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_680),
.B(n_521),
.Y(n_979)
);

INVx4_ASAP7_75t_L g980 ( 
.A(n_743),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_750),
.A2(n_488),
.B1(n_315),
.B2(n_427),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_573),
.B(n_371),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_714),
.A2(n_438),
.B(n_461),
.C(n_435),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_645),
.B(n_510),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_555),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_715),
.B(n_483),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_558),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_573),
.Y(n_988)
);

NOR2xp67_ASAP7_75t_L g989 ( 
.A(n_558),
.B(n_510),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_750),
.A2(n_477),
.B1(n_395),
.B2(n_487),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_646),
.B(n_510),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_717),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_573),
.B(n_371),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_579),
.B(n_371),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_719),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_721),
.B(n_521),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_724),
.B(n_510),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_742),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_559),
.B(n_510),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_559),
.B(n_519),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_561),
.B(n_422),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_579),
.B(n_446),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_702),
.B(n_395),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_561),
.B(n_431),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_564),
.B(n_436),
.Y(n_1005)
);

NOR3xp33_ASAP7_75t_L g1006 ( 
.A(n_676),
.B(n_515),
.C(n_469),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_747),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_622),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_579),
.B(n_446),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_564),
.B(n_566),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_730),
.B(n_515),
.C(n_469),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_638),
.A2(n_444),
.B1(n_445),
.B2(n_436),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_621),
.Y(n_1013)
);

NOR2x1p5_ASAP7_75t_L g1014 ( 
.A(n_743),
.B(n_519),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_747),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_566),
.B(n_444),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_755),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_703),
.B(n_477),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_569),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_569),
.B(n_445),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_572),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_572),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_750),
.A2(n_477),
.B1(n_446),
.B2(n_291),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_543),
.B(n_337),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_755),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_578),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_781),
.A2(n_783),
.B(n_267),
.C(n_758),
.Y(n_1027)
);

INVxp67_ASAP7_75t_SL g1028 ( 
.A(n_579),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_579),
.B(n_521),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_578),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_582),
.B(n_488),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_582),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_730),
.B(n_477),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_583),
.B(n_483),
.Y(n_1034)
);

INVx2_ASAP7_75t_SL g1035 ( 
.A(n_781),
.Y(n_1035)
);

OR2x6_ASAP7_75t_L g1036 ( 
.A(n_743),
.B(n_341),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_694),
.A2(n_527),
.B1(n_519),
.B2(n_238),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_583),
.B(n_519),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_585),
.B(n_519),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_585),
.B(n_519),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_587),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_664),
.A2(n_488),
.B1(n_315),
.B2(n_427),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_587),
.A2(n_526),
.B1(n_530),
.B2(n_516),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_688),
.B(n_337),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_588),
.B(n_527),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_783),
.A2(n_488),
.B1(n_315),
.B2(n_427),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_688),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_688),
.B(n_691),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_588),
.B(n_527),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_688),
.B(n_337),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_688),
.B(n_337),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_591),
.B(n_527),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_591),
.B(n_527),
.Y(n_1053)
);

OR2x2_ASAP7_75t_L g1054 ( 
.A(n_592),
.B(n_485),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_757),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_592),
.B(n_485),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_593),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_757),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_543),
.B(n_419),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_622),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_593),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_758),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_601),
.B(n_527),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_760),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_622),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_571),
.B(n_419),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_760),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_762),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_691),
.B(n_419),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_601),
.B(n_434),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_603),
.B(n_512),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_603),
.B(n_512),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_604),
.B(n_434),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_604),
.B(n_434),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_762),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_614),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_614),
.B(n_427),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_765),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_615),
.B(n_520),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_765),
.Y(n_1080)
);

NOR2xp67_ASAP7_75t_L g1081 ( 
.A(n_615),
.B(n_616),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_616),
.B(n_617),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_647),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_612),
.B(n_520),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_562),
.B(n_528),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_691),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_617),
.B(n_528),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_618),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_691),
.B(n_419),
.Y(n_1089)
);

INVx8_ASAP7_75t_L g1090 ( 
.A(n_691),
.Y(n_1090)
);

NAND3xp33_ASAP7_75t_L g1091 ( 
.A(n_772),
.B(n_262),
.C(n_254),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_618),
.B(n_482),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_772),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_774),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_552),
.A2(n_262),
.B1(n_280),
.B2(n_254),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_562),
.B(n_414),
.Y(n_1096)
);

AO221x1_ASAP7_75t_L g1097 ( 
.A1(n_694),
.A2(n_101),
.B1(n_103),
.B2(n_172),
.C(n_92),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_774),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_776),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_644),
.B(n_414),
.Y(n_1100)
);

NOR2xp67_ASAP7_75t_L g1101 ( 
.A(n_619),
.B(n_267),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_648),
.B(n_414),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_710),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_710),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_870),
.B(n_619),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_973),
.Y(n_1106)
);

INVx11_ASAP7_75t_L g1107 ( 
.A(n_843),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_795),
.A2(n_710),
.B1(n_530),
.B2(n_535),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_905),
.B(n_153),
.Y(n_1109)
);

INVxp67_ASAP7_75t_L g1110 ( 
.A(n_882),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_939),
.A2(n_925),
.B(n_916),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_796),
.B(n_710),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_939),
.A2(n_571),
.B(n_459),
.Y(n_1113)
);

AO21x1_ASAP7_75t_L g1114 ( 
.A1(n_846),
.A2(n_725),
.B(n_647),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_796),
.B(n_710),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_916),
.A2(n_571),
.B(n_459),
.Y(n_1116)
);

INVx3_ASAP7_75t_L g1117 ( 
.A(n_812),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_L g1118 ( 
.A(n_1103),
.B(n_756),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_870),
.B(n_623),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_806),
.Y(n_1120)
);

NOR2xp33_ASAP7_75t_L g1121 ( 
.A(n_786),
.B(n_159),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_890),
.A2(n_1059),
.B(n_875),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_925),
.A2(n_459),
.B(n_419),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_806),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_790),
.B(n_623),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_815),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_799),
.A2(n_459),
.B(n_419),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_954),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_795),
.A2(n_856),
.B1(n_846),
.B2(n_919),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_856),
.A2(n_103),
.B(n_104),
.C(n_101),
.Y(n_1130)
);

OR2x6_ASAP7_75t_L g1131 ( 
.A(n_812),
.B(n_756),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_811),
.A2(n_459),
.B(n_526),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_814),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_791),
.A2(n_106),
.B(n_129),
.C(n_104),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_790),
.B(n_624),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_865),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_901),
.B(n_756),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1024),
.A2(n_459),
.B(n_530),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_SL g1139 ( 
.A(n_814),
.B(n_756),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1024),
.A2(n_535),
.B(n_647),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_854),
.B(n_624),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_794),
.B(n_628),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1066),
.A2(n_535),
.B(n_756),
.Y(n_1143)
);

CKINVDCx16_ASAP7_75t_R g1144 ( 
.A(n_843),
.Y(n_1144)
);

INVx11_ASAP7_75t_L g1145 ( 
.A(n_843),
.Y(n_1145)
);

NOR2xp67_ASAP7_75t_L g1146 ( 
.A(n_801),
.B(n_628),
.Y(n_1146)
);

AOI21x1_ASAP7_75t_L g1147 ( 
.A1(n_894),
.A2(n_754),
.B(n_776),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_983),
.A2(n_129),
.B(n_131),
.C(n_106),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_784),
.B(n_630),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1066),
.A2(n_341),
.B(n_482),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_906),
.A2(n_341),
.B(n_482),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1084),
.A2(n_131),
.B(n_140),
.C(n_134),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_844),
.A2(n_631),
.B1(n_632),
.B2(n_630),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_894),
.A2(n_754),
.B(n_778),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_954),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_802),
.A2(n_341),
.B(n_482),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_954),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_891),
.A2(n_779),
.B(n_780),
.C(n_778),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_959),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_787),
.A2(n_651),
.B(n_650),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_802),
.A2(n_341),
.B(n_492),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1011),
.A2(n_160),
.B1(n_167),
.B2(n_159),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_L g1163 ( 
.A1(n_914),
.A2(n_725),
.B1(n_108),
.B2(n_107),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_784),
.B(n_631),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_810),
.A2(n_134),
.B(n_148),
.C(n_140),
.Y(n_1165)
);

AOI21x1_ASAP7_75t_L g1166 ( 
.A1(n_942),
.A2(n_780),
.B(n_779),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_804),
.B(n_632),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_815),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_845),
.B(n_160),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_804),
.B(n_634),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_816),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_827),
.B(n_238),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_941),
.B(n_634),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_887),
.B(n_245),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_787),
.A2(n_640),
.B(n_642),
.C(n_635),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_942),
.A2(n_401),
.B(n_398),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_803),
.A2(n_341),
.B(n_492),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_812),
.Y(n_1178)
);

OAI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_817),
.A2(n_653),
.B(n_652),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_803),
.A2(n_341),
.B(n_492),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_L g1181 ( 
.A(n_947),
.B(n_245),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_792),
.A2(n_148),
.B(n_156),
.C(n_151),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_800),
.B(n_635),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_844),
.A2(n_642),
.B1(n_679),
.B2(n_640),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_817),
.A2(n_401),
.B(n_403),
.C(n_398),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_785),
.A2(n_403),
.B(n_406),
.C(n_401),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_973),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_865),
.B(n_679),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_959),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_800),
.A2(n_687),
.B1(n_692),
.B2(n_682),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_959),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_892),
.B(n_682),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_937),
.B(n_687),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_964),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_893),
.B(n_245),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_937),
.B(n_692),
.Y(n_1196)
);

AND2x2_ASAP7_75t_SL g1197 ( 
.A(n_834),
.B(n_693),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_861),
.B(n_813),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_819),
.A2(n_495),
.B1(n_443),
.B2(n_88),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_823),
.A2(n_789),
.B1(n_921),
.B2(n_909),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_895),
.B(n_245),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_957),
.B(n_693),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_899),
.A2(n_341),
.B(n_492),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_832),
.B(n_695),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1006),
.A2(n_403),
.B(n_406),
.C(n_401),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_899),
.A2(n_496),
.B(n_493),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_868),
.A2(n_696),
.B(n_697),
.C(n_695),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_801),
.B(n_696),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_903),
.B(n_697),
.Y(n_1209)
);

INVx1_ASAP7_75t_SL g1210 ( 
.A(n_957),
.Y(n_1210)
);

AO21x1_ASAP7_75t_L g1211 ( 
.A1(n_1012),
.A2(n_698),
.B(n_656),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_949),
.A2(n_254),
.B1(n_280),
.B2(n_262),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_812),
.Y(n_1213)
);

NOR2x1p5_ASAP7_75t_SL g1214 ( 
.A(n_863),
.B(n_708),
.Y(n_1214)
);

OAI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_880),
.A2(n_88),
.B1(n_89),
.B2(n_87),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_909),
.A2(n_496),
.B(n_493),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_950),
.A2(n_1012),
.B(n_1085),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_964),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_921),
.A2(n_403),
.B(n_408),
.C(n_406),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_950),
.A2(n_659),
.B(n_654),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_816),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_872),
.B(n_698),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_964),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_866),
.B(n_662),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_911),
.B(n_663),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_L g1226 ( 
.A1(n_1044),
.A2(n_667),
.B(n_670),
.C(n_665),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_866),
.B(n_671),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_840),
.A2(n_496),
.B(n_493),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_823),
.A2(n_486),
.B1(n_494),
.B2(n_480),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_918),
.A2(n_280),
.B1(n_216),
.B2(n_675),
.Y(n_1230)
);

O2A1O1Ixp5_ASAP7_75t_L g1231 ( 
.A1(n_1050),
.A2(n_699),
.B(n_700),
.C(n_678),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_808),
.A2(n_705),
.B(n_701),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_859),
.B(n_245),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_961),
.A2(n_496),
.B(n_493),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_853),
.A2(n_500),
.B(n_497),
.Y(n_1235)
);

INVx4_ASAP7_75t_SL g1236 ( 
.A(n_814),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_967),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_853),
.A2(n_500),
.B(n_497),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1036),
.A2(n_500),
.B(n_497),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_L g1240 ( 
.A(n_958),
.B(n_156),
.C(n_151),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1036),
.A2(n_500),
.B(n_497),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1036),
.A2(n_505),
.B(n_504),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_835),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_926),
.B(n_706),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_835),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_926),
.B(n_707),
.Y(n_1246)
);

AOI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1073),
.A2(n_408),
.B(n_406),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_808),
.A2(n_712),
.B(n_415),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1036),
.A2(n_505),
.B(n_504),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_837),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_855),
.A2(n_933),
.B1(n_971),
.B2(n_938),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_814),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_933),
.B(n_504),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_837),
.Y(n_1254)
);

INVx2_ASAP7_75t_SL g1255 ( 
.A(n_1014),
.Y(n_1255)
);

NOR2xp67_ASAP7_75t_L g1256 ( 
.A(n_801),
.B(n_408),
.Y(n_1256)
);

NOR3xp33_ASAP7_75t_L g1257 ( 
.A(n_966),
.B(n_172),
.C(n_235),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_967),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_797),
.B(n_504),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_847),
.Y(n_1260)
);

OAI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1046),
.A2(n_415),
.B(n_408),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1036),
.A2(n_509),
.B(n_505),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1090),
.Y(n_1263)
);

AOI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1073),
.A2(n_442),
.B(n_415),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1033),
.A2(n_216),
.B1(n_221),
.B2(n_95),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_855),
.A2(n_480),
.B1(n_531),
.B2(n_494),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_812),
.A2(n_509),
.B(n_505),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_797),
.B(n_509),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_976),
.A2(n_517),
.B(n_509),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_911),
.B(n_517),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_809),
.A2(n_235),
.B(n_221),
.C(n_287),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1003),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_801),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_976),
.A2(n_518),
.B(n_517),
.Y(n_1274)
);

O2A1O1Ixp5_ASAP7_75t_L g1275 ( 
.A1(n_1051),
.A2(n_479),
.B(n_475),
.C(n_473),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1046),
.A2(n_981),
.B(n_831),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_976),
.A2(n_518),
.B(n_517),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_981),
.A2(n_442),
.B(n_415),
.Y(n_1278)
);

OR2x2_ASAP7_75t_SL g1279 ( 
.A(n_880),
.B(n_442),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_798),
.B(n_518),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_914),
.A2(n_152),
.B1(n_96),
.B2(n_93),
.Y(n_1281)
);

A2O1A1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_913),
.A2(n_442),
.B(n_448),
.C(n_449),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_798),
.B(n_518),
.Y(n_1283)
);

INVx2_ASAP7_75t_SL g1284 ( 
.A(n_1014),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_973),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_976),
.A2(n_522),
.B(n_486),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_996),
.B(n_311),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_973),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_867),
.B(n_286),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_867),
.B(n_448),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1027),
.A2(n_499),
.B(n_480),
.C(n_486),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_967),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_SL g1293 ( 
.A(n_911),
.B(n_860),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_SL g1294 ( 
.A(n_834),
.B(n_495),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_996),
.B(n_876),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_976),
.A2(n_522),
.B(n_499),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_793),
.A2(n_146),
.B1(n_137),
.B2(n_141),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_911),
.B(n_522),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_877),
.B(n_448),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_890),
.A2(n_522),
.B(n_499),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_885),
.B(n_245),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_881),
.B(n_448),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_L g1303 ( 
.A(n_788),
.B(n_708),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_883),
.B(n_449),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_847),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_849),
.B(n_915),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_952),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_884),
.B(n_449),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1059),
.A2(n_501),
.B(n_494),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_831),
.A2(n_453),
.B(n_449),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_833),
.B(n_453),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1043),
.A2(n_503),
.B(n_501),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_979),
.B(n_311),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1043),
.A2(n_503),
.B(n_501),
.Y(n_1314)
);

NOR2x1_ASAP7_75t_L g1315 ( 
.A(n_828),
.B(n_453),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_879),
.B(n_453),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_913),
.A2(n_463),
.B(n_455),
.C(n_466),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_857),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1018),
.B(n_503),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_973),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_972),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1029),
.A2(n_513),
.B(n_511),
.Y(n_1322)
);

OAI321xp33_ASAP7_75t_L g1323 ( 
.A1(n_1042),
.A2(n_119),
.A3(n_220),
.B1(n_514),
.B2(n_513),
.C(n_511),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_852),
.A2(n_513),
.B(n_511),
.Y(n_1324)
);

BUFx4f_ASAP7_75t_L g1325 ( 
.A(n_842),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_852),
.A2(n_531),
.B(n_514),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_821),
.A2(n_463),
.B(n_455),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_836),
.B(n_986),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_972),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_972),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_821),
.A2(n_463),
.B(n_455),
.Y(n_1331)
);

INVx2_ASAP7_75t_SL g1332 ( 
.A(n_1090),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_948),
.A2(n_1004),
.B(n_1001),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_932),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_822),
.A2(n_463),
.B(n_455),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_948),
.A2(n_1004),
.B(n_1001),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_932),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_L g1338 ( 
.A(n_788),
.B(n_708),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_932),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_952),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_985),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_960),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_979),
.B(n_849),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_849),
.A2(n_267),
.B1(n_495),
.B2(n_443),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_985),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_986),
.B(n_466),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_SL g1347 ( 
.A(n_915),
.B(n_495),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_948),
.A2(n_1016),
.B(n_1005),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_915),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_897),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_805),
.B(n_514),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_985),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_822),
.A2(n_471),
.B(n_466),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_971),
.B(n_920),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_960),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1005),
.A2(n_531),
.B(n_708),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1016),
.A2(n_708),
.B(n_495),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_987),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_842),
.B(n_311),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_824),
.A2(n_471),
.B(n_466),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_824),
.A2(n_1042),
.B(n_1091),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_932),
.B(n_690),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_973),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1094),
.B(n_807),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_962),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1094),
.B(n_471),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_839),
.B(n_471),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1091),
.A2(n_1102),
.B(n_1100),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_962),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_965),
.Y(n_1370)
);

AOI21xp5_ASAP7_75t_L g1371 ( 
.A1(n_1020),
.A2(n_708),
.B(n_495),
.Y(n_1371)
);

AOI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1020),
.A2(n_708),
.B(n_495),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_946),
.B(n_473),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1054),
.B(n_473),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1096),
.A2(n_475),
.B(n_473),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1054),
.B(n_475),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_965),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1072),
.B(n_475),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1072),
.B(n_1031),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1090),
.A2(n_708),
.B(n_495),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_898),
.A2(n_89),
.B(n_87),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1031),
.B(n_479),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_L g1383 ( 
.A1(n_1090),
.A2(n_495),
.B(n_443),
.Y(n_1383)
);

INVx2_ASAP7_75t_SL g1384 ( 
.A(n_1090),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_818),
.A2(n_443),
.B(n_479),
.Y(n_1385)
);

A2O1A1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_898),
.A2(n_479),
.B(n_267),
.C(n_227),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_842),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_820),
.B(n_245),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_829),
.A2(n_443),
.B(n_690),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1077),
.B(n_850),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1077),
.B(n_850),
.Y(n_1391)
);

AO21x1_ASAP7_75t_L g1392 ( 
.A1(n_1097),
.A2(n_292),
.B(n_287),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_SL g1393 ( 
.A(n_990),
.B(n_690),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_970),
.Y(n_1394)
);

AOI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1013),
.A2(n_145),
.B1(n_161),
.B2(n_143),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1069),
.A2(n_443),
.B(n_690),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_987),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_977),
.B(n_737),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_907),
.B(n_245),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1089),
.A2(n_443),
.B(n_737),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_936),
.A2(n_227),
.B(n_220),
.C(n_234),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_904),
.B(n_245),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_SL g1403 ( 
.A(n_1023),
.B(n_1047),
.Y(n_1403)
);

O2A1O1Ixp5_ASAP7_75t_L g1404 ( 
.A1(n_982),
.A2(n_336),
.B(n_320),
.C(n_292),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_988),
.Y(n_1405)
);

INVx4_ASAP7_75t_L g1406 ( 
.A(n_842),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_988),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_842),
.A2(n_1056),
.B(n_1034),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1034),
.A2(n_443),
.B(n_737),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1056),
.A2(n_443),
.B(n_737),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1037),
.A2(n_443),
.B(n_320),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_908),
.B(n_245),
.Y(n_1412)
);

AND2x6_ASAP7_75t_L g1413 ( 
.A(n_1047),
.B(n_245),
.Y(n_1413)
);

OAI21xp33_ASAP7_75t_SL g1414 ( 
.A1(n_936),
.A2(n_320),
.B(n_297),
.Y(n_1414)
);

AOI21xp33_ASAP7_75t_L g1415 ( 
.A1(n_938),
.A2(n_98),
.B(n_97),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1079),
.A2(n_330),
.B(n_297),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_828),
.B(n_245),
.Y(n_1417)
);

BUFx4f_ASAP7_75t_L g1418 ( 
.A(n_1047),
.Y(n_1418)
);

AOI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1081),
.A2(n_330),
.B(n_297),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_910),
.B(n_912),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_917),
.B(n_258),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_924),
.B(n_258),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_927),
.B(n_258),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1008),
.A2(n_336),
.B(n_335),
.C(n_330),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1095),
.A2(n_336),
.B(n_335),
.Y(n_1425)
);

BUFx12f_ASAP7_75t_L g1426 ( 
.A(n_1047),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1079),
.A2(n_335),
.B(n_311),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_970),
.Y(n_1428)
);

O2A1O1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_838),
.A2(n_220),
.B(n_234),
.C(n_329),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1087),
.A2(n_311),
.B(n_293),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1087),
.A2(n_311),
.B(n_293),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1071),
.A2(n_311),
.B(n_293),
.Y(n_1432)
);

NOR2xp33_ASAP7_75t_L g1433 ( 
.A(n_929),
.B(n_258),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_998),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1028),
.A2(n_334),
.B(n_293),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_828),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_SL g1437 ( 
.A(n_828),
.B(n_119),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_998),
.Y(n_1438)
);

BUFx6f_ASAP7_75t_L g1439 ( 
.A(n_1047),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_944),
.B(n_258),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_841),
.B(n_149),
.C(n_144),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1048),
.A2(n_334),
.B(n_293),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_956),
.B(n_258),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1092),
.A2(n_296),
.B(n_288),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_963),
.A2(n_296),
.B(n_288),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_SL g1446 ( 
.A(n_888),
.B(n_119),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_825),
.B(n_258),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_969),
.A2(n_296),
.B(n_288),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_974),
.A2(n_296),
.B(n_288),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_975),
.A2(n_296),
.B(n_288),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1047),
.B(n_258),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_984),
.A2(n_303),
.B(n_302),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_991),
.A2(n_303),
.B(n_302),
.Y(n_1453)
);

AOI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_993),
.A2(n_303),
.B(n_302),
.Y(n_1454)
);

OAI321xp33_ASAP7_75t_L g1455 ( 
.A1(n_1095),
.A2(n_119),
.A3(n_171),
.B1(n_168),
.B2(n_165),
.C(n_164),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_825),
.B(n_258),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_994),
.A2(n_303),
.B(n_302),
.Y(n_1457)
);

CKINVDCx10_ASAP7_75t_R g1458 ( 
.A(n_1097),
.Y(n_1458)
);

AOI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1081),
.A2(n_227),
.B(n_194),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_988),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1086),
.B(n_258),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_825),
.B(n_258),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_826),
.B(n_258),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_826),
.B(n_830),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1010),
.A2(n_194),
.B(n_234),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_826),
.B(n_261),
.Y(n_1466)
);

AOI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1010),
.A2(n_194),
.B(n_234),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_830),
.B(n_229),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1007),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_830),
.B(n_261),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_987),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_848),
.B(n_261),
.Y(n_1472)
);

O2A1O1Ixp33_ASAP7_75t_SL g1473 ( 
.A1(n_1002),
.A2(n_334),
.B(n_333),
.C(n_329),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_SL g1474 ( 
.A(n_1086),
.B(n_261),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_851),
.B(n_261),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_848),
.B(n_864),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_888),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1019),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1007),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1086),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1009),
.A2(n_334),
.B(n_333),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1015),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_848),
.B(n_261),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_864),
.B(n_1070),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_858),
.A2(n_234),
.B(n_333),
.C(n_329),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_999),
.A2(n_334),
.B(n_333),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_864),
.B(n_261),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1070),
.B(n_261),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1019),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_888),
.B(n_261),
.Y(n_1490)
);

AOI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1000),
.A2(n_333),
.B(n_329),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1038),
.A2(n_329),
.B(n_326),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1015),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1017),
.Y(n_1494)
);

AOI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1040),
.A2(n_326),
.B(n_324),
.Y(n_1495)
);

BUFx4f_ASAP7_75t_L g1496 ( 
.A(n_1086),
.Y(n_1496)
);

O2A1O1Ixp5_ASAP7_75t_L g1497 ( 
.A1(n_1008),
.A2(n_234),
.B(n_229),
.C(n_324),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1074),
.B(n_261),
.Y(n_1498)
);

NOR2x1_ASAP7_75t_L g1499 ( 
.A(n_888),
.B(n_302),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_862),
.B(n_261),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_992),
.A2(n_100),
.B1(n_97),
.B2(n_98),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1019),
.Y(n_1502)
);

AOI21xp33_ASAP7_75t_L g1503 ( 
.A1(n_1017),
.A2(n_102),
.B(n_171),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1045),
.A2(n_326),
.B(n_324),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1074),
.B(n_261),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_980),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1049),
.A2(n_326),
.B(n_324),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1025),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1021),
.B(n_266),
.Y(n_1509)
);

INVxp67_ASAP7_75t_L g1510 ( 
.A(n_992),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1025),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_995),
.B(n_878),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1021),
.B(n_266),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_995),
.A2(n_100),
.B1(n_102),
.B2(n_109),
.Y(n_1514)
);

O2A1O1Ixp33_ASAP7_75t_L g1515 ( 
.A1(n_968),
.A2(n_234),
.B(n_324),
.C(n_322),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1212),
.A2(n_1062),
.B1(n_1055),
.B2(n_1099),
.Y(n_1516)
);

AO21x1_ASAP7_75t_L g1517 ( 
.A1(n_1129),
.A2(n_1062),
.B(n_1055),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1128),
.Y(n_1518)
);

AOI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1111),
.A2(n_1113),
.B(n_1150),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1121),
.B(n_878),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1128),
.Y(n_1521)
);

BUFx6f_ASAP7_75t_L g1522 ( 
.A(n_1426),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1110),
.B(n_886),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_SL g1524 ( 
.A(n_1162),
.B(n_1086),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1198),
.B(n_886),
.Y(n_1525)
);

NOR2xp67_ASAP7_75t_L g1526 ( 
.A(n_1133),
.B(n_980),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_SL g1527 ( 
.A(n_1162),
.B(n_1086),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1210),
.B(n_1295),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_SL g1529 ( 
.A(n_1272),
.B(n_1104),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1210),
.B(n_889),
.Y(n_1530)
);

AOI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1176),
.A2(n_1082),
.B(n_1067),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1172),
.B(n_1104),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1138),
.A2(n_1104),
.B(n_980),
.Y(n_1533)
);

AND2x6_ASAP7_75t_L g1534 ( 
.A(n_1117),
.B(n_1104),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1212),
.A2(n_1064),
.B1(n_1068),
.B2(n_1099),
.Y(n_1535)
);

AOI21x1_ASAP7_75t_L g1536 ( 
.A1(n_1176),
.A2(n_1067),
.B(n_1064),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1301),
.B(n_889),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1109),
.B(n_896),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1140),
.A2(n_1104),
.B(n_980),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_L g1540 ( 
.A1(n_1116),
.A2(n_1104),
.B(n_1060),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1129),
.A2(n_119),
.B1(n_900),
.B2(n_923),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_SL g1542 ( 
.A1(n_1219),
.A2(n_1173),
.B(n_1186),
.C(n_1137),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1328),
.B(n_896),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1132),
.A2(n_1127),
.B(n_1123),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1120),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_L g1546 ( 
.A1(n_1165),
.A2(n_923),
.B(n_940),
.C(n_997),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1202),
.B(n_940),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1169),
.B(n_1399),
.Y(n_1548)
);

OA21x2_ASAP7_75t_L g1549 ( 
.A1(n_1217),
.A2(n_1075),
.B(n_1068),
.Y(n_1549)
);

BUFx12f_ASAP7_75t_L g1550 ( 
.A(n_1405),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1202),
.B(n_869),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1354),
.B(n_1379),
.Y(n_1552)
);

AOI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1166),
.A2(n_1151),
.B(n_1147),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1143),
.A2(n_1060),
.B(n_1008),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1120),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1156),
.A2(n_1060),
.B(n_1008),
.Y(n_1556)
);

NOR2xp33_ASAP7_75t_L g1557 ( 
.A(n_1195),
.B(n_266),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1201),
.B(n_869),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1161),
.A2(n_1180),
.B(n_1177),
.Y(n_1559)
);

AOI22x1_ASAP7_75t_L g1560 ( 
.A1(n_1163),
.A2(n_1030),
.B1(n_1022),
.B2(n_1026),
.Y(n_1560)
);

BUFx12f_ASAP7_75t_L g1561 ( 
.A(n_1407),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1293),
.B(n_871),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1350),
.B(n_1281),
.Y(n_1563)
);

AOI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1166),
.A2(n_1078),
.B(n_1075),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1197),
.A2(n_1098),
.B1(n_1078),
.B2(n_1080),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1281),
.B(n_266),
.Y(n_1566)
);

HB1xp67_ASAP7_75t_L g1567 ( 
.A(n_1136),
.Y(n_1567)
);

AO22x1_ASAP7_75t_L g1568 ( 
.A1(n_1240),
.A2(n_1098),
.B1(n_1080),
.B2(n_1035),
.Y(n_1568)
);

AND2x2_ASAP7_75t_SL g1569 ( 
.A(n_1197),
.B(n_1060),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1343),
.B(n_871),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1343),
.B(n_871),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1131),
.B(n_1406),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1152),
.A2(n_1065),
.B(n_1083),
.C(n_955),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1294),
.A2(n_1083),
.B(n_1065),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1125),
.B(n_1021),
.Y(n_1575)
);

AOI21xp5_ASAP7_75t_L g1576 ( 
.A1(n_1294),
.A2(n_1083),
.B(n_1065),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1192),
.B(n_1022),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1276),
.B(n_1022),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_SL g1579 ( 
.A1(n_1163),
.A2(n_133),
.B1(n_110),
.B2(n_112),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1460),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1181),
.B(n_863),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_SL g1582 ( 
.A(n_1263),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_SL g1583 ( 
.A1(n_1319),
.A2(n_1093),
.B(n_1058),
.C(n_1035),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1215),
.B(n_1503),
.Y(n_1584)
);

AOI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1333),
.A2(n_1348),
.B(n_1336),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1426),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1125),
.B(n_1026),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_SL g1588 ( 
.A(n_1174),
.B(n_863),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1408),
.A2(n_1083),
.B(n_1065),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1141),
.B(n_1251),
.Y(n_1590)
);

OAI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1197),
.A2(n_1058),
.B1(n_1093),
.B2(n_1088),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1251),
.B(n_1144),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1318),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1200),
.A2(n_1199),
.B1(n_1209),
.B2(n_1217),
.Y(n_1594)
);

AOI21xp5_ASAP7_75t_L g1595 ( 
.A1(n_1203),
.A2(n_1175),
.B(n_1108),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1128),
.Y(n_1596)
);

AOI22x1_ASAP7_75t_L g1597 ( 
.A1(n_1286),
.A2(n_1026),
.B1(n_1088),
.B2(n_1076),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1510),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1124),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1503),
.B(n_1030),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1155),
.Y(n_1601)
);

O2A1O1Ixp33_ASAP7_75t_L g1602 ( 
.A1(n_1130),
.A2(n_1053),
.B(n_1052),
.C(n_1063),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1287),
.B(n_1030),
.Y(n_1603)
);

AOI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1108),
.A2(n_978),
.B(n_989),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1415),
.A2(n_1088),
.B(n_1076),
.C(n_1061),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1297),
.B(n_1032),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1297),
.B(n_1032),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1381),
.A2(n_1415),
.B(n_1257),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1236),
.B(n_1406),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1200),
.A2(n_1041),
.B1(n_1076),
.B2(n_1061),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1118),
.A2(n_1039),
.B(n_989),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1265),
.B(n_1032),
.Y(n_1612)
);

AOI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1296),
.A2(n_1039),
.B(n_900),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1381),
.A2(n_1276),
.B1(n_1441),
.B2(n_1387),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1144),
.B(n_863),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1460),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1269),
.A2(n_1057),
.B(n_1041),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1265),
.B(n_1041),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1204),
.B(n_1057),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1325),
.A2(n_1061),
.B1(n_1057),
.B2(n_1101),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1359),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1287),
.B(n_873),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1279),
.B(n_266),
.Y(n_1623)
);

AOI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1274),
.A2(n_1277),
.B(n_1261),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1325),
.A2(n_1101),
.B1(n_953),
.B2(n_951),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_R g1626 ( 
.A(n_1133),
.B(n_863),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1261),
.A2(n_928),
.B(n_863),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1124),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1155),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_SL g1630 ( 
.A(n_1351),
.B(n_863),
.Y(n_1630)
);

OAI21xp33_ASAP7_75t_L g1631 ( 
.A1(n_1395),
.A2(n_110),
.B(n_109),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1414),
.A2(n_953),
.B(n_951),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1233),
.B(n_873),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1279),
.B(n_266),
.Y(n_1635)
);

OAI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1325),
.A2(n_1183),
.B1(n_1142),
.B2(n_1170),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1126),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1512),
.B(n_873),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1149),
.B(n_874),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1361),
.B(n_874),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1164),
.B(n_1364),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1414),
.A2(n_953),
.B(n_951),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1126),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_SL g1644 ( 
.A(n_1306),
.B(n_863),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1325),
.A2(n_945),
.B1(n_943),
.B2(n_935),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1278),
.A2(n_863),
.B(n_928),
.Y(n_1646)
);

NAND3xp33_ASAP7_75t_SL g1647 ( 
.A(n_1395),
.B(n_116),
.C(n_168),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_1148),
.A2(n_930),
.B(n_943),
.C(n_935),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1368),
.A2(n_945),
.B(n_943),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1501),
.A2(n_114),
.B(n_165),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1105),
.B(n_874),
.Y(n_1651)
);

INVx3_ASAP7_75t_L g1652 ( 
.A(n_1131),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1480),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1107),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1105),
.B(n_902),
.Y(n_1655)
);

AOI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1441),
.A2(n_119),
.B1(n_928),
.B2(n_164),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1119),
.B(n_902),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1119),
.B(n_902),
.Y(n_1658)
);

BUFx8_ASAP7_75t_SL g1659 ( 
.A(n_1426),
.Y(n_1659)
);

AOI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1230),
.A2(n_158),
.B1(n_155),
.B2(n_154),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1349),
.Y(n_1661)
);

A2O1A1Ixp33_ASAP7_75t_L g1662 ( 
.A1(n_1411),
.A2(n_1455),
.B(n_1368),
.C(n_1134),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1313),
.B(n_922),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1155),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1278),
.A2(n_928),
.B(n_935),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_SL g1666 ( 
.A1(n_1458),
.A2(n_130),
.B1(n_113),
.B2(n_114),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1349),
.Y(n_1667)
);

NOR3xp33_ASAP7_75t_L g1668 ( 
.A(n_1455),
.B(n_1514),
.C(n_1501),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1236),
.B(n_922),
.Y(n_1669)
);

AOI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1147),
.A2(n_945),
.B(n_934),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1306),
.B(n_266),
.Y(n_1671)
);

OAI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1167),
.A2(n_934),
.B1(n_931),
.B2(n_930),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1313),
.B(n_922),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1346),
.A2(n_934),
.B1(n_931),
.B2(n_930),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1306),
.B(n_266),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1168),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1349),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1182),
.B(n_132),
.C(n_113),
.Y(n_1678)
);

NOR2xp67_ASAP7_75t_SL g1679 ( 
.A(n_1323),
.B(n_931),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1168),
.A2(n_130),
.B1(n_116),
.B2(n_117),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1157),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1135),
.B(n_1306),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1135),
.B(n_266),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1411),
.A2(n_928),
.B(n_326),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1248),
.A2(n_928),
.B(n_322),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1255),
.B(n_266),
.Y(n_1686)
);

BUFx4f_ASAP7_75t_L g1687 ( 
.A(n_1131),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1157),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1255),
.B(n_266),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_L g1690 ( 
.A1(n_1248),
.A2(n_928),
.B(n_322),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1375),
.A2(n_928),
.B(n_322),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1244),
.B(n_266),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1244),
.B(n_272),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1171),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1246),
.B(n_272),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1359),
.B(n_1157),
.Y(n_1696)
);

BUFx6f_ASAP7_75t_L g1697 ( 
.A(n_1418),
.Y(n_1697)
);

INVx3_ASAP7_75t_SL g1698 ( 
.A(n_1236),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1246),
.B(n_272),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1375),
.A2(n_928),
.B(n_322),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1284),
.B(n_272),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1380),
.A2(n_319),
.B(n_318),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1160),
.A2(n_319),
.B(n_318),
.Y(n_1703)
);

AOI21x1_ASAP7_75t_L g1704 ( 
.A1(n_1154),
.A2(n_234),
.B(n_229),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1139),
.B(n_112),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1131),
.Y(n_1706)
);

AOI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1154),
.A2(n_234),
.B(n_229),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1139),
.B(n_117),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1420),
.B(n_272),
.Y(n_1709)
);

BUFx2_ASAP7_75t_L g1710 ( 
.A(n_1273),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1117),
.B(n_272),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1230),
.B(n_118),
.C(n_121),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1284),
.B(n_1273),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1361),
.A2(n_118),
.B(n_121),
.C(n_122),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1171),
.A2(n_135),
.B1(n_124),
.B2(n_125),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1273),
.B(n_122),
.Y(n_1716)
);

AOI21x1_ASAP7_75t_L g1717 ( 
.A1(n_1211),
.A2(n_234),
.B(n_229),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1221),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1273),
.B(n_124),
.Y(n_1719)
);

OAI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1221),
.A2(n_138),
.B1(n_126),
.B2(n_132),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1334),
.B(n_272),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1514),
.B(n_272),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1243),
.A2(n_162),
.B1(n_126),
.B2(n_133),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1159),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1334),
.B(n_125),
.Y(n_1725)
);

BUFx8_ASAP7_75t_L g1726 ( 
.A(n_1362),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1159),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1253),
.B(n_272),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1160),
.A2(n_319),
.B(n_318),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1159),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1334),
.B(n_272),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_SL g1732 ( 
.A(n_1334),
.B(n_135),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1337),
.Y(n_1733)
);

O2A1O1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1424),
.A2(n_234),
.B(n_229),
.C(n_319),
.Y(n_1734)
);

BUFx3_ASAP7_75t_L g1735 ( 
.A(n_1418),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1232),
.A2(n_1371),
.B(n_1357),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1189),
.B(n_229),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1337),
.B(n_272),
.Y(n_1738)
);

OAI22xp5_ASAP7_75t_SL g1739 ( 
.A1(n_1458),
.A2(n_163),
.B1(n_162),
.B2(n_138),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1243),
.A2(n_1250),
.B1(n_1254),
.B2(n_1245),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1366),
.Y(n_1741)
);

AO21x1_ASAP7_75t_L g1742 ( 
.A1(n_1190),
.A2(n_229),
.B(n_318),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1409),
.A2(n_163),
.B(n_229),
.C(n_319),
.Y(n_1743)
);

O2A1O1Ixp5_ASAP7_75t_L g1744 ( 
.A1(n_1114),
.A2(n_229),
.B(n_307),
.C(n_303),
.Y(n_1744)
);

NOR3xp33_ASAP7_75t_L g1745 ( 
.A(n_1133),
.B(n_229),
.C(n_208),
.Y(n_1745)
);

AOI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1232),
.A2(n_1372),
.B(n_1418),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1245),
.Y(n_1747)
);

NOR2xp33_ASAP7_75t_R g1748 ( 
.A(n_1303),
.B(n_272),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1250),
.A2(n_1260),
.B1(n_1305),
.B2(n_1254),
.Y(n_1749)
);

OAI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1260),
.A2(n_1305),
.B1(n_1376),
.B2(n_1374),
.Y(n_1750)
);

AOI22xp33_ASAP7_75t_L g1751 ( 
.A1(n_1406),
.A2(n_229),
.B1(n_289),
.B2(n_314),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1382),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1378),
.A2(n_229),
.B1(n_1),
.B2(n_2),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1418),
.A2(n_318),
.B(n_307),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1398),
.A2(n_316),
.B1(n_284),
.B2(n_200),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1337),
.B(n_282),
.Y(n_1756)
);

OAI321xp33_ASAP7_75t_L g1757 ( 
.A1(n_1425),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_8),
.C(n_9),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1253),
.B(n_282),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1222),
.B(n_282),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1496),
.A2(n_307),
.B(n_314),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1337),
.B(n_282),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1307),
.A2(n_1342),
.B1(n_1355),
.B2(n_1340),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1307),
.Y(n_1763)
);

BUFx8_ASAP7_75t_L g1764 ( 
.A(n_1362),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1189),
.B(n_206),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_SL g1766 ( 
.A1(n_1340),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_1766)
);

AOI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1496),
.A2(n_1228),
.B(n_1410),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1496),
.A2(n_307),
.B(n_314),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1323),
.A2(n_1385),
.B(n_1446),
.C(n_1437),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1496),
.A2(n_307),
.B(n_314),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1185),
.A2(n_206),
.B(n_217),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1383),
.A2(n_282),
.B(n_314),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1339),
.B(n_282),
.Y(n_1773)
);

BUFx5_ASAP7_75t_L g1774 ( 
.A(n_1413),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_SL g1775 ( 
.A(n_1133),
.B(n_10),
.Y(n_1775)
);

NOR2xp67_ASAP7_75t_L g1776 ( 
.A(n_1252),
.B(n_10),
.Y(n_1776)
);

OAI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1386),
.A2(n_206),
.B(n_217),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1252),
.B(n_11),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1106),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1189),
.B(n_206),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1191),
.B(n_206),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1191),
.B(n_282),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1356),
.A2(n_282),
.B(n_314),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1437),
.A2(n_314),
.B(n_289),
.C(n_282),
.Y(n_1784)
);

A2O1A1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1446),
.A2(n_314),
.B(n_289),
.C(n_282),
.Y(n_1785)
);

NAND2x1_ASAP7_75t_L g1786 ( 
.A(n_1131),
.B(n_282),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1339),
.B(n_1107),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_SL g1788 ( 
.A(n_1252),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1339),
.B(n_282),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1342),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1191),
.B(n_289),
.Y(n_1791)
);

NAND3xp33_ASAP7_75t_L g1792 ( 
.A(n_1225),
.B(n_314),
.C(n_289),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_1106),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1158),
.A2(n_1207),
.B(n_1338),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1220),
.A2(n_314),
.B(n_289),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1270),
.B(n_314),
.C(n_289),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1220),
.A2(n_314),
.B(n_289),
.Y(n_1797)
);

AOI21xp5_ASAP7_75t_L g1798 ( 
.A1(n_1347),
.A2(n_289),
.B(n_206),
.Y(n_1798)
);

BUFx3_ASAP7_75t_L g1799 ( 
.A(n_1362),
.Y(n_1799)
);

O2A1O1Ixp33_ASAP7_75t_L g1800 ( 
.A1(n_1393),
.A2(n_1403),
.B(n_1205),
.C(n_1115),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_SL g1801 ( 
.A(n_1339),
.B(n_289),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1112),
.A2(n_207),
.B(n_217),
.C(n_206),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1194),
.B(n_289),
.Y(n_1803)
);

NOR2xp67_ASAP7_75t_L g1804 ( 
.A(n_1252),
.B(n_13),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1347),
.A2(n_289),
.B(n_206),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1373),
.A2(n_206),
.B(n_210),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1145),
.B(n_14),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1239),
.A2(n_206),
.B(n_217),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1362),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1355),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1365),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1190),
.A2(n_1389),
.B(n_1396),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1194),
.B(n_316),
.Y(n_1813)
);

OR2x6_ASAP7_75t_L g1814 ( 
.A(n_1406),
.B(n_206),
.Y(n_1814)
);

AND2x2_ASAP7_75t_SL g1815 ( 
.A(n_1117),
.B(n_17),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1145),
.B(n_17),
.Y(n_1816)
);

INVx1_ASAP7_75t_SL g1817 ( 
.A(n_1316),
.Y(n_1817)
);

AOI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1298),
.A2(n_1433),
.B1(n_1188),
.B2(n_1475),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1440),
.B(n_1316),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1194),
.B(n_316),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1218),
.B(n_316),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1440),
.B(n_20),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1218),
.B(n_206),
.Y(n_1823)
);

BUFx6f_ASAP7_75t_L g1824 ( 
.A(n_1106),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1218),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1223),
.B(n_316),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1365),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_SL g1828 ( 
.A(n_1146),
.B(n_206),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1500),
.A2(n_316),
.B1(n_284),
.B2(n_206),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1223),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1223),
.B(n_316),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1400),
.A2(n_210),
.B(n_217),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1237),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1237),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_SL g1835 ( 
.A(n_1263),
.B(n_21),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1311),
.A2(n_210),
.B(n_217),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1237),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1241),
.A2(n_210),
.B(n_217),
.Y(n_1838)
);

INVx2_ASAP7_75t_SL g1839 ( 
.A(n_1106),
.Y(n_1839)
);

AO21x2_ASAP7_75t_L g1840 ( 
.A1(n_1211),
.A2(n_217),
.B(n_210),
.Y(n_1840)
);

AO21x1_ASAP7_75t_L g1841 ( 
.A1(n_1153),
.A2(n_208),
.B(n_217),
.Y(n_1841)
);

INVxp33_ASAP7_75t_SL g1842 ( 
.A(n_1468),
.Y(n_1842)
);

A2O1A1Ixp33_ASAP7_75t_L g1843 ( 
.A1(n_1242),
.A2(n_207),
.B(n_217),
.C(n_26),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1258),
.B(n_316),
.Y(n_1844)
);

AOI21xp5_ASAP7_75t_L g1845 ( 
.A1(n_1249),
.A2(n_210),
.B(n_207),
.Y(n_1845)
);

BUFx6f_ASAP7_75t_L g1846 ( 
.A(n_1106),
.Y(n_1846)
);

AOI21x1_ASAP7_75t_L g1847 ( 
.A1(n_1247),
.A2(n_210),
.B(n_207),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1262),
.A2(n_210),
.B(n_207),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1416),
.A2(n_210),
.B(n_208),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1146),
.B(n_208),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1258),
.B(n_316),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1369),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_1852)
);

O2A1O1Ixp33_ASAP7_75t_L g1853 ( 
.A1(n_1282),
.A2(n_210),
.B(n_31),
.C(n_33),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1484),
.B(n_1299),
.Y(n_1854)
);

A2O1A1Ixp33_ASAP7_75t_L g1855 ( 
.A1(n_1271),
.A2(n_29),
.B(n_34),
.C(n_35),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1258),
.B(n_316),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1267),
.A2(n_208),
.B(n_203),
.Y(n_1857)
);

CKINVDCx14_ASAP7_75t_R g1858 ( 
.A(n_1117),
.Y(n_1858)
);

CKINVDCx8_ASAP7_75t_R g1859 ( 
.A(n_1236),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1292),
.B(n_316),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1369),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1292),
.B(n_208),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1370),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1178),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1302),
.A2(n_208),
.B(n_203),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1292),
.B(n_316),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1321),
.B(n_316),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1321),
.B(n_316),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1208),
.B(n_1256),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1440),
.A2(n_316),
.B1(n_284),
.B2(n_208),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1178),
.Y(n_1871)
);

OAI22x1_ASAP7_75t_L g1872 ( 
.A1(n_1370),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1321),
.Y(n_1873)
);

A2O1A1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1425),
.A2(n_40),
.B(n_42),
.C(n_43),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1329),
.B(n_284),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_SL g1876 ( 
.A(n_1208),
.B(n_208),
.Y(n_1876)
);

BUFx12f_ASAP7_75t_L g1877 ( 
.A(n_1332),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_L g1878 ( 
.A1(n_1179),
.A2(n_43),
.B(n_45),
.C(n_47),
.Y(n_1878)
);

A2O1A1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1179),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1879)
);

AOI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1304),
.A2(n_208),
.B(n_203),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1256),
.B(n_230),
.Y(n_1881)
);

AO22x1_ASAP7_75t_L g1882 ( 
.A1(n_1178),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_1882)
);

AO32x1_ASAP7_75t_L g1883 ( 
.A1(n_1153),
.A2(n_55),
.A3(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_L g1884 ( 
.A(n_1440),
.B(n_56),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_SL g1885 ( 
.A(n_1236),
.B(n_230),
.Y(n_1885)
);

O2A1O1Ixp33_ASAP7_75t_L g1886 ( 
.A1(n_1317),
.A2(n_57),
.B(n_58),
.C(n_59),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1329),
.B(n_284),
.Y(n_1887)
);

AOI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1308),
.A2(n_198),
.B(n_203),
.Y(n_1888)
);

OAI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1122),
.A2(n_284),
.B(n_230),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1327),
.A2(n_198),
.B(n_203),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1332),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1310),
.B(n_230),
.Y(n_1892)
);

BUFx6f_ASAP7_75t_L g1893 ( 
.A(n_1106),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1401),
.A2(n_59),
.B(n_62),
.C(n_65),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1404),
.A2(n_284),
.B(n_233),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_SL g1896 ( 
.A(n_1310),
.B(n_230),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1377),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_SL g1898 ( 
.A(n_1263),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1327),
.A2(n_198),
.B(n_203),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_R g1900 ( 
.A(n_1384),
.B(n_67),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1329),
.B(n_67),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1330),
.B(n_68),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1402),
.B(n_68),
.Y(n_1903)
);

O2A1O1Ixp33_ASAP7_75t_L g1904 ( 
.A1(n_1193),
.A2(n_69),
.B(n_71),
.C(n_72),
.Y(n_1904)
);

AOI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1331),
.A2(n_198),
.B(n_203),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1330),
.B(n_284),
.Y(n_1906)
);

OR2x6_ASAP7_75t_SL g1907 ( 
.A(n_1367),
.B(n_69),
.Y(n_1907)
);

AOI21xp5_ASAP7_75t_L g1908 ( 
.A1(n_1331),
.A2(n_198),
.B(n_203),
.Y(n_1908)
);

OAI22xp5_ASAP7_75t_L g1909 ( 
.A1(n_1377),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1114),
.A2(n_284),
.B1(n_218),
.B2(n_230),
.Y(n_1910)
);

NAND2x1_ASAP7_75t_L g1911 ( 
.A(n_1178),
.B(n_284),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1224),
.B(n_230),
.Y(n_1912)
);

AOI21xp5_ASAP7_75t_L g1913 ( 
.A1(n_1335),
.A2(n_198),
.B(n_203),
.Y(n_1913)
);

AOI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1519),
.A2(n_1353),
.B(n_1335),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1552),
.B(n_1394),
.Y(n_1915)
);

OAI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1584),
.A2(n_1493),
.B1(n_1482),
.B2(n_1511),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1641),
.B(n_1394),
.Y(n_1917)
);

INVx4_ASAP7_75t_L g1918 ( 
.A(n_1698),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1520),
.B(n_1428),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1548),
.B(n_1428),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1549),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1528),
.B(n_1434),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1530),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1624),
.A2(n_1360),
.B(n_1353),
.Y(n_1924)
);

AOI21xp5_ASAP7_75t_L g1925 ( 
.A1(n_1585),
.A2(n_1360),
.B(n_1229),
.Y(n_1925)
);

BUFx2_ASAP7_75t_L g1926 ( 
.A(n_1710),
.Y(n_1926)
);

OAI21x1_ASAP7_75t_L g1927 ( 
.A1(n_1544),
.A2(n_1122),
.B(n_1247),
.Y(n_1927)
);

AO31x2_ASAP7_75t_L g1928 ( 
.A1(n_1517),
.A2(n_1392),
.A3(n_1184),
.B(n_1266),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1549),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_L g1930 ( 
.A(n_1608),
.B(n_1438),
.C(n_1434),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1559),
.A2(n_1229),
.B(n_1427),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1594),
.A2(n_1291),
.B(n_1266),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1621),
.B(n_1213),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1741),
.B(n_1438),
.Y(n_1934)
);

BUFx2_ASAP7_75t_SL g1935 ( 
.A(n_1859),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1752),
.B(n_1469),
.Y(n_1936)
);

OAI21x1_ASAP7_75t_L g1937 ( 
.A1(n_1812),
.A2(n_1264),
.B(n_1275),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1662),
.A2(n_1231),
.B(n_1226),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1767),
.A2(n_1264),
.B(n_1213),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1696),
.B(n_1213),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1632),
.B(n_1469),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1682),
.B(n_1479),
.Y(n_1942)
);

OA21x2_ASAP7_75t_L g1943 ( 
.A1(n_1595),
.A2(n_1392),
.B(n_1314),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1553),
.A2(n_1213),
.B(n_1312),
.Y(n_1944)
);

AOI221xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1608),
.A2(n_1184),
.B1(n_1322),
.B2(n_1508),
.C(n_1493),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1594),
.A2(n_1894),
.B(n_1769),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1538),
.B(n_1479),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1736),
.A2(n_1234),
.B(n_1508),
.Y(n_1948)
);

AOI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1646),
.A2(n_1627),
.B(n_1539),
.Y(n_1949)
);

NOR2xp67_ASAP7_75t_SL g1950 ( 
.A(n_1757),
.B(n_1263),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1525),
.B(n_1482),
.Y(n_1951)
);

AOI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1794),
.A2(n_1206),
.B(n_1216),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1543),
.B(n_1494),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1549),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1523),
.B(n_1494),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1563),
.B(n_1636),
.Y(n_1956)
);

OAI21x1_ASAP7_75t_L g1957 ( 
.A1(n_1553),
.A2(n_1670),
.B(n_1597),
.Y(n_1957)
);

O2A1O1Ixp5_ASAP7_75t_L g1958 ( 
.A1(n_1855),
.A2(n_1451),
.B(n_1474),
.C(n_1461),
.Y(n_1958)
);

A2O1A1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1668),
.A2(n_1214),
.B(n_1344),
.C(n_1497),
.Y(n_1959)
);

OAI21xp33_ASAP7_75t_L g1960 ( 
.A1(n_1631),
.A2(n_1511),
.B(n_1227),
.Y(n_1960)
);

AND2x6_ASAP7_75t_L g1961 ( 
.A(n_1609),
.B(n_1697),
.Y(n_1961)
);

OA21x2_ASAP7_75t_L g1962 ( 
.A1(n_1517),
.A2(n_1467),
.B(n_1300),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1670),
.A2(n_1309),
.B(n_1459),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1567),
.B(n_1330),
.Y(n_1964)
);

AO31x2_ASAP7_75t_L g1965 ( 
.A1(n_1565),
.A2(n_1484),
.A3(n_1358),
.B(n_1345),
.Y(n_1965)
);

AO21x1_ASAP7_75t_L g1966 ( 
.A1(n_1886),
.A2(n_1853),
.B(n_1835),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1579),
.A2(n_1290),
.B1(n_1283),
.B2(n_1280),
.Y(n_1967)
);

AO21x1_ASAP7_75t_L g1968 ( 
.A1(n_1835),
.A2(n_1196),
.B(n_1476),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1649),
.Y(n_1969)
);

A2O1A1Ixp33_ASAP7_75t_L g1970 ( 
.A1(n_1647),
.A2(n_1214),
.B(n_1235),
.C(n_1238),
.Y(n_1970)
);

A2O1A1Ixp33_ASAP7_75t_L g1971 ( 
.A1(n_1712),
.A2(n_1324),
.B(n_1326),
.C(n_1506),
.Y(n_1971)
);

INVxp67_ASAP7_75t_L g1972 ( 
.A(n_1598),
.Y(n_1972)
);

A2O1A1Ixp33_ASAP7_75t_L g1973 ( 
.A1(n_1712),
.A2(n_1436),
.B(n_1506),
.C(n_1477),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1570),
.B(n_1341),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1549),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1696),
.B(n_1621),
.Y(n_1976)
);

AO31x2_ASAP7_75t_L g1977 ( 
.A1(n_1565),
.A2(n_1397),
.A3(n_1358),
.B(n_1352),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1545),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1571),
.B(n_1341),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1666),
.B(n_1412),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1817),
.B(n_1341),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1597),
.A2(n_1459),
.B(n_1467),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1817),
.B(n_1345),
.Y(n_1983)
);

AOI21x1_ASAP7_75t_L g1984 ( 
.A1(n_1531),
.A2(n_1419),
.B(n_1315),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1590),
.B(n_1345),
.Y(n_1985)
);

BUFx10_ASAP7_75t_L g1986 ( 
.A(n_1582),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1854),
.B(n_1352),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1533),
.A2(n_1430),
.B(n_1431),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_1710),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1545),
.Y(n_1990)
);

AO31x2_ASAP7_75t_L g1991 ( 
.A1(n_1591),
.A2(n_1478),
.A3(n_1397),
.B(n_1489),
.Y(n_1991)
);

OAI21x1_ASAP7_75t_L g1992 ( 
.A1(n_1531),
.A2(n_1540),
.B(n_1556),
.Y(n_1992)
);

BUFx3_ASAP7_75t_L g1993 ( 
.A(n_1859),
.Y(n_1993)
);

A2O1A1Ixp33_ASAP7_75t_L g1994 ( 
.A1(n_1714),
.A2(n_1477),
.B(n_1436),
.C(n_1506),
.Y(n_1994)
);

BUFx2_ASAP7_75t_SL g1995 ( 
.A(n_1582),
.Y(n_1995)
);

OAI21x1_ASAP7_75t_L g1996 ( 
.A1(n_1536),
.A2(n_1315),
.B(n_1419),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1578),
.B(n_1352),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1555),
.Y(n_1998)
);

OAI21x1_ASAP7_75t_L g1999 ( 
.A1(n_1536),
.A2(n_1589),
.B(n_1746),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_SL g2000 ( 
.A(n_1636),
.B(n_1436),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1569),
.B(n_1358),
.Y(n_2001)
);

AO31x2_ASAP7_75t_L g2002 ( 
.A1(n_1591),
.A2(n_1397),
.A3(n_1478),
.B(n_1489),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1555),
.Y(n_2003)
);

OAI21x1_ASAP7_75t_L g2004 ( 
.A1(n_1564),
.A2(n_1432),
.B(n_1444),
.Y(n_2004)
);

OAI21x1_ASAP7_75t_SL g2005 ( 
.A1(n_1742),
.A2(n_1283),
.B(n_1268),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1599),
.Y(n_2006)
);

OAI21x1_ASAP7_75t_L g2007 ( 
.A1(n_1564),
.A2(n_1486),
.B(n_1491),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1854),
.B(n_1471),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_L g2009 ( 
.A1(n_1878),
.A2(n_1388),
.B(n_1492),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1750),
.B(n_1471),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1750),
.B(n_1471),
.Y(n_2011)
);

OAI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1579),
.A2(n_1268),
.B1(n_1259),
.B2(n_1280),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1616),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1603),
.B(n_1619),
.Y(n_2014)
);

AOI21xp5_ASAP7_75t_L g2015 ( 
.A1(n_1784),
.A2(n_1436),
.B(n_1506),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1599),
.Y(n_2016)
);

INVx3_ASAP7_75t_L g2017 ( 
.A(n_1609),
.Y(n_2017)
);

O2A1O1Ixp5_ASAP7_75t_L g2018 ( 
.A1(n_1879),
.A2(n_1874),
.B(n_1592),
.C(n_1568),
.Y(n_2018)
);

OAI21x1_ASAP7_75t_L g2019 ( 
.A1(n_1554),
.A2(n_1495),
.B(n_1504),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1603),
.B(n_1578),
.Y(n_2020)
);

BUFx6f_ASAP7_75t_L g2021 ( 
.A(n_1698),
.Y(n_2021)
);

A2O1A1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1566),
.A2(n_1477),
.B(n_1429),
.C(n_1384),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1649),
.Y(n_2023)
);

NOR2x1_ASAP7_75t_SL g2024 ( 
.A(n_1572),
.B(n_1187),
.Y(n_2024)
);

NOR2xp67_ASAP7_75t_L g2025 ( 
.A(n_1864),
.B(n_1477),
.Y(n_2025)
);

NAND2x1p5_ASAP7_75t_L g2026 ( 
.A(n_1687),
.B(n_1187),
.Y(n_2026)
);

HB1xp67_ASAP7_75t_L g2027 ( 
.A(n_1580),
.Y(n_2027)
);

AOI21xp5_ASAP7_75t_L g2028 ( 
.A1(n_1785),
.A2(n_1488),
.B(n_1498),
.Y(n_2028)
);

OAI21x1_ASAP7_75t_L g2029 ( 
.A1(n_1665),
.A2(n_1507),
.B(n_1453),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1666),
.B(n_1421),
.Y(n_2030)
);

INVx4_ASAP7_75t_L g2031 ( 
.A(n_1698),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1614),
.A2(n_1445),
.B(n_1452),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1622),
.B(n_1478),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1622),
.B(n_1489),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1569),
.B(n_1502),
.Y(n_2035)
);

AOI21xp5_ASAP7_75t_L g2036 ( 
.A1(n_1613),
.A2(n_1488),
.B(n_1505),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1628),
.Y(n_2037)
);

NOR2xp67_ASAP7_75t_L g2038 ( 
.A(n_1864),
.B(n_1502),
.Y(n_2038)
);

OAI21x1_ASAP7_75t_L g2039 ( 
.A1(n_1847),
.A2(n_1449),
.B(n_1448),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_1580),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1775),
.B(n_1502),
.Y(n_2041)
);

OAI21x1_ASAP7_75t_L g2042 ( 
.A1(n_1847),
.A2(n_1450),
.B(n_1442),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1663),
.B(n_1476),
.Y(n_2043)
);

NOR4xp25_ASAP7_75t_L g2044 ( 
.A(n_1757),
.B(n_1464),
.C(n_1259),
.D(n_1505),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_1739),
.B(n_1422),
.Y(n_2045)
);

A2O1A1Ixp33_ASAP7_75t_L g2046 ( 
.A1(n_1660),
.A2(n_1423),
.B(n_1443),
.C(n_1490),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1611),
.A2(n_1498),
.B(n_1417),
.Y(n_2047)
);

AOI221x1_ASAP7_75t_L g2048 ( 
.A1(n_1872),
.A2(n_1363),
.B1(n_1439),
.B2(n_1288),
.C(n_1320),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1617),
.A2(n_1417),
.B(n_1363),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1663),
.B(n_1363),
.Y(n_2050)
);

OA21x2_ASAP7_75t_L g2051 ( 
.A1(n_1744),
.A2(n_1457),
.B(n_1454),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_1575),
.B(n_1320),
.Y(n_2052)
);

NAND2x1_ASAP7_75t_L g2053 ( 
.A(n_1609),
.B(n_1320),
.Y(n_2053)
);

AOI21xp5_ASAP7_75t_L g2054 ( 
.A1(n_1626),
.A2(n_1417),
.B(n_1363),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1575),
.B(n_1320),
.Y(n_2055)
);

AOI21xp33_ASAP7_75t_L g2056 ( 
.A1(n_1753),
.A2(n_1465),
.B(n_1513),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1537),
.B(n_1320),
.Y(n_2057)
);

OAI21x1_ASAP7_75t_L g2058 ( 
.A1(n_1704),
.A2(n_1481),
.B(n_1435),
.Y(n_2058)
);

OAI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1843),
.A2(n_1499),
.B(n_1513),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1609),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1628),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1739),
.A2(n_1468),
.B1(n_1490),
.B2(n_1289),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1637),
.Y(n_2063)
);

INVx5_ASAP7_75t_L g2064 ( 
.A(n_1534),
.Y(n_2064)
);

NOR2xp33_ASAP7_75t_L g2065 ( 
.A(n_1593),
.B(n_1285),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_L g2066 ( 
.A1(n_1704),
.A2(n_1499),
.B(n_1509),
.Y(n_2066)
);

AND3x4_ASAP7_75t_L g2067 ( 
.A(n_1776),
.B(n_1490),
.C(n_1285),
.Y(n_2067)
);

OAI21x1_ASAP7_75t_L g2068 ( 
.A1(n_1707),
.A2(n_1509),
.B(n_1470),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1775),
.B(n_1187),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1707),
.A2(n_1470),
.B(n_1487),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1748),
.B(n_1187),
.Y(n_2071)
);

NAND3xp33_ASAP7_75t_L g2072 ( 
.A(n_1660),
.B(n_1485),
.C(n_1487),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1573),
.A2(n_1466),
.B(n_1472),
.Y(n_2073)
);

AOI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1626),
.A2(n_1417),
.B(n_1320),
.Y(n_2074)
);

AND2x2_ASAP7_75t_L g2075 ( 
.A(n_1569),
.B(n_1819),
.Y(n_2075)
);

AOI21x1_ASAP7_75t_L g2076 ( 
.A1(n_1679),
.A2(n_1466),
.B(n_1472),
.Y(n_2076)
);

AOI21x1_ASAP7_75t_SL g2077 ( 
.A1(n_1600),
.A2(n_1490),
.B(n_1483),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1649),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1903),
.B(n_1483),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1637),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1822),
.B(n_1288),
.Y(n_2081)
);

CKINVDCx6p67_ASAP7_75t_R g2082 ( 
.A(n_1550),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1884),
.B(n_1288),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1638),
.B(n_1288),
.Y(n_2084)
);

NOR2xp33_ASAP7_75t_L g2085 ( 
.A(n_1593),
.B(n_1288),
.Y(n_2085)
);

OAI21x1_ASAP7_75t_L g2086 ( 
.A1(n_1574),
.A2(n_1447),
.B(n_1456),
.Y(n_2086)
);

CKINVDCx20_ASAP7_75t_R g2087 ( 
.A(n_1654),
.Y(n_2087)
);

OAI21x1_ASAP7_75t_L g2088 ( 
.A1(n_1576),
.A2(n_1462),
.B(n_1463),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1547),
.B(n_1187),
.Y(n_2089)
);

AOI221xp5_ASAP7_75t_SL g2090 ( 
.A1(n_1766),
.A2(n_1515),
.B1(n_1439),
.B2(n_1363),
.C(n_1288),
.Y(n_2090)
);

INVxp67_ASAP7_75t_L g2091 ( 
.A(n_1653),
.Y(n_2091)
);

NOR2xp67_ASAP7_75t_SL g2092 ( 
.A(n_1550),
.B(n_1187),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_1542),
.A2(n_1687),
.B(n_1620),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_1864),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_1633),
.A2(n_1285),
.B(n_1439),
.Y(n_2095)
);

AO31x2_ASAP7_75t_L g2096 ( 
.A1(n_1841),
.A2(n_1742),
.A3(n_1645),
.B(n_1620),
.Y(n_2096)
);

AOI22xp5_ASAP7_75t_L g2097 ( 
.A1(n_1815),
.A2(n_1465),
.B1(n_1417),
.B2(n_1413),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1643),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_1633),
.A2(n_1439),
.B(n_1363),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1587),
.B(n_1285),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1640),
.B(n_1439),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1642),
.A2(n_1717),
.B(n_1604),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1643),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1551),
.B(n_1285),
.Y(n_2104)
);

NOR2xp33_ASAP7_75t_L g2105 ( 
.A(n_1631),
.B(n_1550),
.Y(n_2105)
);

OAI21x1_ASAP7_75t_L g2106 ( 
.A1(n_1642),
.A2(n_1439),
.B(n_1285),
.Y(n_2106)
);

BUFx6f_ASAP7_75t_L g2107 ( 
.A(n_1779),
.Y(n_2107)
);

OAI21x1_ASAP7_75t_L g2108 ( 
.A1(n_1717),
.A2(n_1473),
.B(n_1413),
.Y(n_2108)
);

OAI21x1_ASAP7_75t_L g2109 ( 
.A1(n_1684),
.A2(n_1413),
.B(n_1465),
.Y(n_2109)
);

OAI21x1_ASAP7_75t_L g2110 ( 
.A1(n_1685),
.A2(n_1413),
.B(n_284),
.Y(n_2110)
);

OA21x2_ASAP7_75t_L g2111 ( 
.A1(n_1560),
.A2(n_1413),
.B(n_75),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_L g2112 ( 
.A(n_1561),
.B(n_73),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1661),
.Y(n_2113)
);

NAND2x1p5_ASAP7_75t_L g2114 ( 
.A(n_1687),
.B(n_1413),
.Y(n_2114)
);

INVx1_ASAP7_75t_SL g2115 ( 
.A(n_1667),
.Y(n_2115)
);

INVx2_ASAP7_75t_SL g2116 ( 
.A(n_1779),
.Y(n_2116)
);

AOI21x1_ASAP7_75t_SL g2117 ( 
.A1(n_1606),
.A2(n_75),
.B(n_76),
.Y(n_2117)
);

AOI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1581),
.A2(n_198),
.B(n_212),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1562),
.B(n_77),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_1815),
.B(n_77),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1818),
.B(n_218),
.Y(n_2121)
);

AOI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1815),
.A2(n_284),
.B1(n_79),
.B2(n_80),
.Y(n_2122)
);

AOI21xp5_ASAP7_75t_L g2123 ( 
.A1(n_1588),
.A2(n_203),
.B(n_212),
.Y(n_2123)
);

AOI21xp5_ASAP7_75t_L g2124 ( 
.A1(n_1625),
.A2(n_203),
.B(n_212),
.Y(n_2124)
);

OA21x2_ASAP7_75t_L g2125 ( 
.A1(n_1560),
.A2(n_78),
.B(n_81),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1690),
.A2(n_284),
.B(n_82),
.Y(n_2126)
);

OAI21x1_ASAP7_75t_SL g2127 ( 
.A1(n_1841),
.A2(n_1800),
.B(n_1535),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1524),
.B(n_81),
.Y(n_2128)
);

OAI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_1907),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_1864),
.B(n_84),
.Y(n_2130)
);

CKINVDCx20_ASAP7_75t_R g2131 ( 
.A(n_1654),
.Y(n_2131)
);

AO31x2_ASAP7_75t_L g2132 ( 
.A1(n_1645),
.A2(n_86),
.A3(n_284),
.B(n_228),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_1691),
.A2(n_284),
.B(n_218),
.Y(n_2133)
);

BUFx3_ASAP7_75t_L g2134 ( 
.A(n_1534),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_1640),
.B(n_218),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_SL g2136 ( 
.A1(n_1516),
.A2(n_233),
.B(n_228),
.Y(n_2136)
);

NOR2x1_ASAP7_75t_L g2137 ( 
.A(n_1577),
.B(n_218),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1676),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_1871),
.B(n_218),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_1676),
.B(n_1694),
.Y(n_2140)
);

OAI21xp5_ASAP7_75t_L g2141 ( 
.A1(n_1743),
.A2(n_233),
.B(n_228),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1733),
.Y(n_2142)
);

AOI221xp5_ASAP7_75t_L g2143 ( 
.A1(n_1650),
.A2(n_218),
.B1(n_230),
.B2(n_212),
.C(n_198),
.Y(n_2143)
);

BUFx3_ASAP7_75t_L g2144 ( 
.A(n_1534),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1625),
.A2(n_198),
.B(n_203),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1700),
.A2(n_218),
.B(n_230),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_1871),
.B(n_218),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1694),
.B(n_1718),
.Y(n_2148)
);

OAI21xp5_ASAP7_75t_L g2149 ( 
.A1(n_1612),
.A2(n_233),
.B(n_228),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_1529),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1871),
.B(n_218),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_1818),
.B(n_218),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_1618),
.A2(n_233),
.B(n_228),
.Y(n_2153)
);

NOR3xp33_ASAP7_75t_L g2154 ( 
.A(n_1678),
.B(n_233),
.C(n_228),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1718),
.B(n_218),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1747),
.B(n_1763),
.Y(n_2156)
);

BUFx12f_ASAP7_75t_L g2157 ( 
.A(n_1891),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_1747),
.B(n_1763),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_1532),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_L g2160 ( 
.A1(n_1702),
.A2(n_218),
.B(n_230),
.Y(n_2160)
);

OR2x2_ASAP7_75t_L g2161 ( 
.A(n_1871),
.B(n_218),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1674),
.A2(n_1672),
.B(n_1832),
.Y(n_2162)
);

AOI21x1_ASAP7_75t_L g2163 ( 
.A1(n_1679),
.A2(n_233),
.B(n_228),
.Y(n_2163)
);

OAI21xp5_ASAP7_75t_SL g2164 ( 
.A1(n_1650),
.A2(n_218),
.B(n_230),
.Y(n_2164)
);

AO31x2_ASAP7_75t_L g2165 ( 
.A1(n_1740),
.A2(n_233),
.A3(n_228),
.B(n_218),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1795),
.A2(n_198),
.B(n_203),
.Y(n_2166)
);

AOI21xp33_ASAP7_75t_L g2167 ( 
.A1(n_1753),
.A2(n_218),
.B(n_230),
.Y(n_2167)
);

OAI21x1_ASAP7_75t_L g2168 ( 
.A1(n_1674),
.A2(n_218),
.B(n_230),
.Y(n_2168)
);

BUFx3_ASAP7_75t_L g2169 ( 
.A(n_1534),
.Y(n_2169)
);

OAI21x1_ASAP7_75t_L g2170 ( 
.A1(n_1672),
.A2(n_218),
.B(n_230),
.Y(n_2170)
);

OAI21x1_ASAP7_75t_L g2171 ( 
.A1(n_1610),
.A2(n_230),
.B(n_203),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_1610),
.A2(n_230),
.B(n_203),
.Y(n_2172)
);

OA22x2_ASAP7_75t_L g2173 ( 
.A1(n_1766),
.A2(n_230),
.B1(n_233),
.B2(n_228),
.Y(n_2173)
);

OAI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_1907),
.A2(n_230),
.B1(n_233),
.B2(n_228),
.Y(n_2174)
);

INVx1_ASAP7_75t_SL g2175 ( 
.A(n_1634),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1797),
.A2(n_198),
.B(n_203),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1607),
.A2(n_228),
.B(n_233),
.Y(n_2177)
);

OAI21x1_ASAP7_75t_L g2178 ( 
.A1(n_1889),
.A2(n_230),
.B(n_203),
.Y(n_2178)
);

OAI21x1_ASAP7_75t_L g2179 ( 
.A1(n_1889),
.A2(n_230),
.B(n_203),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_1810),
.B(n_230),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_1583),
.A2(n_198),
.B(n_203),
.Y(n_2181)
);

OAI21x1_ASAP7_75t_SL g2182 ( 
.A1(n_1516),
.A2(n_1535),
.B(n_1740),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_1659),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1810),
.B(n_198),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_1652),
.B(n_198),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_1811),
.B(n_198),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_1792),
.A2(n_198),
.B(n_203),
.Y(n_2187)
);

HB1xp67_ASAP7_75t_L g2188 ( 
.A(n_1677),
.Y(n_2188)
);

NOR2xp33_ASAP7_75t_L g2189 ( 
.A(n_1842),
.B(n_198),
.Y(n_2189)
);

BUFx6f_ASAP7_75t_L g2190 ( 
.A(n_1779),
.Y(n_2190)
);

NAND2xp33_ASAP7_75t_L g2191 ( 
.A(n_1900),
.B(n_198),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1811),
.B(n_198),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1891),
.B(n_198),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_1652),
.B(n_198),
.Y(n_2194)
);

AOI21xp5_ASAP7_75t_L g2195 ( 
.A1(n_1792),
.A2(n_203),
.B(n_212),
.Y(n_2195)
);

AOI21x1_ASAP7_75t_L g2196 ( 
.A1(n_1568),
.A2(n_228),
.B(n_233),
.Y(n_2196)
);

OAI21x1_ASAP7_75t_L g2197 ( 
.A1(n_1648),
.A2(n_1783),
.B(n_1762),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_1749),
.A2(n_212),
.B(n_228),
.Y(n_2198)
);

OA21x2_ASAP7_75t_L g2199 ( 
.A1(n_1863),
.A2(n_1897),
.B(n_1762),
.Y(n_2199)
);

AOI21x1_ASAP7_75t_L g2200 ( 
.A1(n_1615),
.A2(n_228),
.B(n_233),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_SL g2201 ( 
.A1(n_1904),
.A2(n_212),
.B(n_228),
.Y(n_2201)
);

OAI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1602),
.A2(n_228),
.B(n_233),
.Y(n_2202)
);

AOI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_1869),
.A2(n_212),
.B(n_215),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1863),
.B(n_1897),
.Y(n_2204)
);

OAI21x1_ASAP7_75t_L g2205 ( 
.A1(n_1749),
.A2(n_212),
.B(n_228),
.Y(n_2205)
);

OAI21x1_ASAP7_75t_L g2206 ( 
.A1(n_1703),
.A2(n_212),
.B(n_228),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1807),
.B(n_212),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1673),
.B(n_212),
.Y(n_2208)
);

INVxp67_ASAP7_75t_SL g2209 ( 
.A(n_1558),
.Y(n_2209)
);

INVx1_ASAP7_75t_SL g2210 ( 
.A(n_1788),
.Y(n_2210)
);

OAI21x1_ASAP7_75t_L g2211 ( 
.A1(n_1729),
.A2(n_212),
.B(n_228),
.Y(n_2211)
);

OAI21xp33_ASAP7_75t_L g2212 ( 
.A1(n_1872),
.A2(n_212),
.B(n_228),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_1652),
.B(n_212),
.Y(n_2213)
);

AOI21xp5_ASAP7_75t_L g2214 ( 
.A1(n_1796),
.A2(n_212),
.B(n_215),
.Y(n_2214)
);

OAI21x1_ASAP7_75t_L g2215 ( 
.A1(n_1786),
.A2(n_212),
.B(n_228),
.Y(n_2215)
);

OAI21xp5_ASAP7_75t_L g2216 ( 
.A1(n_1546),
.A2(n_228),
.B(n_233),
.Y(n_2216)
);

AOI211x1_ASAP7_75t_L g2217 ( 
.A1(n_1882),
.A2(n_228),
.B(n_233),
.C(n_212),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_1527),
.B(n_1713),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_L g2219 ( 
.A1(n_1786),
.A2(n_212),
.B(n_233),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1518),
.Y(n_2220)
);

AND2x2_ASAP7_75t_L g2221 ( 
.A(n_1652),
.B(n_212),
.Y(n_2221)
);

OAI22xp5_ASAP7_75t_SL g2222 ( 
.A1(n_1790),
.A2(n_233),
.B1(n_212),
.B2(n_215),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_1816),
.B(n_1705),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_1796),
.A2(n_215),
.B(n_233),
.Y(n_2224)
);

AOI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_1790),
.A2(n_215),
.B1(n_233),
.B2(n_1827),
.Y(n_2225)
);

A2O1A1Ixp33_ASAP7_75t_L g2226 ( 
.A1(n_1656),
.A2(n_215),
.B(n_233),
.C(n_1776),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1827),
.A2(n_215),
.B1(n_233),
.B2(n_1852),
.Y(n_2227)
);

OAI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_1541),
.A2(n_1852),
.B1(n_1861),
.B2(n_1909),
.Y(n_2228)
);

AOI21xp5_ASAP7_75t_L g2229 ( 
.A1(n_1644),
.A2(n_215),
.B(n_233),
.Y(n_2229)
);

OAI21x1_ASAP7_75t_L g2230 ( 
.A1(n_1838),
.A2(n_1848),
.B(n_1845),
.Y(n_2230)
);

OAI21xp5_ASAP7_75t_L g2231 ( 
.A1(n_1605),
.A2(n_215),
.B(n_1772),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1518),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1901),
.B(n_215),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1706),
.A2(n_215),
.B(n_1849),
.Y(n_2234)
);

INVx2_ASAP7_75t_SL g2235 ( 
.A(n_1779),
.Y(n_2235)
);

AO31x2_ASAP7_75t_L g2236 ( 
.A1(n_1861),
.A2(n_215),
.A3(n_1909),
.B(n_1518),
.Y(n_2236)
);

AO31x2_ASAP7_75t_L g2237 ( 
.A1(n_1521),
.A2(n_215),
.A3(n_1601),
.B(n_1596),
.Y(n_2237)
);

AOI21xp33_ASAP7_75t_L g2238 ( 
.A1(n_1722),
.A2(n_215),
.B(n_1623),
.Y(n_2238)
);

BUFx2_ASAP7_75t_L g2239 ( 
.A(n_1572),
.Y(n_2239)
);

NAND3xp33_ASAP7_75t_SL g2240 ( 
.A(n_1708),
.B(n_215),
.C(n_1680),
.Y(n_2240)
);

OAI21x1_ASAP7_75t_L g2241 ( 
.A1(n_1706),
.A2(n_215),
.B(n_1521),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_1706),
.A2(n_215),
.B(n_1521),
.Y(n_2242)
);

BUFx3_ASAP7_75t_L g2243 ( 
.A(n_1534),
.Y(n_2243)
);

OAI21x1_ASAP7_75t_L g2244 ( 
.A1(n_1706),
.A2(n_215),
.B(n_1596),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_1557),
.A2(n_215),
.B1(n_1858),
.B2(n_1715),
.Y(n_2245)
);

OAI21x1_ASAP7_75t_L g2246 ( 
.A1(n_1596),
.A2(n_215),
.B(n_1601),
.Y(n_2246)
);

OAI21x1_ASAP7_75t_L g2247 ( 
.A1(n_1601),
.A2(n_215),
.B(n_1629),
.Y(n_2247)
);

AO32x2_ASAP7_75t_L g2248 ( 
.A1(n_1883),
.A2(n_215),
.A3(n_1839),
.B1(n_1715),
.B2(n_1720),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1901),
.B(n_215),
.Y(n_2249)
);

OAI21xp5_ASAP7_75t_L g2250 ( 
.A1(n_1808),
.A2(n_1719),
.B(n_1716),
.Y(n_2250)
);

OAI21x1_ASAP7_75t_L g2251 ( 
.A1(n_1629),
.A2(n_1681),
.B(n_1664),
.Y(n_2251)
);

AO21x1_ASAP7_75t_L g2252 ( 
.A1(n_1630),
.A2(n_1883),
.B(n_1635),
.Y(n_2252)
);

AOI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_1892),
.A2(n_1896),
.B(n_1572),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_1808),
.A2(n_1732),
.B(n_1725),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1902),
.B(n_1639),
.Y(n_2255)
);

AO21x1_ASAP7_75t_L g2256 ( 
.A1(n_1883),
.A2(n_1655),
.B(n_1651),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1779),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_1572),
.A2(n_1526),
.B(n_1883),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_1582),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_SL g2260 ( 
.A(n_1778),
.B(n_1804),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1902),
.B(n_1572),
.Y(n_2261)
);

OAI21x1_ASAP7_75t_L g2262 ( 
.A1(n_1629),
.A2(n_1830),
.B(n_1730),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_1669),
.B(n_1799),
.Y(n_2263)
);

NAND2x1p5_ASAP7_75t_L g2264 ( 
.A(n_1669),
.B(n_1526),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1657),
.B(n_1658),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1664),
.Y(n_2266)
);

OAI21x1_ASAP7_75t_L g2267 ( 
.A1(n_1664),
.A2(n_1834),
.B(n_1837),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2098),
.Y(n_2268)
);

INVxp67_ASAP7_75t_L g2269 ( 
.A(n_2013),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2261),
.B(n_1940),
.Y(n_2270)
);

AND2x4_ASAP7_75t_L g2271 ( 
.A(n_2024),
.B(n_1669),
.Y(n_2271)
);

OAI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2122),
.A2(n_1778),
.B1(n_1804),
.B2(n_1787),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_1925),
.A2(n_1883),
.B(n_1882),
.Y(n_2273)
);

O2A1O1Ixp33_ASAP7_75t_SL g2274 ( 
.A1(n_2129),
.A2(n_1720),
.B(n_1723),
.C(n_1680),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2098),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_2223),
.B(n_1799),
.Y(n_2276)
);

AOI21xp5_ASAP7_75t_L g2277 ( 
.A1(n_1931),
.A2(n_1801),
.B(n_1669),
.Y(n_2277)
);

OAI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2122),
.A2(n_1735),
.B1(n_1809),
.B2(n_1799),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2098),
.Y(n_2279)
);

NOR2x1_ASAP7_75t_SL g2280 ( 
.A(n_2064),
.B(n_1840),
.Y(n_2280)
);

AO31x2_ASAP7_75t_L g2281 ( 
.A1(n_2048),
.A2(n_1837),
.A3(n_1724),
.B(n_1727),
.Y(n_2281)
);

OAI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2062),
.A2(n_1735),
.B1(n_1809),
.B2(n_1586),
.Y(n_2282)
);

INVx2_ASAP7_75t_SL g2283 ( 
.A(n_2060),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_2027),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2209),
.B(n_1681),
.Y(n_2285)
);

AND2x4_ASAP7_75t_L g2286 ( 
.A(n_2024),
.B(n_1534),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1978),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2017),
.B(n_1534),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2261),
.B(n_1840),
.Y(n_2289)
);

AOI22xp33_ASAP7_75t_L g2290 ( 
.A1(n_1956),
.A2(n_1809),
.B1(n_1814),
.B2(n_1745),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1923),
.B(n_2175),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1978),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_1940),
.B(n_1840),
.Y(n_2293)
);

INVx3_ASAP7_75t_L g2294 ( 
.A(n_2017),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1990),
.Y(n_2295)
);

O2A1O1Ixp33_ASAP7_75t_L g2296 ( 
.A1(n_2129),
.A2(n_1723),
.B(n_1689),
.C(n_1686),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1990),
.Y(n_2297)
);

A2O1A1Ixp33_ASAP7_75t_SL g2298 ( 
.A1(n_2105),
.A2(n_1701),
.B(n_1675),
.C(n_1671),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2175),
.B(n_1681),
.Y(n_2299)
);

INVxp33_ASAP7_75t_L g2300 ( 
.A(n_2065),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_1998),
.Y(n_2301)
);

NAND2x1_ASAP7_75t_L g2302 ( 
.A(n_2259),
.B(n_1688),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_2157),
.Y(n_2303)
);

CKINVDCx20_ASAP7_75t_R g2304 ( 
.A(n_2087),
.Y(n_2304)
);

BUFx3_ASAP7_75t_L g2305 ( 
.A(n_2157),
.Y(n_2305)
);

AND2x4_ASAP7_75t_L g2306 ( 
.A(n_2017),
.B(n_1839),
.Y(n_2306)
);

BUFx6f_ASAP7_75t_L g2307 ( 
.A(n_2021),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_1924),
.A2(n_1692),
.B(n_1695),
.Y(n_2308)
);

OAI22xp5_ASAP7_75t_L g2309 ( 
.A1(n_2062),
.A2(n_1735),
.B1(n_1586),
.B2(n_1755),
.Y(n_2309)
);

BUFx2_ASAP7_75t_L g2310 ( 
.A(n_2239),
.Y(n_2310)
);

OR2x2_ASAP7_75t_L g2311 ( 
.A(n_2239),
.B(n_1688),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_1976),
.B(n_1688),
.Y(n_2312)
);

AO21x2_ASAP7_75t_L g2313 ( 
.A1(n_1988),
.A2(n_1724),
.B(n_1830),
.Y(n_2313)
);

CKINVDCx20_ASAP7_75t_R g2314 ( 
.A(n_2131),
.Y(n_2314)
);

INVx4_ASAP7_75t_L g2315 ( 
.A(n_2259),
.Y(n_2315)
);

O2A1O1Ixp33_ASAP7_75t_L g2316 ( 
.A1(n_1946),
.A2(n_1709),
.B(n_1885),
.C(n_1814),
.Y(n_2316)
);

INVx4_ASAP7_75t_L g2317 ( 
.A(n_2259),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_1942),
.B(n_1724),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_1976),
.B(n_1727),
.Y(n_2319)
);

NAND2xp33_ASAP7_75t_L g2320 ( 
.A(n_1960),
.B(n_1774),
.Y(n_2320)
);

AND2x4_ASAP7_75t_L g2321 ( 
.A(n_2017),
.B(n_1793),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2094),
.B(n_1727),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_1998),
.Y(n_2323)
);

AOI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_1914),
.A2(n_1699),
.B(n_1693),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2094),
.B(n_1730),
.Y(n_2325)
);

OAI21x1_ASAP7_75t_L g2326 ( 
.A1(n_1957),
.A2(n_1873),
.B(n_1825),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_2157),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_1926),
.Y(n_2328)
);

OAI22xp33_ASAP7_75t_L g2329 ( 
.A1(n_1946),
.A2(n_1697),
.B1(n_1755),
.B2(n_1522),
.Y(n_2329)
);

NAND2x1p5_ASAP7_75t_L g2330 ( 
.A(n_2064),
.B(n_1793),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_1949),
.A2(n_1759),
.B(n_1770),
.Y(n_2331)
);

INVx4_ASAP7_75t_L g2332 ( 
.A(n_2259),
.Y(n_2332)
);

BUFx2_ASAP7_75t_L g2333 ( 
.A(n_1926),
.Y(n_2333)
);

AOI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_1932),
.A2(n_1760),
.B(n_1768),
.Y(n_2334)
);

NAND2x1p5_ASAP7_75t_L g2335 ( 
.A(n_2064),
.B(n_1793),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2040),
.B(n_1730),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2040),
.B(n_1825),
.Y(n_2337)
);

AND2x4_ASAP7_75t_L g2338 ( 
.A(n_2064),
.B(n_1793),
.Y(n_2338)
);

AND2x2_ASAP7_75t_L g2339 ( 
.A(n_2001),
.B(n_1825),
.Y(n_2339)
);

OAI22xp5_ASAP7_75t_L g2340 ( 
.A1(n_1980),
.A2(n_1586),
.B1(n_1697),
.B2(n_1522),
.Y(n_2340)
);

CKINVDCx8_ASAP7_75t_R g2341 ( 
.A(n_1935),
.Y(n_2341)
);

INVx2_ASAP7_75t_SL g2342 ( 
.A(n_2060),
.Y(n_2342)
);

BUFx2_ASAP7_75t_R g2343 ( 
.A(n_1935),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2014),
.B(n_1830),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2003),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2003),
.Y(n_2346)
);

INVx5_ASAP7_75t_L g2347 ( 
.A(n_2021),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2006),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2014),
.B(n_1833),
.Y(n_2349)
);

AO32x1_ASAP7_75t_L g2350 ( 
.A1(n_2228),
.A2(n_1834),
.A3(n_1837),
.B1(n_1833),
.B2(n_1873),
.Y(n_2350)
);

NAND2xp5_ASAP7_75t_L g2351 ( 
.A(n_2255),
.B(n_1833),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1920),
.B(n_1834),
.Y(n_2352)
);

AOI21xp5_ASAP7_75t_L g2353 ( 
.A1(n_2093),
.A2(n_1913),
.B(n_1890),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2218),
.B(n_1873),
.Y(n_2354)
);

NAND2xp5_ASAP7_75t_L g2355 ( 
.A(n_1922),
.B(n_1683),
.Y(n_2355)
);

OAI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_2030),
.A2(n_1697),
.B1(n_1522),
.B2(n_1898),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2113),
.Y(n_2357)
);

NAND2x1p5_ASAP7_75t_L g2358 ( 
.A(n_2064),
.B(n_2111),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2001),
.B(n_1793),
.Y(n_2359)
);

INVx3_ASAP7_75t_L g2360 ( 
.A(n_2060),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2064),
.B(n_1824),
.Y(n_2361)
);

NAND2xp5_ASAP7_75t_L g2362 ( 
.A(n_2265),
.B(n_1824),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2134),
.B(n_1824),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1934),
.B(n_1824),
.Y(n_2364)
);

BUFx2_ASAP7_75t_L g2365 ( 
.A(n_1989),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2006),
.Y(n_2366)
);

OAI21x1_ASAP7_75t_L g2367 ( 
.A1(n_1957),
.A2(n_1857),
.B(n_1777),
.Y(n_2367)
);

AND2x2_ASAP7_75t_L g2368 ( 
.A(n_2035),
.B(n_1824),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2016),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2035),
.B(n_1846),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2075),
.B(n_1846),
.Y(n_2371)
);

INVx4_ASAP7_75t_L g2372 ( 
.A(n_2021),
.Y(n_2372)
);

NOR2xp33_ASAP7_75t_L g2373 ( 
.A(n_2091),
.B(n_1726),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2016),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2037),
.Y(n_2375)
);

AOI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2049),
.A2(n_1899),
.B(n_1905),
.Y(n_2376)
);

INVx3_ASAP7_75t_SL g2377 ( 
.A(n_2082),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_R g2378 ( 
.A(n_2183),
.B(n_1522),
.Y(n_2378)
);

AND2x4_ASAP7_75t_L g2379 ( 
.A(n_2134),
.B(n_1846),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2057),
.B(n_1846),
.Y(n_2380)
);

INVx1_ASAP7_75t_SL g2381 ( 
.A(n_2210),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2057),
.B(n_1846),
.Y(n_2382)
);

O2A1O1Ixp5_ASAP7_75t_L g2383 ( 
.A1(n_1966),
.A2(n_1911),
.B(n_1912),
.C(n_1881),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2037),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2061),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1936),
.B(n_1893),
.Y(n_2386)
);

AOI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2071),
.A2(n_1908),
.B(n_1728),
.Y(n_2387)
);

AND2x4_ASAP7_75t_L g2388 ( 
.A(n_2134),
.B(n_1893),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_1972),
.B(n_1893),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2061),
.Y(n_2390)
);

AND2x6_ASAP7_75t_L g2391 ( 
.A(n_2144),
.B(n_1697),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2063),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2075),
.B(n_1893),
.Y(n_2393)
);

CKINVDCx5p33_ASAP7_75t_R g2394 ( 
.A(n_2082),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_1917),
.B(n_1893),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2107),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2063),
.Y(n_2397)
);

INVx5_ASAP7_75t_L g2398 ( 
.A(n_2021),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2079),
.B(n_1522),
.Y(n_2399)
);

CKINVDCx20_ASAP7_75t_R g2400 ( 
.A(n_2085),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2020),
.B(n_1774),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_2021),
.Y(n_2402)
);

INVx3_ASAP7_75t_SL g2403 ( 
.A(n_1986),
.Y(n_2403)
);

CKINVDCx20_ASAP7_75t_R g2404 ( 
.A(n_2210),
.Y(n_2404)
);

AO21x1_ASAP7_75t_L g2405 ( 
.A1(n_2228),
.A2(n_1711),
.B(n_1721),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2080),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_2080),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2103),
.Y(n_2408)
);

AND2x4_ASAP7_75t_L g2409 ( 
.A(n_2144),
.B(n_1814),
.Y(n_2409)
);

BUFx3_ASAP7_75t_L g2410 ( 
.A(n_2107),
.Y(n_2410)
);

OR2x6_ASAP7_75t_SL g2411 ( 
.A(n_1930),
.B(n_1898),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_SL g2412 ( 
.A1(n_2112),
.A2(n_1877),
.B1(n_1711),
.B2(n_1814),
.Y(n_2412)
);

AOI21xp33_ASAP7_75t_SL g2413 ( 
.A1(n_2045),
.A2(n_1711),
.B(n_1814),
.Y(n_2413)
);

INVx5_ASAP7_75t_L g2414 ( 
.A(n_2021),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2103),
.Y(n_2415)
);

INVx3_ASAP7_75t_L g2416 ( 
.A(n_2107),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2020),
.B(n_1774),
.Y(n_2417)
);

AND2x4_ASAP7_75t_L g2418 ( 
.A(n_2144),
.B(n_2169),
.Y(n_2418)
);

AOI21xp5_ASAP7_75t_L g2419 ( 
.A1(n_1930),
.A2(n_1758),
.B(n_1798),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2084),
.B(n_1823),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_1915),
.B(n_1823),
.Y(n_2421)
);

AOI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2015),
.A2(n_1805),
.B(n_1777),
.Y(n_2422)
);

O2A1O1Ixp5_ASAP7_75t_SL g2423 ( 
.A1(n_1921),
.A2(n_1876),
.B(n_1850),
.C(n_1828),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2138),
.Y(n_2424)
);

AND2x4_ASAP7_75t_L g2425 ( 
.A(n_2169),
.B(n_1911),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_1919),
.B(n_1781),
.Y(n_2426)
);

BUFx6f_ASAP7_75t_L g2427 ( 
.A(n_1986),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_1941),
.B(n_1964),
.Y(n_2428)
);

BUFx2_ASAP7_75t_L g2429 ( 
.A(n_1989),
.Y(n_2429)
);

CKINVDCx5p33_ASAP7_75t_R g2430 ( 
.A(n_1995),
.Y(n_2430)
);

AOI21xp5_ASAP7_75t_L g2431 ( 
.A1(n_1952),
.A2(n_1754),
.B(n_1731),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1955),
.B(n_1781),
.Y(n_2432)
);

BUFx3_ASAP7_75t_L g2433 ( 
.A(n_2107),
.Y(n_2433)
);

NAND2x1p5_ASAP7_75t_L g2434 ( 
.A(n_2111),
.B(n_1774),
.Y(n_2434)
);

OAI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_2067),
.A2(n_1898),
.B1(n_1829),
.B2(n_1877),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2138),
.B(n_1774),
.Y(n_2436)
);

OAI21xp5_ASAP7_75t_L g2437 ( 
.A1(n_2018),
.A2(n_1789),
.B(n_1773),
.Y(n_2437)
);

A2O1A1Ixp33_ASAP7_75t_L g2438 ( 
.A1(n_1960),
.A2(n_1761),
.B(n_1738),
.C(n_1756),
.Y(n_2438)
);

AND2x4_ASAP7_75t_L g2439 ( 
.A(n_2169),
.B(n_1765),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2115),
.B(n_1780),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_2107),
.Y(n_2441)
);

INVx4_ASAP7_75t_L g2442 ( 
.A(n_1986),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2199),
.Y(n_2443)
);

INVx4_ASAP7_75t_L g2444 ( 
.A(n_1986),
.Y(n_2444)
);

INVx6_ASAP7_75t_L g2445 ( 
.A(n_1918),
.Y(n_2445)
);

AOI21xp5_ASAP7_75t_L g2446 ( 
.A1(n_2047),
.A2(n_1966),
.B(n_2041),
.Y(n_2446)
);

BUFx2_ASAP7_75t_L g2447 ( 
.A(n_2199),
.Y(n_2447)
);

INVx4_ASAP7_75t_L g2448 ( 
.A(n_1918),
.Y(n_2448)
);

INVx2_ASAP7_75t_SL g2449 ( 
.A(n_2115),
.Y(n_2449)
);

INVx3_ASAP7_75t_L g2450 ( 
.A(n_2107),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1947),
.B(n_1780),
.Y(n_2451)
);

INVx1_ASAP7_75t_SL g2452 ( 
.A(n_2052),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2089),
.B(n_1765),
.Y(n_2453)
);

BUFx4f_ASAP7_75t_L g2454 ( 
.A(n_2067),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1953),
.B(n_1726),
.Y(n_2455)
);

INVx1_ASAP7_75t_L g2456 ( 
.A(n_2199),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_1933),
.B(n_1774),
.Y(n_2457)
);

OAI321xp33_ASAP7_75t_L g2458 ( 
.A1(n_2120),
.A2(n_1870),
.A3(n_1771),
.B1(n_1829),
.B2(n_1895),
.C(n_1737),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2207),
.B(n_1726),
.Y(n_2459)
);

AOI22xp33_ASAP7_75t_L g2460 ( 
.A1(n_2120),
.A2(n_1726),
.B1(n_1764),
.B2(n_1877),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_2190),
.Y(n_2461)
);

INVx2_ASAP7_75t_SL g2462 ( 
.A(n_2190),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2199),
.Y(n_2463)
);

BUFx12f_ASAP7_75t_L g2464 ( 
.A(n_2130),
.Y(n_2464)
);

AND2x2_ASAP7_75t_L g2465 ( 
.A(n_1933),
.B(n_1774),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1951),
.B(n_1764),
.Y(n_2466)
);

BUFx6f_ASAP7_75t_L g2467 ( 
.A(n_2190),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2243),
.B(n_1737),
.Y(n_2468)
);

OAI22xp5_ASAP7_75t_L g2469 ( 
.A1(n_2067),
.A2(n_1870),
.B1(n_1751),
.B2(n_1910),
.Y(n_2469)
);

A2O1A1Ixp33_ASAP7_75t_L g2470 ( 
.A1(n_2090),
.A2(n_1734),
.B(n_1806),
.C(n_1895),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2140),
.Y(n_2471)
);

OR2x6_ASAP7_75t_L g2472 ( 
.A(n_1995),
.B(n_1774),
.Y(n_2472)
);

AOI21xp5_ASAP7_75t_SL g2473 ( 
.A1(n_2069),
.A2(n_1764),
.B(n_1771),
.Y(n_2473)
);

OAI22xp5_ASAP7_75t_L g2474 ( 
.A1(n_2097),
.A2(n_1851),
.B1(n_1887),
.B2(n_1875),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2100),
.B(n_1764),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2101),
.B(n_1774),
.Y(n_2476)
);

AND2x2_ASAP7_75t_SL g2477 ( 
.A(n_2111),
.B(n_1862),
.Y(n_2477)
);

OAI21xp33_ASAP7_75t_L g2478 ( 
.A1(n_2128),
.A2(n_1844),
.B(n_1868),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2190),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2140),
.Y(n_2480)
);

AO21x2_ASAP7_75t_L g2481 ( 
.A1(n_1938),
.A2(n_1836),
.B(n_1888),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2148),
.Y(n_2482)
);

BUFx4_ASAP7_75t_SL g2483 ( 
.A(n_1993),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2267),
.Y(n_2484)
);

OR2x6_ASAP7_75t_L g2485 ( 
.A(n_2114),
.B(n_1782),
.Y(n_2485)
);

HB1xp67_ASAP7_75t_L g2486 ( 
.A(n_2142),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2081),
.B(n_1856),
.Y(n_2487)
);

O2A1O1Ixp5_ASAP7_75t_L g2488 ( 
.A1(n_1968),
.A2(n_1950),
.B(n_2260),
.C(n_2000),
.Y(n_2488)
);

AOI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2054),
.A2(n_2074),
.B(n_1971),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2174),
.B(n_1802),
.C(n_1831),
.Y(n_2490)
);

O2A1O1Ixp33_ASAP7_75t_L g2491 ( 
.A1(n_1967),
.A2(n_1906),
.B(n_1860),
.C(n_1813),
.Y(n_2491)
);

AOI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2036),
.A2(n_1791),
.B(n_1803),
.Y(n_2492)
);

BUFx3_ASAP7_75t_L g2493 ( 
.A(n_2190),
.Y(n_2493)
);

NAND2x1_ASAP7_75t_L g2494 ( 
.A(n_1918),
.B(n_1862),
.Y(n_2494)
);

HB1xp67_ASAP7_75t_L g2495 ( 
.A(n_2188),
.Y(n_2495)
);

OR2x2_ASAP7_75t_L g2496 ( 
.A(n_1965),
.B(n_1820),
.Y(n_2496)
);

NOR2x1_ASAP7_75t_R g2497 ( 
.A(n_1918),
.B(n_1821),
.Y(n_2497)
);

AND2x4_ASAP7_75t_L g2498 ( 
.A(n_2243),
.B(n_1826),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2267),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2190),
.Y(n_2500)
);

NOR2xp33_ASAP7_75t_SL g2501 ( 
.A(n_2031),
.B(n_1866),
.Y(n_2501)
);

AND2x4_ASAP7_75t_L g2502 ( 
.A(n_2243),
.B(n_1867),
.Y(n_2502)
);

AO21x1_ASAP7_75t_L g2503 ( 
.A1(n_1916),
.A2(n_1865),
.B(n_1880),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_1973),
.A2(n_1938),
.B(n_2022),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2148),
.Y(n_2505)
);

BUFx3_ASAP7_75t_L g2506 ( 
.A(n_2257),
.Y(n_2506)
);

INVx3_ASAP7_75t_L g2507 ( 
.A(n_2257),
.Y(n_2507)
);

BUFx6f_ASAP7_75t_L g2508 ( 
.A(n_2257),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_2104),
.B(n_2159),
.Y(n_2509)
);

INVx2_ASAP7_75t_L g2510 ( 
.A(n_2251),
.Y(n_2510)
);

CKINVDCx8_ASAP7_75t_R g2511 ( 
.A(n_1961),
.Y(n_2511)
);

BUFx6f_ASAP7_75t_L g2512 ( 
.A(n_2257),
.Y(n_2512)
);

BUFx6f_ASAP7_75t_L g2513 ( 
.A(n_2257),
.Y(n_2513)
);

AOI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2028),
.A2(n_1970),
.B(n_2048),
.Y(n_2514)
);

AND2x4_ASAP7_75t_L g2515 ( 
.A(n_2263),
.B(n_2095),
.Y(n_2515)
);

BUFx2_ASAP7_75t_L g2516 ( 
.A(n_2095),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_1965),
.B(n_2101),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2099),
.Y(n_2518)
);

AOI21xp5_ASAP7_75t_L g2519 ( 
.A1(n_2197),
.A2(n_1968),
.B(n_2253),
.Y(n_2519)
);

BUFx3_ASAP7_75t_L g2520 ( 
.A(n_2257),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_SL g2521 ( 
.A(n_1967),
.B(n_2012),
.Y(n_2521)
);

OA21x2_ASAP7_75t_L g2522 ( 
.A1(n_1999),
.A2(n_1992),
.B(n_1927),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2053),
.Y(n_2523)
);

AND2x6_ASAP7_75t_L g2524 ( 
.A(n_1993),
.B(n_2097),
.Y(n_2524)
);

AOI21xp5_ASAP7_75t_L g2525 ( 
.A1(n_2197),
.A2(n_1948),
.B(n_1994),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2053),
.Y(n_2526)
);

INVx3_ASAP7_75t_L g2527 ( 
.A(n_1961),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2156),
.Y(n_2528)
);

AOI22xp33_ASAP7_75t_SL g2529 ( 
.A1(n_2182),
.A2(n_2127),
.B1(n_2012),
.B2(n_2174),
.Y(n_2529)
);

AOI21xp5_ASAP7_75t_L g2530 ( 
.A1(n_1948),
.A2(n_2111),
.B(n_2032),
.Y(n_2530)
);

CKINVDCx8_ASAP7_75t_R g2531 ( 
.A(n_1961),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_1965),
.B(n_2263),
.Y(n_2532)
);

OA21x2_ASAP7_75t_L g2533 ( 
.A1(n_1999),
.A2(n_1992),
.B(n_1927),
.Y(n_2533)
);

AOI22xp5_ASAP7_75t_L g2534 ( 
.A1(n_2240),
.A2(n_2090),
.B1(n_2245),
.B2(n_1950),
.Y(n_2534)
);

AOI21xp5_ASAP7_75t_L g2535 ( 
.A1(n_1948),
.A2(n_2032),
.B(n_2046),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2156),
.Y(n_2536)
);

OR2x2_ASAP7_75t_L g2537 ( 
.A(n_1965),
.B(n_1921),
.Y(n_2537)
);

INVx4_ASAP7_75t_L g2538 ( 
.A(n_2031),
.Y(n_2538)
);

AND2x4_ASAP7_75t_L g2539 ( 
.A(n_2263),
.B(n_2099),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_L g2540 ( 
.A(n_2159),
.B(n_1987),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_1993),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2106),
.Y(n_2542)
);

A2O1A1Ixp33_ASAP7_75t_L g2543 ( 
.A1(n_2191),
.A2(n_2201),
.B(n_2254),
.C(n_2250),
.Y(n_2543)
);

AND2x2_ASAP7_75t_L g2544 ( 
.A(n_1965),
.B(n_2263),
.Y(n_2544)
);

NOR2xp33_ASAP7_75t_SL g2545 ( 
.A(n_2031),
.B(n_2092),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_1987),
.B(n_2008),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2158),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_1948),
.A2(n_2073),
.B(n_1943),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2008),
.B(n_2052),
.Y(n_2549)
);

AOI21xp5_ASAP7_75t_L g2550 ( 
.A1(n_2073),
.A2(n_1943),
.B(n_2044),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_L g2551 ( 
.A(n_2055),
.B(n_2083),
.Y(n_2551)
);

OAI22xp5_ASAP7_75t_L g2552 ( 
.A1(n_2072),
.A2(n_2227),
.B1(n_2114),
.B2(n_2150),
.Y(n_2552)
);

OR2x2_ASAP7_75t_SL g2553 ( 
.A(n_2125),
.B(n_1943),
.Y(n_2553)
);

OAI22xp5_ASAP7_75t_L g2554 ( 
.A1(n_2072),
.A2(n_2227),
.B1(n_2114),
.B2(n_2150),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2158),
.Y(n_2555)
);

NAND2x1p5_ASAP7_75t_L g2556 ( 
.A(n_2031),
.B(n_2092),
.Y(n_2556)
);

HB1xp67_ASAP7_75t_L g2557 ( 
.A(n_1997),
.Y(n_2557)
);

NAND2xp5_ASAP7_75t_L g2558 ( 
.A(n_2055),
.B(n_2043),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2251),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2262),
.Y(n_2560)
);

AOI21xp5_ASAP7_75t_L g2561 ( 
.A1(n_1943),
.A2(n_2044),
.B(n_2250),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2262),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_SL g2563 ( 
.A(n_2254),
.B(n_2119),
.Y(n_2563)
);

OAI22xp5_ASAP7_75t_L g2564 ( 
.A1(n_2225),
.A2(n_2201),
.B1(n_1959),
.B2(n_2245),
.Y(n_2564)
);

NOR2xp33_ASAP7_75t_L g2565 ( 
.A(n_2189),
.B(n_2050),
.Y(n_2565)
);

OAI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2226),
.A2(n_2203),
.B(n_2229),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2204),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2043),
.B(n_1981),
.Y(n_2568)
);

INVx3_ASAP7_75t_SL g2569 ( 
.A(n_2116),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_L g2570 ( 
.A1(n_2182),
.A2(n_2009),
.B(n_2127),
.Y(n_2570)
);

INVx2_ASAP7_75t_L g2571 ( 
.A(n_2220),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2204),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_1929),
.Y(n_2573)
);

OAI22xp5_ASAP7_75t_SL g2574 ( 
.A1(n_2125),
.A2(n_2026),
.B1(n_2264),
.B2(n_1916),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_1929),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2026),
.A2(n_2173),
.B1(n_2212),
.B2(n_1985),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_1954),
.Y(n_2577)
);

AOI21xp5_ASAP7_75t_L g2578 ( 
.A1(n_2009),
.A2(n_1958),
.B(n_2059),
.Y(n_2578)
);

BUFx3_ASAP7_75t_L g2579 ( 
.A(n_1961),
.Y(n_2579)
);

INVx1_ASAP7_75t_SL g2580 ( 
.A(n_2050),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2059),
.A2(n_2125),
.B(n_2011),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_1983),
.B(n_1985),
.Y(n_2582)
);

INVx2_ASAP7_75t_SL g2583 ( 
.A(n_2116),
.Y(n_2583)
);

OAI22xp5_ASAP7_75t_L g2584 ( 
.A1(n_2026),
.A2(n_2173),
.B1(n_2212),
.B2(n_2264),
.Y(n_2584)
);

INVxp67_ASAP7_75t_L g2585 ( 
.A(n_2033),
.Y(n_2585)
);

AND2x4_ASAP7_75t_L g2586 ( 
.A(n_2106),
.B(n_1961),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_1954),
.Y(n_2587)
);

AND2x4_ASAP7_75t_L g2588 ( 
.A(n_1961),
.B(n_2220),
.Y(n_2588)
);

INVx1_ASAP7_75t_SL g2589 ( 
.A(n_1997),
.Y(n_2589)
);

BUFx6f_ASAP7_75t_L g2590 ( 
.A(n_1961),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_1974),
.B(n_1979),
.Y(n_2591)
);

OAI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2238),
.A2(n_2126),
.B(n_2241),
.Y(n_2592)
);

AOI22xp5_ASAP7_75t_L g2593 ( 
.A1(n_2173),
.A2(n_2222),
.B1(n_2154),
.B2(n_1945),
.Y(n_2593)
);

OAI21xp5_ASAP7_75t_L g2594 ( 
.A1(n_2238),
.A2(n_2126),
.B(n_2241),
.Y(n_2594)
);

BUFx6f_ASAP7_75t_L g2595 ( 
.A(n_2264),
.Y(n_2595)
);

AOI21xp5_ASAP7_75t_L g2596 ( 
.A1(n_2125),
.A2(n_2011),
.B(n_2010),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_2033),
.B(n_2034),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_1965),
.B(n_2130),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_1975),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2232),
.Y(n_2600)
);

AOI22xp5_ASAP7_75t_L g2601 ( 
.A1(n_2222),
.A2(n_1945),
.B1(n_2152),
.B2(n_2121),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_2034),
.B(n_2010),
.Y(n_2602)
);

CKINVDCx16_ASAP7_75t_R g2603 ( 
.A(n_2235),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2213),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2235),
.Y(n_2605)
);

AOI21xp5_ASAP7_75t_L g2606 ( 
.A1(n_1939),
.A2(n_2019),
.B(n_2102),
.Y(n_2606)
);

NAND2x1p5_ASAP7_75t_L g2607 ( 
.A(n_2102),
.B(n_1939),
.Y(n_2607)
);

HB1xp67_ASAP7_75t_L g2608 ( 
.A(n_2038),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2242),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2232),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1975),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2266),
.Y(n_2612)
);

BUFx6f_ASAP7_75t_L g2613 ( 
.A(n_2242),
.Y(n_2613)
);

CKINVDCx11_ASAP7_75t_R g2614 ( 
.A(n_2266),
.Y(n_2614)
);

AOI21xp5_ASAP7_75t_L g2615 ( 
.A1(n_2019),
.A2(n_2029),
.B(n_2056),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_1991),
.B(n_2002),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_1991),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_2135),
.B(n_2038),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2025),
.B(n_1991),
.Y(n_2619)
);

AO21x1_ASAP7_75t_L g2620 ( 
.A1(n_2258),
.A2(n_2056),
.B(n_2076),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_1991),
.Y(n_2621)
);

OAI22xp5_ASAP7_75t_L g2622 ( 
.A1(n_2193),
.A2(n_2164),
.B1(n_2217),
.B2(n_2025),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_1991),
.Y(n_2623)
);

AND2x4_ASAP7_75t_L g2624 ( 
.A(n_1991),
.B(n_2002),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2002),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2454),
.A2(n_2217),
.B1(n_2164),
.B2(n_2249),
.Y(n_2626)
);

BUFx2_ASAP7_75t_L g2627 ( 
.A(n_2515),
.Y(n_2627)
);

OAI22xp5_ASAP7_75t_L g2628 ( 
.A1(n_2454),
.A2(n_2233),
.B1(n_2149),
.B2(n_2153),
.Y(n_2628)
);

BUFx6f_ASAP7_75t_L g2629 ( 
.A(n_2427),
.Y(n_2629)
);

AOI22xp33_ASAP7_75t_L g2630 ( 
.A1(n_2521),
.A2(n_2136),
.B1(n_2177),
.B2(n_2149),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2573),
.Y(n_2631)
);

INVx6_ASAP7_75t_L g2632 ( 
.A(n_2347),
.Y(n_2632)
);

AOI22xp33_ASAP7_75t_L g2633 ( 
.A1(n_2564),
.A2(n_2136),
.B1(n_2177),
.B2(n_2153),
.Y(n_2633)
);

BUFx3_ASAP7_75t_L g2634 ( 
.A(n_2526),
.Y(n_2634)
);

AOI22xp33_ASAP7_75t_L g2635 ( 
.A1(n_2566),
.A2(n_2216),
.B1(n_2202),
.B2(n_2252),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2274),
.A2(n_2252),
.B1(n_2216),
.B2(n_2202),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2573),
.Y(n_2637)
);

BUFx10_ASAP7_75t_L g2638 ( 
.A(n_2394),
.Y(n_2638)
);

INVx3_ASAP7_75t_SL g2639 ( 
.A(n_2394),
.Y(n_2639)
);

BUFx6f_ASAP7_75t_L g2640 ( 
.A(n_2427),
.Y(n_2640)
);

INVx1_ASAP7_75t_SL g2641 ( 
.A(n_2328),
.Y(n_2641)
);

BUFx4_ASAP7_75t_R g2642 ( 
.A(n_2303),
.Y(n_2642)
);

OAI22xp5_ASAP7_75t_L g2643 ( 
.A1(n_2454),
.A2(n_2135),
.B1(n_2137),
.B2(n_2200),
.Y(n_2643)
);

OAI22xp5_ASAP7_75t_L g2644 ( 
.A1(n_2290),
.A2(n_2137),
.B1(n_2200),
.B2(n_2214),
.Y(n_2644)
);

AOI22xp33_ASAP7_75t_SL g2645 ( 
.A1(n_2524),
.A2(n_2117),
.B1(n_2005),
.B2(n_2231),
.Y(n_2645)
);

BUFx8_ASAP7_75t_L g2646 ( 
.A(n_2427),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_2552),
.A2(n_2256),
.B1(n_2234),
.B2(n_2244),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2515),
.Y(n_2648)
);

OAI21xp33_ASAP7_75t_L g2649 ( 
.A1(n_2563),
.A2(n_2076),
.B(n_2231),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2524),
.A2(n_2234),
.B1(n_2141),
.B2(n_2244),
.Y(n_2650)
);

OAI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2543),
.A2(n_2180),
.B1(n_2155),
.B2(n_2194),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2291),
.B(n_2551),
.Y(n_2652)
);

OAI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2341),
.A2(n_2180),
.B1(n_2155),
.B2(n_2194),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2575),
.Y(n_2654)
);

OAI22xp33_ASAP7_75t_SL g2655 ( 
.A1(n_2411),
.A2(n_2248),
.B1(n_2185),
.B2(n_2132),
.Y(n_2655)
);

INVx6_ASAP7_75t_L g2656 ( 
.A(n_2347),
.Y(n_2656)
);

OAI22xp5_ASAP7_75t_L g2657 ( 
.A1(n_2341),
.A2(n_2185),
.B1(n_2141),
.B2(n_2208),
.Y(n_2657)
);

INVx1_ASAP7_75t_SL g2658 ( 
.A(n_2328),
.Y(n_2658)
);

BUFx8_ASAP7_75t_L g2659 ( 
.A(n_2427),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2524),
.A2(n_2205),
.B1(n_2198),
.B2(n_2005),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2575),
.Y(n_2661)
);

INVx2_ASAP7_75t_SL g2662 ( 
.A(n_2347),
.Y(n_2662)
);

OAI21xp33_ASAP7_75t_L g2663 ( 
.A1(n_2578),
.A2(n_1969),
.B(n_2023),
.Y(n_2663)
);

INVxp33_ASAP7_75t_L g2664 ( 
.A(n_2378),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2577),
.Y(n_2665)
);

AOI22xp33_ASAP7_75t_L g2666 ( 
.A1(n_2524),
.A2(n_2205),
.B1(n_2198),
.B2(n_2256),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2577),
.Y(n_2667)
);

CKINVDCx11_ASAP7_75t_R g2668 ( 
.A(n_2304),
.Y(n_2668)
);

INVx6_ASAP7_75t_L g2669 ( 
.A(n_2347),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2587),
.Y(n_2670)
);

AOI22xp33_ASAP7_75t_L g2671 ( 
.A1(n_2524),
.A2(n_2246),
.B1(n_2247),
.B2(n_2167),
.Y(n_2671)
);

AOI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2524),
.A2(n_2246),
.B1(n_2247),
.B2(n_2167),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2587),
.Y(n_2673)
);

BUFx12f_ASAP7_75t_L g2674 ( 
.A(n_2430),
.Y(n_2674)
);

AOI22xp33_ASAP7_75t_L g2675 ( 
.A1(n_2524),
.A2(n_2221),
.B1(n_2213),
.B2(n_2211),
.Y(n_2675)
);

CKINVDCx11_ASAP7_75t_R g2676 ( 
.A(n_2314),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_2490),
.A2(n_2221),
.B1(n_2206),
.B2(n_2211),
.Y(n_2677)
);

INVx8_ASAP7_75t_L g2678 ( 
.A(n_2391),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2599),
.Y(n_2679)
);

AOI22xp33_ASAP7_75t_SL g2680 ( 
.A1(n_2412),
.A2(n_2272),
.B1(n_2504),
.B2(n_2554),
.Y(n_2680)
);

BUFx6f_ASAP7_75t_L g2681 ( 
.A(n_2427),
.Y(n_2681)
);

AND2x2_ASAP7_75t_L g2682 ( 
.A(n_2270),
.B(n_2532),
.Y(n_2682)
);

BUFx3_ASAP7_75t_L g2683 ( 
.A(n_2526),
.Y(n_2683)
);

AO22x1_ASAP7_75t_L g2684 ( 
.A1(n_2430),
.A2(n_2078),
.B1(n_2023),
.B2(n_1969),
.Y(n_2684)
);

AOI22xp5_ASAP7_75t_L g2685 ( 
.A1(n_2329),
.A2(n_2088),
.B1(n_2086),
.B2(n_2109),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_SL g2686 ( 
.A1(n_2412),
.A2(n_2162),
.B1(n_2248),
.B2(n_2109),
.Y(n_2686)
);

AOI22xp33_ASAP7_75t_L g2687 ( 
.A1(n_2529),
.A2(n_2206),
.B1(n_2224),
.B2(n_2230),
.Y(n_2687)
);

CKINVDCx11_ASAP7_75t_R g2688 ( 
.A(n_2404),
.Y(n_2688)
);

INVx1_ASAP7_75t_SL g2689 ( 
.A(n_2333),
.Y(n_2689)
);

INVx6_ASAP7_75t_L g2690 ( 
.A(n_2347),
.Y(n_2690)
);

NAND2xp5_ASAP7_75t_L g2691 ( 
.A(n_2568),
.B(n_2002),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2526),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_2405),
.A2(n_2230),
.B1(n_2051),
.B2(n_2215),
.Y(n_2693)
);

OAI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2411),
.A2(n_2208),
.B1(n_2196),
.B2(n_2184),
.Y(n_2694)
);

CKINVDCx11_ASAP7_75t_R g2695 ( 
.A(n_2377),
.Y(n_2695)
);

BUFx2_ASAP7_75t_L g2696 ( 
.A(n_2515),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2515),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2599),
.Y(n_2698)
);

AOI22xp33_ASAP7_75t_L g2699 ( 
.A1(n_2498),
.A2(n_2051),
.B1(n_2215),
.B2(n_2219),
.Y(n_2699)
);

INVxp67_ASAP7_75t_SL g2700 ( 
.A(n_2608),
.Y(n_2700)
);

CKINVDCx11_ASAP7_75t_R g2701 ( 
.A(n_2377),
.Y(n_2701)
);

INVx3_ASAP7_75t_L g2702 ( 
.A(n_2539),
.Y(n_2702)
);

INVx4_ASAP7_75t_L g2703 ( 
.A(n_2403),
.Y(n_2703)
);

AOI22xp33_ASAP7_75t_L g2704 ( 
.A1(n_2498),
.A2(n_2051),
.B1(n_2219),
.B2(n_2110),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2611),
.Y(n_2705)
);

AOI22xp33_ASAP7_75t_L g2706 ( 
.A1(n_2498),
.A2(n_2051),
.B1(n_2110),
.B2(n_2151),
.Y(n_2706)
);

AOI22xp33_ASAP7_75t_L g2707 ( 
.A1(n_2502),
.A2(n_2139),
.B1(n_2151),
.B2(n_2088),
.Y(n_2707)
);

AOI22xp33_ASAP7_75t_SL g2708 ( 
.A1(n_2570),
.A2(n_2162),
.B1(n_2248),
.B2(n_1962),
.Y(n_2708)
);

AOI22xp33_ASAP7_75t_L g2709 ( 
.A1(n_2502),
.A2(n_2613),
.B1(n_2609),
.B2(n_2464),
.Y(n_2709)
);

INVx2_ASAP7_75t_L g2710 ( 
.A(n_2611),
.Y(n_2710)
);

OAI22xp5_ASAP7_75t_L g2711 ( 
.A1(n_2534),
.A2(n_2196),
.B1(n_2186),
.B2(n_2184),
.Y(n_2711)
);

INVx6_ASAP7_75t_L g2712 ( 
.A(n_2347),
.Y(n_2712)
);

OAI22xp33_ASAP7_75t_L g2713 ( 
.A1(n_2534),
.A2(n_2192),
.B1(n_2186),
.B2(n_2161),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2287),
.Y(n_2714)
);

OAI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2446),
.A2(n_1944),
.B(n_2029),
.Y(n_2715)
);

AOI22xp33_ASAP7_75t_L g2716 ( 
.A1(n_2502),
.A2(n_2139),
.B1(n_2086),
.B2(n_1962),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2279),
.Y(n_2717)
);

AOI22xp33_ASAP7_75t_L g2718 ( 
.A1(n_2609),
.A2(n_1962),
.B1(n_2124),
.B2(n_2145),
.Y(n_2718)
);

OAI22xp33_ASAP7_75t_L g2719 ( 
.A1(n_2601),
.A2(n_2192),
.B1(n_2147),
.B2(n_2161),
.Y(n_2719)
);

INVx3_ASAP7_75t_L g2720 ( 
.A(n_2539),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_L g2721 ( 
.A1(n_2609),
.A2(n_1962),
.B1(n_2023),
.B2(n_2078),
.Y(n_2721)
);

INVx8_ASAP7_75t_L g2722 ( 
.A(n_2391),
.Y(n_2722)
);

AOI22xp33_ASAP7_75t_L g2723 ( 
.A1(n_2609),
.A2(n_1969),
.B1(n_2078),
.B2(n_2123),
.Y(n_2723)
);

OAI22xp5_ASAP7_75t_SL g2724 ( 
.A1(n_2400),
.A2(n_2248),
.B1(n_1928),
.B2(n_2132),
.Y(n_2724)
);

AND2x2_ASAP7_75t_L g2725 ( 
.A(n_2270),
.B(n_1977),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2287),
.Y(n_2726)
);

BUFx2_ASAP7_75t_L g2727 ( 
.A(n_2539),
.Y(n_2727)
);

INVx2_ASAP7_75t_L g2728 ( 
.A(n_2279),
.Y(n_2728)
);

BUFx2_ASAP7_75t_L g2729 ( 
.A(n_2539),
.Y(n_2729)
);

BUFx10_ASAP7_75t_L g2730 ( 
.A(n_2445),
.Y(n_2730)
);

BUFx12f_ASAP7_75t_L g2731 ( 
.A(n_2614),
.Y(n_2731)
);

AOI22xp33_ASAP7_75t_L g2732 ( 
.A1(n_2609),
.A2(n_2118),
.B1(n_2058),
.B2(n_1944),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2469),
.A2(n_2108),
.B1(n_2066),
.B2(n_2068),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2268),
.Y(n_2734)
);

INVx2_ASAP7_75t_L g2735 ( 
.A(n_2268),
.Y(n_2735)
);

OAI22xp33_ASAP7_75t_L g2736 ( 
.A1(n_2601),
.A2(n_2147),
.B1(n_2163),
.B2(n_2077),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2292),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2275),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2275),
.Y(n_2739)
);

AOI22xp33_ASAP7_75t_L g2740 ( 
.A1(n_2613),
.A2(n_2058),
.B1(n_2166),
.B2(n_2176),
.Y(n_2740)
);

AOI22xp33_ASAP7_75t_L g2741 ( 
.A1(n_2613),
.A2(n_2108),
.B1(n_2066),
.B2(n_2039),
.Y(n_2741)
);

BUFx6f_ASAP7_75t_L g2742 ( 
.A(n_2307),
.Y(n_2742)
);

OAI22xp33_ASAP7_75t_L g2743 ( 
.A1(n_2501),
.A2(n_2163),
.B1(n_2248),
.B2(n_1984),
.Y(n_2743)
);

INVx4_ASAP7_75t_L g2744 ( 
.A(n_2403),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_SL g2745 ( 
.A1(n_2320),
.A2(n_2248),
.B1(n_2132),
.B2(n_1928),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2292),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2495),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2295),
.Y(n_2748)
);

BUFx2_ASAP7_75t_L g2749 ( 
.A(n_2586),
.Y(n_2749)
);

BUFx10_ASAP7_75t_L g2750 ( 
.A(n_2445),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2295),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2297),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2333),
.Y(n_2753)
);

INVx3_ASAP7_75t_L g2754 ( 
.A(n_2586),
.Y(n_2754)
);

BUFx4f_ASAP7_75t_SL g2755 ( 
.A(n_2377),
.Y(n_2755)
);

OAI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2460),
.A2(n_2181),
.B1(n_1984),
.B2(n_2195),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_2398),
.Y(n_2757)
);

BUFx4_ASAP7_75t_R g2758 ( 
.A(n_2303),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2483),
.Y(n_2759)
);

AOI22xp33_ASAP7_75t_SL g2760 ( 
.A1(n_2320),
.A2(n_2132),
.B1(n_1928),
.B2(n_1996),
.Y(n_2760)
);

INVx8_ASAP7_75t_L g2761 ( 
.A(n_2391),
.Y(n_2761)
);

AND2x2_ASAP7_75t_L g2762 ( 
.A(n_2532),
.B(n_1977),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_SL g2763 ( 
.A1(n_2514),
.A2(n_2132),
.B1(n_1928),
.B2(n_1996),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2365),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2484),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2613),
.A2(n_2039),
.B1(n_2068),
.B2(n_2007),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2484),
.Y(n_2767)
);

OAI22xp5_ASAP7_75t_L g2768 ( 
.A1(n_2343),
.A2(n_2435),
.B1(n_2473),
.B2(n_2541),
.Y(n_2768)
);

OAI22xp5_ASAP7_75t_L g2769 ( 
.A1(n_2473),
.A2(n_2187),
.B1(n_1928),
.B2(n_2096),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2297),
.Y(n_2770)
);

CKINVDCx5p33_ASAP7_75t_R g2771 ( 
.A(n_2381),
.Y(n_2771)
);

INVx4_ASAP7_75t_L g2772 ( 
.A(n_2403),
.Y(n_2772)
);

BUFx8_ASAP7_75t_L g2773 ( 
.A(n_2305),
.Y(n_2773)
);

CKINVDCx20_ASAP7_75t_R g2774 ( 
.A(n_2305),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2366),
.Y(n_2775)
);

AOI22xp33_ASAP7_75t_L g2776 ( 
.A1(n_2613),
.A2(n_2007),
.B1(n_2070),
.B2(n_2042),
.Y(n_2776)
);

AOI22xp5_ASAP7_75t_SL g2777 ( 
.A1(n_2489),
.A2(n_1928),
.B1(n_2132),
.B2(n_2096),
.Y(n_2777)
);

AOI22xp33_ASAP7_75t_L g2778 ( 
.A1(n_2464),
.A2(n_2070),
.B1(n_2042),
.B2(n_1937),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2366),
.Y(n_2779)
);

CKINVDCx6p67_ASAP7_75t_R g2780 ( 
.A(n_2327),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2307),
.Y(n_2781)
);

AOI22xp33_ASAP7_75t_L g2782 ( 
.A1(n_2474),
.A2(n_1937),
.B1(n_2143),
.B2(n_2004),
.Y(n_2782)
);

INVx1_ASAP7_75t_SL g2783 ( 
.A(n_2365),
.Y(n_2783)
);

BUFx4f_ASAP7_75t_L g2784 ( 
.A(n_2556),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2499),
.Y(n_2785)
);

OAI22xp5_ASAP7_75t_L g2786 ( 
.A1(n_2541),
.A2(n_2096),
.B1(n_2236),
.B2(n_2165),
.Y(n_2786)
);

AOI22xp33_ASAP7_75t_SL g2787 ( 
.A1(n_2278),
.A2(n_2096),
.B1(n_1982),
.B2(n_2004),
.Y(n_2787)
);

AOI22xp33_ASAP7_75t_L g2788 ( 
.A1(n_2478),
.A2(n_2133),
.B1(n_1982),
.B2(n_2170),
.Y(n_2788)
);

INVx6_ASAP7_75t_L g2789 ( 
.A(n_2398),
.Y(n_2789)
);

AOI22xp33_ASAP7_75t_L g2790 ( 
.A1(n_2478),
.A2(n_2300),
.B1(n_2584),
.B2(n_2282),
.Y(n_2790)
);

AOI22xp5_ASAP7_75t_L g2791 ( 
.A1(n_2309),
.A2(n_2133),
.B1(n_2170),
.B2(n_2168),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2369),
.Y(n_2792)
);

CKINVDCx11_ASAP7_75t_R g2793 ( 
.A(n_2327),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2369),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2374),
.Y(n_2795)
);

INVx1_ASAP7_75t_SL g2796 ( 
.A(n_2429),
.Y(n_2796)
);

AOI22xp33_ASAP7_75t_L g2797 ( 
.A1(n_2422),
.A2(n_2168),
.B1(n_2146),
.B2(n_2160),
.Y(n_2797)
);

BUFx12f_ASAP7_75t_L g2798 ( 
.A(n_2442),
.Y(n_2798)
);

INVx5_ASAP7_75t_L g2799 ( 
.A(n_2472),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2374),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2459),
.A2(n_2487),
.B1(n_2468),
.B2(n_2576),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_SL g2802 ( 
.A1(n_2574),
.A2(n_2477),
.B1(n_2273),
.B2(n_2545),
.Y(n_2802)
);

BUFx3_ASAP7_75t_L g2803 ( 
.A(n_2526),
.Y(n_2803)
);

INVx2_ASAP7_75t_SL g2804 ( 
.A(n_2398),
.Y(n_2804)
);

INVx1_ASAP7_75t_L g2805 ( 
.A(n_2385),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2385),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2499),
.Y(n_2807)
);

BUFx2_ASAP7_75t_L g2808 ( 
.A(n_2586),
.Y(n_2808)
);

AOI22xp33_ASAP7_75t_L g2809 ( 
.A1(n_2468),
.A2(n_2146),
.B1(n_2160),
.B2(n_1963),
.Y(n_2809)
);

INVx3_ASAP7_75t_SL g2810 ( 
.A(n_2442),
.Y(n_2810)
);

INVx2_ASAP7_75t_L g2811 ( 
.A(n_2510),
.Y(n_2811)
);

OAI22x1_ASAP7_75t_L g2812 ( 
.A1(n_2310),
.A2(n_2449),
.B1(n_2269),
.B2(n_2357),
.Y(n_2812)
);

AND2x4_ASAP7_75t_L g2813 ( 
.A(n_2586),
.B(n_2002),
.Y(n_2813)
);

CKINVDCx6p67_ASAP7_75t_R g2814 ( 
.A(n_2398),
.Y(n_2814)
);

OAI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2276),
.A2(n_2593),
.B1(n_2466),
.B2(n_2455),
.Y(n_2815)
);

INVx6_ASAP7_75t_L g2816 ( 
.A(n_2398),
.Y(n_2816)
);

CKINVDCx20_ASAP7_75t_R g2817 ( 
.A(n_2284),
.Y(n_2817)
);

CKINVDCx5p33_ASAP7_75t_R g2818 ( 
.A(n_2486),
.Y(n_2818)
);

INVx2_ASAP7_75t_L g2819 ( 
.A(n_2510),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2390),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2544),
.B(n_1977),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2565),
.A2(n_2593),
.B1(n_2622),
.B2(n_2399),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2390),
.Y(n_2823)
);

AOI22xp33_ASAP7_75t_L g2824 ( 
.A1(n_2468),
.A2(n_1963),
.B1(n_2171),
.B2(n_2172),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2397),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2397),
.Y(n_2826)
);

BUFx2_ASAP7_75t_SL g2827 ( 
.A(n_2398),
.Y(n_2827)
);

CKINVDCx6p67_ASAP7_75t_R g2828 ( 
.A(n_2414),
.Y(n_2828)
);

CKINVDCx11_ASAP7_75t_R g2829 ( 
.A(n_2307),
.Y(n_2829)
);

OAI22xp5_ASAP7_75t_L g2830 ( 
.A1(n_2296),
.A2(n_2096),
.B1(n_2236),
.B2(n_2165),
.Y(n_2830)
);

INVx6_ASAP7_75t_L g2831 ( 
.A(n_2414),
.Y(n_2831)
);

BUFx2_ASAP7_75t_L g2832 ( 
.A(n_2310),
.Y(n_2832)
);

AOI22xp33_ASAP7_75t_L g2833 ( 
.A1(n_2468),
.A2(n_2425),
.B1(n_2439),
.B2(n_2409),
.Y(n_2833)
);

BUFx2_ASAP7_75t_SL g2834 ( 
.A(n_2414),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2406),
.Y(n_2835)
);

BUFx2_ASAP7_75t_L g2836 ( 
.A(n_2588),
.Y(n_2836)
);

CKINVDCx14_ASAP7_75t_R g2837 ( 
.A(n_2371),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2559),
.Y(n_2838)
);

BUFx12f_ASAP7_75t_L g2839 ( 
.A(n_2442),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2406),
.Y(n_2840)
);

BUFx2_ASAP7_75t_L g2841 ( 
.A(n_2588),
.Y(n_2841)
);

INVx1_ASAP7_75t_SL g2842 ( 
.A(n_2429),
.Y(n_2842)
);

INVx6_ASAP7_75t_L g2843 ( 
.A(n_2414),
.Y(n_2843)
);

OAI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2413),
.A2(n_2096),
.B1(n_2236),
.B2(n_2165),
.Y(n_2844)
);

AOI22xp33_ASAP7_75t_L g2845 ( 
.A1(n_2425),
.A2(n_2172),
.B1(n_2171),
.B2(n_2179),
.Y(n_2845)
);

BUFx12f_ASAP7_75t_L g2846 ( 
.A(n_2444),
.Y(n_2846)
);

AND2x2_ASAP7_75t_L g2847 ( 
.A(n_2544),
.B(n_1977),
.Y(n_2847)
);

BUFx6f_ASAP7_75t_L g2848 ( 
.A(n_2307),
.Y(n_2848)
);

BUFx4f_ASAP7_75t_SL g2849 ( 
.A(n_2449),
.Y(n_2849)
);

AOI22xp33_ASAP7_75t_L g2850 ( 
.A1(n_2425),
.A2(n_2178),
.B1(n_2179),
.B2(n_2236),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2559),
.Y(n_2851)
);

AOI22xp33_ASAP7_75t_L g2852 ( 
.A1(n_2425),
.A2(n_2178),
.B1(n_2236),
.B2(n_2165),
.Y(n_2852)
);

AOI22xp33_ASAP7_75t_L g2853 ( 
.A1(n_2439),
.A2(n_2236),
.B1(n_2165),
.B2(n_2237),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2408),
.Y(n_2854)
);

AOI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2439),
.A2(n_2165),
.B1(n_2237),
.B2(n_2002),
.Y(n_2855)
);

OAI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2413),
.A2(n_1977),
.B1(n_2237),
.B2(n_2438),
.Y(n_2856)
);

INVx6_ASAP7_75t_L g2857 ( 
.A(n_2414),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2560),
.Y(n_2858)
);

CKINVDCx6p67_ASAP7_75t_R g2859 ( 
.A(n_2414),
.Y(n_2859)
);

NAND2x1p5_ASAP7_75t_L g2860 ( 
.A(n_2477),
.B(n_1977),
.Y(n_2860)
);

BUFx2_ASAP7_75t_L g2861 ( 
.A(n_2588),
.Y(n_2861)
);

INVx11_ASAP7_75t_L g2862 ( 
.A(n_2391),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_L g2863 ( 
.A1(n_2439),
.A2(n_2237),
.B1(n_2409),
.B2(n_2373),
.Y(n_2863)
);

AOI22xp33_ASAP7_75t_L g2864 ( 
.A1(n_2409),
.A2(n_2237),
.B1(n_2475),
.B2(n_2485),
.Y(n_2864)
);

AOI22xp33_ASAP7_75t_L g2865 ( 
.A1(n_2409),
.A2(n_2237),
.B1(n_2485),
.B2(n_2437),
.Y(n_2865)
);

AOI22xp33_ASAP7_75t_L g2866 ( 
.A1(n_2485),
.A2(n_2592),
.B1(n_2594),
.B2(n_2604),
.Y(n_2866)
);

OAI22xp33_ASAP7_75t_L g2867 ( 
.A1(n_2494),
.A2(n_2485),
.B1(n_2334),
.B2(n_2458),
.Y(n_2867)
);

AOI22xp5_ASAP7_75t_L g2868 ( 
.A1(n_2356),
.A2(n_2340),
.B1(n_2470),
.B2(n_2535),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2408),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2415),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2415),
.Y(n_2871)
);

BUFx3_ASAP7_75t_L g2872 ( 
.A(n_2526),
.Y(n_2872)
);

BUFx12f_ASAP7_75t_L g2873 ( 
.A(n_2444),
.Y(n_2873)
);

BUFx4_ASAP7_75t_SL g2874 ( 
.A(n_2410),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2424),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2424),
.Y(n_2876)
);

AOI22xp33_ASAP7_75t_SL g2877 ( 
.A1(n_2477),
.A2(n_2561),
.B1(n_2550),
.B2(n_2445),
.Y(n_2877)
);

AOI22xp33_ASAP7_75t_SL g2878 ( 
.A1(n_2445),
.A2(n_2519),
.B1(n_2581),
.B2(n_2590),
.Y(n_2878)
);

AOI22xp33_ASAP7_75t_SL g2879 ( 
.A1(n_2590),
.A2(n_2598),
.B1(n_2556),
.B2(n_2579),
.Y(n_2879)
);

BUFx3_ASAP7_75t_L g2880 ( 
.A(n_2595),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2604),
.A2(n_2503),
.B1(n_2308),
.B2(n_2324),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2301),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2301),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2560),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2562),
.Y(n_2885)
);

BUFx2_ASAP7_75t_SL g2886 ( 
.A(n_2511),
.Y(n_2886)
);

AOI22xp33_ASAP7_75t_L g2887 ( 
.A1(n_2604),
.A2(n_2503),
.B1(n_2401),
.B2(n_2417),
.Y(n_2887)
);

BUFx3_ASAP7_75t_L g2888 ( 
.A(n_2595),
.Y(n_2888)
);

BUFx2_ASAP7_75t_SL g2889 ( 
.A(n_2511),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_2428),
.B(n_2509),
.Y(n_2890)
);

INVx2_ASAP7_75t_L g2891 ( 
.A(n_2562),
.Y(n_2891)
);

BUFx3_ASAP7_75t_L g2892 ( 
.A(n_2595),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2571),
.Y(n_2893)
);

OAI22xp33_ASAP7_75t_R g2894 ( 
.A1(n_2452),
.A2(n_2580),
.B1(n_2517),
.B2(n_2589),
.Y(n_2894)
);

BUFx12f_ASAP7_75t_L g2895 ( 
.A(n_2444),
.Y(n_2895)
);

OAI22xp33_ASAP7_75t_L g2896 ( 
.A1(n_2494),
.A2(n_2531),
.B1(n_2556),
.B2(n_2419),
.Y(n_2896)
);

INVx1_ASAP7_75t_L g2897 ( 
.A(n_2323),
.Y(n_2897)
);

INVx6_ASAP7_75t_L g2898 ( 
.A(n_2372),
.Y(n_2898)
);

INVx6_ASAP7_75t_L g2899 ( 
.A(n_2372),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2323),
.Y(n_2900)
);

INVx6_ASAP7_75t_L g2901 ( 
.A(n_2372),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2558),
.B(n_2549),
.Y(n_2902)
);

AOI22xp33_ASAP7_75t_L g2903 ( 
.A1(n_2401),
.A2(n_2417),
.B1(n_2418),
.B2(n_2289),
.Y(n_2903)
);

NAND2x1p5_ASAP7_75t_L g2904 ( 
.A(n_2448),
.B(n_2538),
.Y(n_2904)
);

CKINVDCx5p33_ASAP7_75t_R g2905 ( 
.A(n_2389),
.Y(n_2905)
);

INVx2_ASAP7_75t_L g2906 ( 
.A(n_2571),
.Y(n_2906)
);

INVx2_ASAP7_75t_SL g2907 ( 
.A(n_2605),
.Y(n_2907)
);

INVx2_ASAP7_75t_L g2908 ( 
.A(n_2600),
.Y(n_2908)
);

OAI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2531),
.A2(n_2538),
.B1(n_2448),
.B2(n_2421),
.Y(n_2909)
);

OAI22xp5_ASAP7_75t_L g2910 ( 
.A1(n_2316),
.A2(n_2355),
.B1(n_2426),
.B2(n_2451),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2432),
.A2(n_2420),
.B1(n_2391),
.B2(n_2453),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2345),
.Y(n_2912)
);

CKINVDCx6p67_ASAP7_75t_R g2913 ( 
.A(n_2569),
.Y(n_2913)
);

AOI22xp33_ASAP7_75t_SL g2914 ( 
.A1(n_2590),
.A2(n_2598),
.B1(n_2579),
.B2(n_2286),
.Y(n_2914)
);

BUFx4f_ASAP7_75t_SL g2915 ( 
.A(n_2605),
.Y(n_2915)
);

AOI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2418),
.A2(n_2289),
.B1(n_2476),
.B2(n_2590),
.Y(n_2916)
);

BUFx2_ASAP7_75t_L g2917 ( 
.A(n_2588),
.Y(n_2917)
);

INVx4_ASAP7_75t_L g2918 ( 
.A(n_2315),
.Y(n_2918)
);

OAI22xp33_ASAP7_75t_L g2919 ( 
.A1(n_2448),
.A2(n_2538),
.B1(n_2402),
.B2(n_2307),
.Y(n_2919)
);

INVxp33_ASAP7_75t_L g2920 ( 
.A(n_2371),
.Y(n_2920)
);

AOI211xp5_ASAP7_75t_L g2921 ( 
.A1(n_2620),
.A2(n_2298),
.B(n_2596),
.C(n_2431),
.Y(n_2921)
);

INVx2_ASAP7_75t_L g2922 ( 
.A(n_2600),
.Y(n_2922)
);

BUFx8_ASAP7_75t_L g2923 ( 
.A(n_2402),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2345),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2590),
.A2(n_2286),
.B1(n_2402),
.B2(n_2391),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2585),
.B(n_2540),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2346),
.Y(n_2927)
);

INVx2_ASAP7_75t_R g2928 ( 
.A(n_2443),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2418),
.A2(n_2476),
.B1(n_2595),
.B2(n_2315),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2346),
.Y(n_2930)
);

CKINVDCx6p67_ASAP7_75t_R g2931 ( 
.A(n_2569),
.Y(n_2931)
);

BUFx6f_ASAP7_75t_L g2932 ( 
.A(n_2402),
.Y(n_2932)
);

INVx4_ASAP7_75t_L g2933 ( 
.A(n_2315),
.Y(n_2933)
);

OAI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2440),
.A2(n_2402),
.B1(n_2602),
.B2(n_2271),
.Y(n_2934)
);

BUFx3_ASAP7_75t_L g2935 ( 
.A(n_2595),
.Y(n_2935)
);

CKINVDCx6p67_ASAP7_75t_R g2936 ( 
.A(n_2569),
.Y(n_2936)
);

AND2x4_ASAP7_75t_SL g2937 ( 
.A(n_2286),
.B(n_2271),
.Y(n_2937)
);

BUFx8_ASAP7_75t_L g2938 ( 
.A(n_2391),
.Y(n_2938)
);

AOI22xp33_ASAP7_75t_SL g2939 ( 
.A1(n_2286),
.A2(n_2271),
.B1(n_2317),
.B2(n_2332),
.Y(n_2939)
);

AOI22xp33_ASAP7_75t_L g2940 ( 
.A1(n_2418),
.A2(n_2317),
.B1(n_2332),
.B2(n_2331),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2605),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_SL g2942 ( 
.A1(n_2271),
.A2(n_2317),
.B1(n_2332),
.B2(n_2527),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2517),
.Y(n_2943)
);

INVx8_ASAP7_75t_L g2944 ( 
.A(n_2472),
.Y(n_2944)
);

AOI22xp33_ASAP7_75t_L g2945 ( 
.A1(n_2288),
.A2(n_2277),
.B1(n_2393),
.B2(n_2457),
.Y(n_2945)
);

INVx4_ASAP7_75t_L g2946 ( 
.A(n_2472),
.Y(n_2946)
);

NAND2xp5_ASAP7_75t_L g2947 ( 
.A(n_2591),
.B(n_2597),
.Y(n_2947)
);

AND2x2_ASAP7_75t_L g2948 ( 
.A(n_2359),
.B(n_2368),
.Y(n_2948)
);

INVx4_ASAP7_75t_L g2949 ( 
.A(n_2472),
.Y(n_2949)
);

AOI22xp33_ASAP7_75t_L g2950 ( 
.A1(n_2288),
.A2(n_2393),
.B1(n_2457),
.B2(n_2465),
.Y(n_2950)
);

BUFx3_ASAP7_75t_L g2951 ( 
.A(n_2523),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2557),
.B(n_2582),
.Y(n_2952)
);

OAI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2387),
.A2(n_2527),
.B1(n_2618),
.B2(n_2285),
.Y(n_2953)
);

AOI22xp33_ASAP7_75t_L g2954 ( 
.A1(n_2288),
.A2(n_2465),
.B1(n_2481),
.B2(n_2353),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_L g2955 ( 
.A(n_2362),
.B(n_2546),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2348),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2364),
.B(n_2386),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2610),
.Y(n_2958)
);

AOI22xp33_ASAP7_75t_SL g2959 ( 
.A1(n_2527),
.A2(n_2288),
.B1(n_2358),
.B2(n_2280),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2348),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2481),
.A2(n_2360),
.B1(n_2620),
.B2(n_2388),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2375),
.Y(n_2962)
);

OAI21xp5_ASAP7_75t_SL g2963 ( 
.A1(n_2376),
.A2(n_2358),
.B(n_2530),
.Y(n_2963)
);

INVx6_ASAP7_75t_L g2964 ( 
.A(n_2338),
.Y(n_2964)
);

CKINVDCx5p33_ASAP7_75t_R g2965 ( 
.A(n_2603),
.Y(n_2965)
);

INVx6_ASAP7_75t_L g2966 ( 
.A(n_2338),
.Y(n_2966)
);

BUFx2_ASAP7_75t_SL g2967 ( 
.A(n_2583),
.Y(n_2967)
);

AOI22xp33_ASAP7_75t_L g2968 ( 
.A1(n_2481),
.A2(n_2360),
.B1(n_2379),
.B2(n_2388),
.Y(n_2968)
);

OAI22xp5_ASAP7_75t_SL g2969 ( 
.A1(n_2553),
.A2(n_2358),
.B1(n_2603),
.B2(n_2434),
.Y(n_2969)
);

OAI22xp5_ASAP7_75t_L g2970 ( 
.A1(n_2283),
.A2(n_2342),
.B1(n_2380),
.B2(n_2382),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2375),
.Y(n_2971)
);

BUFx8_ASAP7_75t_SL g2972 ( 
.A(n_2605),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2384),
.Y(n_2973)
);

OA22x2_ASAP7_75t_L g2974 ( 
.A1(n_2283),
.A2(n_2342),
.B1(n_2388),
.B2(n_2379),
.Y(n_2974)
);

CKINVDCx5p33_ASAP7_75t_R g2975 ( 
.A(n_2605),
.Y(n_2975)
);

AOI22xp33_ASAP7_75t_SL g2976 ( 
.A1(n_2280),
.A2(n_2434),
.B1(n_2523),
.B2(n_2447),
.Y(n_2976)
);

CKINVDCx20_ASAP7_75t_R g2977 ( 
.A(n_2359),
.Y(n_2977)
);

AOI22xp33_ASAP7_75t_L g2978 ( 
.A1(n_2360),
.A2(n_2388),
.B1(n_2379),
.B2(n_2363),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2384),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2392),
.Y(n_2980)
);

AOI22xp33_ASAP7_75t_L g2981 ( 
.A1(n_2363),
.A2(n_2379),
.B1(n_2293),
.B2(n_2492),
.Y(n_2981)
);

INVx3_ASAP7_75t_L g2982 ( 
.A(n_2619),
.Y(n_2982)
);

CKINVDCx20_ASAP7_75t_R g2983 ( 
.A(n_2368),
.Y(n_2983)
);

BUFx12f_ASAP7_75t_L g2984 ( 
.A(n_2467),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2610),
.Y(n_2985)
);

BUFx3_ASAP7_75t_L g2986 ( 
.A(n_2523),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2392),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2407),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2395),
.B(n_2471),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2407),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2537),
.Y(n_2991)
);

BUFx3_ASAP7_75t_L g2992 ( 
.A(n_2467),
.Y(n_2992)
);

INVx3_ASAP7_75t_L g2993 ( 
.A(n_2619),
.Y(n_2993)
);

INVxp67_ASAP7_75t_SL g2994 ( 
.A(n_2299),
.Y(n_2994)
);

OAI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_2491),
.A2(n_2352),
.B1(n_2363),
.B2(n_2547),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2537),
.Y(n_2996)
);

OAI31xp33_ASAP7_75t_SL g2997 ( 
.A1(n_2680),
.A2(n_2363),
.A3(n_2616),
.B(n_2370),
.Y(n_2997)
);

OAI22xp5_ASAP7_75t_L g2998 ( 
.A1(n_2822),
.A2(n_2335),
.B1(n_2330),
.B2(n_2536),
.Y(n_2998)
);

BUFx3_ASAP7_75t_L g2999 ( 
.A(n_2695),
.Y(n_2999)
);

AOI21x1_ASAP7_75t_SL g3000 ( 
.A1(n_2691),
.A2(n_2338),
.B(n_2361),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2682),
.B(n_2294),
.Y(n_3001)
);

AOI21xp5_ASAP7_75t_L g3002 ( 
.A1(n_2867),
.A2(n_2488),
.B(n_2525),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2943),
.B(n_2516),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2667),
.Y(n_3004)
);

BUFx6f_ASAP7_75t_L g3005 ( 
.A(n_2701),
.Y(n_3005)
);

AND2x4_ASAP7_75t_L g3006 ( 
.A(n_2937),
.B(n_2619),
.Y(n_3006)
);

O2A1O1Ixp5_ASAP7_75t_L g3007 ( 
.A1(n_2896),
.A2(n_2953),
.B(n_2995),
.C(n_2909),
.Y(n_3007)
);

O2A1O1Ixp33_ASAP7_75t_L g3008 ( 
.A1(n_2921),
.A2(n_2383),
.B(n_2354),
.C(n_2548),
.Y(n_3008)
);

AOI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2921),
.A2(n_2497),
.B(n_2615),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2994),
.B(n_2471),
.Y(n_3010)
);

AOI221xp5_ASAP7_75t_L g3011 ( 
.A1(n_2802),
.A2(n_2480),
.B1(n_2482),
.B2(n_2572),
.C(n_2505),
.Y(n_3011)
);

NOR2xp67_ASAP7_75t_L g3012 ( 
.A(n_2799),
.B(n_2443),
.Y(n_3012)
);

OAI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2822),
.A2(n_2335),
.B1(n_2330),
.B2(n_2572),
.Y(n_3013)
);

OA21x2_ASAP7_75t_L g3014 ( 
.A1(n_2963),
.A2(n_2456),
.B(n_2463),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2682),
.B(n_2294),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_2902),
.B(n_2480),
.Y(n_3016)
);

HB1xp67_ASAP7_75t_L g3017 ( 
.A(n_2753),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2755),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_2667),
.Y(n_3019)
);

AOI21x1_ASAP7_75t_SL g3020 ( 
.A1(n_2762),
.A2(n_2361),
.B(n_2338),
.Y(n_3020)
);

CKINVDCx16_ASAP7_75t_R g3021 ( 
.A(n_2731),
.Y(n_3021)
);

AND2x4_ASAP7_75t_L g3022 ( 
.A(n_2937),
.B(n_2982),
.Y(n_3022)
);

INVx2_ASAP7_75t_L g3023 ( 
.A(n_2667),
.Y(n_3023)
);

OA21x2_ASAP7_75t_L g3024 ( 
.A1(n_2963),
.A2(n_2456),
.B(n_2463),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2749),
.B(n_2294),
.Y(n_3025)
);

OAI22xp5_ASAP7_75t_L g3026 ( 
.A1(n_2868),
.A2(n_2335),
.B1(n_2330),
.B2(n_2528),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2670),
.Y(n_3027)
);

OR2x2_ASAP7_75t_L g3028 ( 
.A(n_2943),
.B(n_2516),
.Y(n_3028)
);

O2A1O1Ixp5_ASAP7_75t_L g3029 ( 
.A1(n_2784),
.A2(n_2302),
.B(n_2555),
.C(n_2567),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_L g3030 ( 
.A(n_2652),
.B(n_2482),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2947),
.B(n_2505),
.Y(n_3031)
);

A2O1A1Ixp33_ASAP7_75t_L g3032 ( 
.A1(n_2868),
.A2(n_2447),
.B(n_2302),
.C(n_2616),
.Y(n_3032)
);

OAI22xp5_ASAP7_75t_L g3033 ( 
.A1(n_2790),
.A2(n_2567),
.B1(n_2555),
.B2(n_2528),
.Y(n_3033)
);

AND2x4_ASAP7_75t_L g3034 ( 
.A(n_2937),
.B(n_2461),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2951),
.Y(n_3035)
);

AOI21xp5_ASAP7_75t_SL g3036 ( 
.A1(n_2768),
.A2(n_2497),
.B(n_2361),
.Y(n_3036)
);

OAI22xp5_ASAP7_75t_L g3037 ( 
.A1(n_2801),
.A2(n_2496),
.B1(n_2361),
.B2(n_2553),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2951),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2670),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2749),
.B(n_2542),
.Y(n_3040)
);

AND2x4_ASAP7_75t_L g3041 ( 
.A(n_2982),
.B(n_2441),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2808),
.B(n_2542),
.Y(n_3042)
);

AOI21xp5_ASAP7_75t_SL g3043 ( 
.A1(n_2769),
.A2(n_2434),
.B(n_2619),
.Y(n_3043)
);

O2A1O1Ixp5_ASAP7_75t_L g3044 ( 
.A1(n_2784),
.A2(n_2351),
.B(n_2349),
.C(n_2344),
.Y(n_3044)
);

AOI21xp5_ASAP7_75t_SL g3045 ( 
.A1(n_2812),
.A2(n_2624),
.B(n_2306),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2670),
.Y(n_3046)
);

AOI21xp5_ASAP7_75t_L g3047 ( 
.A1(n_2881),
.A2(n_2606),
.B(n_2350),
.Y(n_3047)
);

NOR2xp67_ASAP7_75t_L g3048 ( 
.A(n_2799),
.B(n_2623),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_L g3049 ( 
.A(n_2890),
.B(n_2955),
.Y(n_3049)
);

AOI21x1_ASAP7_75t_SL g3050 ( 
.A1(n_2762),
.A2(n_2336),
.B(n_2337),
.Y(n_3050)
);

O2A1O1Ixp33_ASAP7_75t_L g3051 ( 
.A1(n_2815),
.A2(n_2655),
.B(n_2736),
.C(n_2830),
.Y(n_3051)
);

HB1xp67_ASAP7_75t_L g3052 ( 
.A(n_2764),
.Y(n_3052)
);

O2A1O1Ixp5_ASAP7_75t_L g3053 ( 
.A1(n_2784),
.A2(n_2450),
.B(n_2396),
.C(n_2416),
.Y(n_3053)
);

AND2x2_ASAP7_75t_L g3054 ( 
.A(n_2808),
.B(n_2627),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_2991),
.B(n_2518),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2627),
.B(n_2518),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2926),
.B(n_2339),
.Y(n_3057)
);

AND2x4_ASAP7_75t_L g3058 ( 
.A(n_2982),
.B(n_2506),
.Y(n_3058)
);

AND2x4_ASAP7_75t_L g3059 ( 
.A(n_2982),
.B(n_2462),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2649),
.A2(n_2784),
.B(n_2711),
.Y(n_3060)
);

AND2x6_ASAP7_75t_L g3061 ( 
.A(n_2629),
.B(n_2436),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_L g3062 ( 
.A(n_2952),
.B(n_2747),
.Y(n_3062)
);

OAI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2630),
.A2(n_2321),
.B1(n_2311),
.B2(n_2306),
.Y(n_3063)
);

NOR2xp67_ASAP7_75t_L g3064 ( 
.A(n_2799),
.B(n_2621),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2673),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2993),
.B(n_2462),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2673),
.Y(n_3067)
);

AND2x2_ASAP7_75t_L g3068 ( 
.A(n_2696),
.B(n_2370),
.Y(n_3068)
);

AOI21xp5_ASAP7_75t_L g3069 ( 
.A1(n_2649),
.A2(n_2350),
.B(n_2313),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_2696),
.B(n_2436),
.Y(n_3070)
);

NOR2xp67_ASAP7_75t_L g3071 ( 
.A(n_2799),
.B(n_2621),
.Y(n_3071)
);

A2O1A1Ixp33_ASAP7_75t_L g3072 ( 
.A1(n_2777),
.A2(n_2624),
.B(n_2367),
.C(n_2493),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2951),
.Y(n_3073)
);

NOR2xp67_ASAP7_75t_L g3074 ( 
.A(n_2799),
.B(n_2623),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_L g3075 ( 
.A(n_2957),
.B(n_2339),
.Y(n_3075)
);

AOI21xp5_ASAP7_75t_L g3076 ( 
.A1(n_2777),
.A2(n_2350),
.B(n_2313),
.Y(n_3076)
);

O2A1O1Ixp33_ASAP7_75t_L g3077 ( 
.A1(n_2655),
.A2(n_2607),
.B(n_2479),
.C(n_2583),
.Y(n_3077)
);

OAI22xp5_ASAP7_75t_L g3078 ( 
.A1(n_2633),
.A2(n_2321),
.B1(n_2311),
.B2(n_2306),
.Y(n_3078)
);

AOI21xp5_ASAP7_75t_SL g3079 ( 
.A1(n_2812),
.A2(n_2624),
.B(n_2306),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2673),
.Y(n_3080)
);

AOI21xp5_ASAP7_75t_L g3081 ( 
.A1(n_2628),
.A2(n_2350),
.B(n_2313),
.Y(n_3081)
);

AND2x4_ASAP7_75t_L g3082 ( 
.A(n_2993),
.B(n_2479),
.Y(n_3082)
);

O2A1O1Ixp33_ASAP7_75t_L g3083 ( 
.A1(n_2910),
.A2(n_2607),
.B(n_2416),
.C(n_2450),
.Y(n_3083)
);

A2O1A1Ixp33_ASAP7_75t_L g3084 ( 
.A1(n_2877),
.A2(n_2624),
.B(n_2367),
.C(n_2441),
.Y(n_3084)
);

AOI211xp5_ASAP7_75t_L g3085 ( 
.A1(n_2969),
.A2(n_2894),
.B(n_2724),
.C(n_2919),
.Y(n_3085)
);

AOI21x1_ASAP7_75t_SL g3086 ( 
.A1(n_2821),
.A2(n_2321),
.B(n_2293),
.Y(n_3086)
);

O2A1O1Ixp5_ASAP7_75t_L g3087 ( 
.A1(n_2934),
.A2(n_2450),
.B(n_2507),
.C(n_2416),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2849),
.A2(n_2321),
.B1(n_2396),
.B2(n_2507),
.Y(n_3088)
);

OA21x2_ASAP7_75t_L g3089 ( 
.A1(n_2715),
.A2(n_2625),
.B(n_2617),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2989),
.B(n_2905),
.Y(n_3090)
);

OAI22xp5_ASAP7_75t_L g3091 ( 
.A1(n_2645),
.A2(n_2507),
.B1(n_2396),
.B2(n_2520),
.Y(n_3091)
);

AOI21x1_ASAP7_75t_SL g3092 ( 
.A1(n_2821),
.A2(n_2322),
.B(n_2325),
.Y(n_3092)
);

BUFx4f_ASAP7_75t_L g3093 ( 
.A(n_2639),
.Y(n_3093)
);

AND2x2_ASAP7_75t_L g3094 ( 
.A(n_2697),
.B(n_2727),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2700),
.B(n_2818),
.Y(n_3095)
);

NOR2xp33_ASAP7_75t_L g3096 ( 
.A(n_2668),
.B(n_2676),
.Y(n_3096)
);

AOI21xp5_ASAP7_75t_L g3097 ( 
.A1(n_2644),
.A2(n_2350),
.B(n_2318),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2865),
.A2(n_2433),
.B1(n_2506),
.B2(n_2520),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2697),
.B(n_2727),
.Y(n_3099)
);

AOI21xp5_ASAP7_75t_L g3100 ( 
.A1(n_2694),
.A2(n_2607),
.B(n_2522),
.Y(n_3100)
);

CKINVDCx16_ASAP7_75t_R g3101 ( 
.A(n_2731),
.Y(n_3101)
);

HB1xp67_ASAP7_75t_L g3102 ( 
.A(n_2832),
.Y(n_3102)
);

OR2x2_ASAP7_75t_L g3103 ( 
.A(n_2991),
.B(n_2625),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2710),
.Y(n_3104)
);

O2A1O1Ixp5_ASAP7_75t_L g3105 ( 
.A1(n_2946),
.A2(n_2617),
.B(n_2312),
.C(n_2319),
.Y(n_3105)
);

OAI22xp5_ASAP7_75t_L g3106 ( 
.A1(n_2863),
.A2(n_2461),
.B1(n_2493),
.B2(n_2433),
.Y(n_3106)
);

AOI21xp5_ASAP7_75t_L g3107 ( 
.A1(n_2626),
.A2(n_2522),
.B(n_2533),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2710),
.Y(n_3108)
);

AND2x4_ASAP7_75t_L g3109 ( 
.A(n_2993),
.B(n_2410),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2729),
.B(n_2325),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_2993),
.B(n_2500),
.Y(n_3111)
);

INVx1_ASAP7_75t_SL g3112 ( 
.A(n_2688),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2729),
.B(n_2322),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2710),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_2911),
.B(n_2312),
.Y(n_3115)
);

O2A1O1Ixp5_ASAP7_75t_L g3116 ( 
.A1(n_2946),
.A2(n_2319),
.B(n_2423),
.C(n_2612),
.Y(n_3116)
);

OA21x2_ASAP7_75t_L g3117 ( 
.A1(n_2961),
.A2(n_2663),
.B(n_2887),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_2911),
.A2(n_2612),
.B1(n_2508),
.B2(n_2512),
.Y(n_3118)
);

BUFx6f_ASAP7_75t_L g3119 ( 
.A(n_2793),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_2836),
.B(n_2508),
.Y(n_3120)
);

AND2x2_ASAP7_75t_L g3121 ( 
.A(n_2836),
.B(n_2508),
.Y(n_3121)
);

INVxp67_ASAP7_75t_SL g3122 ( 
.A(n_2894),
.Y(n_3122)
);

NAND2xp5_ASAP7_75t_L g3123 ( 
.A(n_2641),
.B(n_2508),
.Y(n_3123)
);

CKINVDCx20_ASAP7_75t_R g3124 ( 
.A(n_2759),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2731),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2841),
.B(n_2508),
.Y(n_3126)
);

AOI21x1_ASAP7_75t_SL g3127 ( 
.A1(n_2847),
.A2(n_2423),
.B(n_2513),
.Y(n_3127)
);

OAI22xp5_ASAP7_75t_L g3128 ( 
.A1(n_2833),
.A2(n_2512),
.B1(n_2513),
.B2(n_2467),
.Y(n_3128)
);

OAI22xp5_ASAP7_75t_SL g3129 ( 
.A1(n_2817),
.A2(n_2512),
.B1(n_2513),
.B2(n_2467),
.Y(n_3129)
);

AOI21x1_ASAP7_75t_L g3130 ( 
.A1(n_2684),
.A2(n_2533),
.B(n_2522),
.Y(n_3130)
);

OAI22xp5_ASAP7_75t_L g3131 ( 
.A1(n_2864),
.A2(n_2512),
.B1(n_2513),
.B2(n_2467),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2631),
.Y(n_3132)
);

INVx1_ASAP7_75t_SL g3133 ( 
.A(n_2639),
.Y(n_3133)
);

NAND2xp5_ASAP7_75t_L g3134 ( 
.A(n_2641),
.B(n_2500),
.Y(n_3134)
);

AOI21x1_ASAP7_75t_SL g3135 ( 
.A1(n_2847),
.A2(n_2500),
.B(n_2512),
.Y(n_3135)
);

CKINVDCx5p33_ASAP7_75t_R g3136 ( 
.A(n_2674),
.Y(n_3136)
);

O2A1O1Ixp5_ASAP7_75t_L g3137 ( 
.A1(n_2946),
.A2(n_2500),
.B(n_2513),
.C(n_2522),
.Y(n_3137)
);

OR2x2_ASAP7_75t_L g3138 ( 
.A(n_2996),
.B(n_2281),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2658),
.B(n_2500),
.Y(n_3139)
);

OR2x2_ASAP7_75t_L g3140 ( 
.A(n_2996),
.B(n_2281),
.Y(n_3140)
);

CKINVDCx5p33_ASAP7_75t_R g3141 ( 
.A(n_2674),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2658),
.B(n_2281),
.Y(n_3142)
);

OAI22xp5_ASAP7_75t_L g3143 ( 
.A1(n_2853),
.A2(n_2533),
.B1(n_2281),
.B2(n_2326),
.Y(n_3143)
);

BUFx12f_ASAP7_75t_L g3144 ( 
.A(n_2638),
.Y(n_3144)
);

OA21x2_ASAP7_75t_L g3145 ( 
.A1(n_2663),
.A2(n_2326),
.B(n_2533),
.Y(n_3145)
);

AND2x2_ASAP7_75t_L g3146 ( 
.A(n_2841),
.B(n_2281),
.Y(n_3146)
);

O2A1O1Ixp5_ASAP7_75t_L g3147 ( 
.A1(n_2946),
.A2(n_2949),
.B(n_2970),
.C(n_2684),
.Y(n_3147)
);

NOR2xp67_ASAP7_75t_L g3148 ( 
.A(n_2799),
.B(n_2949),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_2949),
.B(n_2813),
.Y(n_3149)
);

A2O1A1Ixp33_ASAP7_75t_L g3150 ( 
.A1(n_2878),
.A2(n_2636),
.B(n_2866),
.C(n_2745),
.Y(n_3150)
);

OAI22xp5_ASAP7_75t_L g3151 ( 
.A1(n_2709),
.A2(n_2636),
.B1(n_2639),
.B2(n_2780),
.Y(n_3151)
);

O2A1O1Ixp33_ASAP7_75t_L g3152 ( 
.A1(n_2786),
.A2(n_2844),
.B(n_2719),
.C(n_2856),
.Y(n_3152)
);

AOI21x1_ASAP7_75t_SL g3153 ( 
.A1(n_2813),
.A2(n_2725),
.B(n_2642),
.Y(n_3153)
);

A2O1A1Ixp33_ASAP7_75t_L g3154 ( 
.A1(n_2763),
.A2(n_2981),
.B(n_2954),
.C(n_2787),
.Y(n_3154)
);

CKINVDCx11_ASAP7_75t_R g3155 ( 
.A(n_2638),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2631),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2689),
.B(n_2783),
.Y(n_3157)
);

AND2x2_ASAP7_75t_L g3158 ( 
.A(n_2861),
.B(n_2917),
.Y(n_3158)
);

AOI21xp5_ASAP7_75t_L g3159 ( 
.A1(n_2713),
.A2(n_2635),
.B(n_2687),
.Y(n_3159)
);

AND2x2_ASAP7_75t_L g3160 ( 
.A(n_2861),
.B(n_2917),
.Y(n_3160)
);

NAND2xp5_ASAP7_75t_L g3161 ( 
.A(n_2689),
.B(n_2783),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2796),
.B(n_2842),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2648),
.B(n_2702),
.Y(n_3163)
);

O2A1O1Ixp33_ASAP7_75t_L g3164 ( 
.A1(n_2651),
.A2(n_2756),
.B(n_2860),
.C(n_2743),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2796),
.B(n_2842),
.Y(n_3165)
);

OR2x2_ASAP7_75t_L g3166 ( 
.A(n_2832),
.B(n_2725),
.Y(n_3166)
);

AOI21x1_ASAP7_75t_SL g3167 ( 
.A1(n_2813),
.A2(n_2758),
.B(n_2913),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2940),
.A2(n_2657),
.B(n_2643),
.Y(n_3168)
);

INVx1_ASAP7_75t_L g3169 ( 
.A(n_2637),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_2637),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_2654),
.Y(n_3171)
);

AOI21x1_ASAP7_75t_SL g3172 ( 
.A1(n_2813),
.A2(n_2931),
.B(n_2913),
.Y(n_3172)
);

AND2x4_ASAP7_75t_L g3173 ( 
.A(n_2949),
.B(n_2754),
.Y(n_3173)
);

OR2x2_ASAP7_75t_L g3174 ( 
.A(n_2860),
.B(n_2648),
.Y(n_3174)
);

A2O1A1Ixp33_ASAP7_75t_L g3175 ( 
.A1(n_2760),
.A2(n_2879),
.B(n_2686),
.C(n_2945),
.Y(n_3175)
);

NAND2xp5_ASAP7_75t_L g3176 ( 
.A(n_2948),
.B(n_2903),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2948),
.B(n_2950),
.Y(n_3177)
);

NAND2xp5_ASAP7_75t_L g3178 ( 
.A(n_2920),
.B(n_2916),
.Y(n_3178)
);

AOI21x1_ASAP7_75t_SL g3179 ( 
.A1(n_2931),
.A2(n_2936),
.B(n_2780),
.Y(n_3179)
);

NAND2xp5_ASAP7_75t_L g3180 ( 
.A(n_2882),
.B(n_2883),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2654),
.Y(n_3181)
);

AOI21xp5_ASAP7_75t_L g3182 ( 
.A1(n_2724),
.A2(n_2650),
.B(n_2677),
.Y(n_3182)
);

OAI22xp5_ASAP7_75t_L g3183 ( 
.A1(n_2886),
.A2(n_2889),
.B1(n_2965),
.B2(n_2978),
.Y(n_3183)
);

A2O1A1Ixp33_ASAP7_75t_L g3184 ( 
.A1(n_2976),
.A2(n_2944),
.B(n_2968),
.C(n_2733),
.Y(n_3184)
);

AOI21xp5_ASAP7_75t_L g3185 ( 
.A1(n_2969),
.A2(n_2672),
.B(n_2671),
.Y(n_3185)
);

OA22x2_ASAP7_75t_L g3186 ( 
.A1(n_2771),
.A2(n_2889),
.B1(n_2886),
.B2(n_2662),
.Y(n_3186)
);

AOI21xp5_ASAP7_75t_SL g3187 ( 
.A1(n_2904),
.A2(n_2757),
.B(n_2662),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2653),
.A2(n_2647),
.B(n_2782),
.Y(n_3188)
);

OAI22xp5_ASAP7_75t_L g3189 ( 
.A1(n_2929),
.A2(n_2862),
.B1(n_2852),
.B2(n_2664),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2661),
.Y(n_3190)
);

AOI21xp5_ASAP7_75t_SL g3191 ( 
.A1(n_2904),
.A2(n_2804),
.B(n_2757),
.Y(n_3191)
);

AND2x2_ASAP7_75t_L g3192 ( 
.A(n_2648),
.B(n_2702),
.Y(n_3192)
);

INVx3_ASAP7_75t_L g3193 ( 
.A(n_2634),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2882),
.B(n_2883),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_2661),
.Y(n_3195)
);

AND2x4_ASAP7_75t_L g3196 ( 
.A(n_2754),
.B(n_2648),
.Y(n_3196)
);

OA21x2_ASAP7_75t_L g3197 ( 
.A1(n_2721),
.A2(n_2767),
.B(n_2765),
.Y(n_3197)
);

INVx2_ASAP7_75t_L g3198 ( 
.A(n_2734),
.Y(n_3198)
);

O2A1O1Ixp5_ASAP7_75t_L g3199 ( 
.A1(n_2703),
.A2(n_2772),
.B(n_2744),
.C(n_2918),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2862),
.A2(n_2675),
.B1(n_2674),
.B2(n_2774),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2897),
.B(n_2900),
.Y(n_3201)
);

OA21x2_ASAP7_75t_L g3202 ( 
.A1(n_2765),
.A2(n_2785),
.B(n_2767),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2702),
.B(n_2720),
.Y(n_3203)
);

NOR2xp33_ASAP7_75t_L g3204 ( 
.A(n_2638),
.B(n_2773),
.Y(n_3204)
);

BUFx3_ASAP7_75t_L g3205 ( 
.A(n_2638),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2665),
.Y(n_3206)
);

NAND2xp5_ASAP7_75t_L g3207 ( 
.A(n_2897),
.B(n_2900),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2702),
.B(n_2720),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2720),
.B(n_2754),
.Y(n_3209)
);

O2A1O1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2860),
.A2(n_2810),
.B(n_2904),
.C(n_2804),
.Y(n_3210)
);

OR2x2_ASAP7_75t_L g3211 ( 
.A(n_2720),
.B(n_2754),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2634),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2647),
.A2(n_2944),
.B(n_2693),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_2912),
.B(n_2924),
.Y(n_3214)
);

A2O1A1Ixp33_ASAP7_75t_L g3215 ( 
.A1(n_2944),
.A2(n_2733),
.B(n_2761),
.C(n_2678),
.Y(n_3215)
);

A2O1A1Ixp33_ASAP7_75t_L g3216 ( 
.A1(n_2944),
.A2(n_2761),
.B(n_2678),
.C(n_2722),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_2912),
.B(n_2924),
.Y(n_3217)
);

CKINVDCx16_ASAP7_75t_R g3218 ( 
.A(n_2837),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_2665),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_2927),
.B(n_2930),
.Y(n_3220)
);

O2A1O1Ixp5_ASAP7_75t_L g3221 ( 
.A1(n_2703),
.A2(n_2772),
.B(n_2744),
.C(n_2918),
.Y(n_3221)
);

AOI21xp5_ASAP7_75t_L g3222 ( 
.A1(n_2944),
.A2(n_2740),
.B(n_2660),
.Y(n_3222)
);

OAI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_2914),
.A2(n_2855),
.B1(n_2850),
.B2(n_2707),
.Y(n_3223)
);

O2A1O1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_2810),
.A2(n_2778),
.B(n_2692),
.C(n_2634),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_2927),
.B(n_2930),
.Y(n_3225)
);

AND2x2_ASAP7_75t_L g3226 ( 
.A(n_2974),
.B(n_2986),
.Y(n_3226)
);

OA22x2_ASAP7_75t_L g3227 ( 
.A1(n_2967),
.A2(n_2975),
.B1(n_2834),
.B2(n_2827),
.Y(n_3227)
);

NAND2xp5_ASAP7_75t_L g3228 ( 
.A(n_2956),
.B(n_2960),
.Y(n_3228)
);

INVx1_ASAP7_75t_SL g3229 ( 
.A(n_2874),
.Y(n_3229)
);

O2A1O1Ixp5_ASAP7_75t_L g3230 ( 
.A1(n_2703),
.A2(n_2744),
.B(n_2772),
.C(n_2933),
.Y(n_3230)
);

INVx1_ASAP7_75t_SL g3231 ( 
.A(n_2972),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2974),
.B(n_2986),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2734),
.Y(n_3233)
);

INVx4_ASAP7_75t_SL g3234 ( 
.A(n_2669),
.Y(n_3234)
);

AND2x4_ASAP7_75t_L g3235 ( 
.A(n_2986),
.B(n_2683),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2734),
.Y(n_3236)
);

HB1xp67_ASAP7_75t_L g3237 ( 
.A(n_2679),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_2735),
.Y(n_3238)
);

AND2x2_ASAP7_75t_L g3239 ( 
.A(n_2974),
.B(n_2959),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_2880),
.B(n_2888),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2679),
.Y(n_3241)
);

OR2x2_ASAP7_75t_L g3242 ( 
.A(n_2717),
.B(n_2728),
.Y(n_3242)
);

O2A1O1Ixp5_ASAP7_75t_L g3243 ( 
.A1(n_2703),
.A2(n_2772),
.B(n_2744),
.C(n_2918),
.Y(n_3243)
);

AND2x4_ASAP7_75t_L g3244 ( 
.A(n_2683),
.B(n_2692),
.Y(n_3244)
);

OAI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_2936),
.A2(n_2723),
.B1(n_2925),
.B2(n_2666),
.Y(n_3245)
);

A2O1A1Ixp33_ASAP7_75t_L g3246 ( 
.A1(n_2678),
.A2(n_2722),
.B(n_2761),
.C(n_2685),
.Y(n_3246)
);

AOI21x1_ASAP7_75t_SL g3247 ( 
.A1(n_2773),
.A2(n_2828),
.B(n_2814),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_2773),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2685),
.A2(n_2732),
.B(n_2716),
.Y(n_3249)
);

AOI21x1_ASAP7_75t_SL g3250 ( 
.A1(n_2773),
.A2(n_2828),
.B(n_2814),
.Y(n_3250)
);

HB1xp67_ASAP7_75t_L g3251 ( 
.A(n_2698),
.Y(n_3251)
);

OAI22xp5_ASAP7_75t_L g3252 ( 
.A1(n_2939),
.A2(n_2983),
.B1(n_2977),
.B2(n_2708),
.Y(n_3252)
);

BUFx3_ASAP7_75t_L g3253 ( 
.A(n_2683),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2698),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_2705),
.Y(n_3255)
);

BUFx2_ASAP7_75t_L g3256 ( 
.A(n_2692),
.Y(n_3256)
);

OR2x6_ASAP7_75t_L g3257 ( 
.A(n_2678),
.B(n_2722),
.Y(n_3257)
);

AND2x2_ASAP7_75t_L g3258 ( 
.A(n_2880),
.B(n_2888),
.Y(n_3258)
);

OAI22xp5_ASAP7_75t_L g3259 ( 
.A1(n_2942),
.A2(n_2791),
.B1(n_2789),
.B2(n_2857),
.Y(n_3259)
);

OAI22xp5_ASAP7_75t_L g3260 ( 
.A1(n_2791),
.A2(n_2789),
.B1(n_2712),
.B2(n_2857),
.Y(n_3260)
);

INVxp67_ASAP7_75t_L g3261 ( 
.A(n_2803),
.Y(n_3261)
);

O2A1O1Ixp5_ASAP7_75t_L g3262 ( 
.A1(n_2918),
.A2(n_2933),
.B(n_2705),
.C(n_2806),
.Y(n_3262)
);

AND2x4_ASAP7_75t_L g3263 ( 
.A(n_2803),
.B(n_2872),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2735),
.Y(n_3264)
);

OAI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_2669),
.A2(n_2789),
.B1(n_2712),
.B2(n_2857),
.Y(n_3265)
);

OA21x2_ASAP7_75t_L g3266 ( 
.A1(n_2765),
.A2(n_2851),
.B(n_2838),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_2766),
.A2(n_2776),
.B(n_2722),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2956),
.B(n_2960),
.Y(n_3268)
);

OA21x2_ASAP7_75t_L g3269 ( 
.A1(n_2767),
.A2(n_2891),
.B(n_2885),
.Y(n_3269)
);

INVx2_ASAP7_75t_L g3270 ( 
.A(n_2735),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_2738),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2738),
.Y(n_3272)
);

O2A1O1Ixp5_ASAP7_75t_L g3273 ( 
.A1(n_2933),
.A2(n_2820),
.B(n_2876),
.C(n_2794),
.Y(n_3273)
);

AOI21x1_ASAP7_75t_SL g3274 ( 
.A1(n_2859),
.A2(n_2810),
.B(n_2632),
.Y(n_3274)
);

AND2x2_ASAP7_75t_L g3275 ( 
.A(n_2880),
.B(n_2888),
.Y(n_3275)
);

AND2x2_ASAP7_75t_L g3276 ( 
.A(n_2892),
.B(n_2935),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_2738),
.Y(n_3277)
);

BUFx12f_ASAP7_75t_L g3278 ( 
.A(n_2829),
.Y(n_3278)
);

AND2x2_ASAP7_75t_L g3279 ( 
.A(n_2892),
.B(n_2935),
.Y(n_3279)
);

BUFx12f_ASAP7_75t_L g3280 ( 
.A(n_2798),
.Y(n_3280)
);

O2A1O1Ixp33_ASAP7_75t_L g3281 ( 
.A1(n_2803),
.A2(n_2872),
.B(n_2907),
.C(n_2941),
.Y(n_3281)
);

OR2x2_ASAP7_75t_L g3282 ( 
.A(n_2717),
.B(n_2728),
.Y(n_3282)
);

O2A1O1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_2872),
.A2(n_2941),
.B(n_2907),
.C(n_2935),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_2892),
.B(n_2964),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_2739),
.Y(n_3285)
);

O2A1O1Ixp33_ASAP7_75t_L g3286 ( 
.A1(n_2785),
.A2(n_2807),
.B(n_2891),
.C(n_2885),
.Y(n_3286)
);

INVx2_ASAP7_75t_SL g3287 ( 
.A(n_2964),
.Y(n_3287)
);

AOI21xp5_ASAP7_75t_L g3288 ( 
.A1(n_2678),
.A2(n_2722),
.B(n_2761),
.Y(n_3288)
);

OR2x2_ASAP7_75t_L g3289 ( 
.A(n_2717),
.B(n_2728),
.Y(n_3289)
);

AOI21xp5_ASAP7_75t_SL g3290 ( 
.A1(n_2933),
.A2(n_2629),
.B(n_2681),
.Y(n_3290)
);

HB1xp67_ASAP7_75t_L g3291 ( 
.A(n_2739),
.Y(n_3291)
);

OR2x6_ASAP7_75t_L g3292 ( 
.A(n_2761),
.B(n_2827),
.Y(n_3292)
);

BUFx2_ASAP7_75t_L g3293 ( 
.A(n_2938),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_2797),
.A2(n_2699),
.B(n_2718),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_2739),
.Y(n_3295)
);

BUFx3_ASAP7_75t_L g3296 ( 
.A(n_2992),
.Y(n_3296)
);

OR2x2_ASAP7_75t_L g3297 ( 
.A(n_2893),
.B(n_2906),
.Y(n_3297)
);

OAI22xp5_ASAP7_75t_L g3298 ( 
.A1(n_2669),
.A2(n_2857),
.B1(n_2712),
.B2(n_2789),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_2893),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2714),
.Y(n_3300)
);

OAI22xp5_ASAP7_75t_L g3301 ( 
.A1(n_2669),
.A2(n_2857),
.B1(n_2712),
.B2(n_2789),
.Y(n_3301)
);

OAI22xp5_ASAP7_75t_L g3302 ( 
.A1(n_2669),
.A2(n_2712),
.B1(n_2859),
.B2(n_2964),
.Y(n_3302)
);

OR2x2_ASAP7_75t_L g3303 ( 
.A(n_2893),
.B(n_2906),
.Y(n_3303)
);

OR2x2_ASAP7_75t_L g3304 ( 
.A(n_2906),
.B(n_2908),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2714),
.Y(n_3305)
);

O2A1O1Ixp5_ASAP7_75t_L g3306 ( 
.A1(n_2726),
.A2(n_2820),
.B(n_2823),
.C(n_2825),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_2962),
.B(n_2971),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_2964),
.B(n_2966),
.Y(n_3308)
);

AOI21xp5_ASAP7_75t_L g3309 ( 
.A1(n_2704),
.A2(n_2788),
.B(n_2741),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2962),
.B(n_2971),
.Y(n_3310)
);

AND2x2_ASAP7_75t_L g3311 ( 
.A(n_2966),
.B(n_2992),
.Y(n_3311)
);

BUFx3_ASAP7_75t_L g3312 ( 
.A(n_2992),
.Y(n_3312)
);

HB1xp67_ASAP7_75t_L g3313 ( 
.A(n_2973),
.Y(n_3313)
);

OA21x2_ASAP7_75t_L g3314 ( 
.A1(n_2785),
.A2(n_2838),
.B(n_2891),
.Y(n_3314)
);

AND2x2_ASAP7_75t_L g3315 ( 
.A(n_2966),
.B(n_2908),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_2966),
.B(n_2908),
.Y(n_3316)
);

OAI22xp5_ASAP7_75t_L g3317 ( 
.A1(n_2632),
.A2(n_2690),
.B1(n_2816),
.B2(n_2843),
.Y(n_3317)
);

AOI21xp5_ASAP7_75t_L g3318 ( 
.A1(n_2706),
.A2(n_2809),
.B(n_2824),
.Y(n_3318)
);

AOI21x1_ASAP7_75t_SL g3319 ( 
.A1(n_2632),
.A2(n_2816),
.B(n_2831),
.Y(n_3319)
);

AOI21x1_ASAP7_75t_SL g3320 ( 
.A1(n_2632),
.A2(n_2816),
.B(n_2831),
.Y(n_3320)
);

A2O1A1Ixp33_ASAP7_75t_L g3321 ( 
.A1(n_2834),
.A2(n_2967),
.B(n_2640),
.C(n_2629),
.Y(n_3321)
);

OR2x2_ASAP7_75t_L g3322 ( 
.A(n_2922),
.B(n_2958),
.Y(n_3322)
);

OR2x2_ASAP7_75t_L g3323 ( 
.A(n_2922),
.B(n_2958),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_SL g3324 ( 
.A1(n_2629),
.A2(n_2640),
.B(n_2681),
.Y(n_3324)
);

OAI22xp5_ASAP7_75t_L g3325 ( 
.A1(n_2656),
.A2(n_2816),
.B1(n_2831),
.B2(n_2843),
.Y(n_3325)
);

OAI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_2656),
.A2(n_2831),
.B1(n_2843),
.B2(n_2690),
.Y(n_3326)
);

AND2x2_ASAP7_75t_L g3327 ( 
.A(n_2922),
.B(n_2958),
.Y(n_3327)
);

AND2x4_ASAP7_75t_L g3328 ( 
.A(n_2742),
.B(n_2781),
.Y(n_3328)
);

OAI22xp5_ASAP7_75t_L g3329 ( 
.A1(n_2656),
.A2(n_2843),
.B1(n_2690),
.B2(n_2915),
.Y(n_3329)
);

AOI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_2845),
.A2(n_2629),
.B(n_2640),
.Y(n_3330)
);

AOI21xp5_ASAP7_75t_L g3331 ( 
.A1(n_2629),
.A2(n_2640),
.B(n_2681),
.Y(n_3331)
);

BUFx2_ASAP7_75t_L g3332 ( 
.A(n_2938),
.Y(n_3332)
);

CKINVDCx16_ASAP7_75t_R g3333 ( 
.A(n_2984),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_2985),
.B(n_2973),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2979),
.B(n_2990),
.Y(n_3335)
);

AND2x2_ASAP7_75t_L g3336 ( 
.A(n_2985),
.B(n_2990),
.Y(n_3336)
);

INVx2_ASAP7_75t_L g3337 ( 
.A(n_2985),
.Y(n_3337)
);

OAI22xp5_ASAP7_75t_L g3338 ( 
.A1(n_2656),
.A2(n_2690),
.B1(n_2898),
.B2(n_2899),
.Y(n_3338)
);

HB1xp67_ASAP7_75t_L g3339 ( 
.A(n_2979),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_2980),
.B(n_2988),
.Y(n_3340)
);

OA21x2_ASAP7_75t_L g3341 ( 
.A1(n_2807),
.A2(n_2851),
.B(n_2885),
.Y(n_3341)
);

AOI211xp5_ASAP7_75t_L g3342 ( 
.A1(n_2640),
.A2(n_2681),
.B(n_2932),
.C(n_2781),
.Y(n_3342)
);

AND2x2_ASAP7_75t_L g3343 ( 
.A(n_2980),
.B(n_2988),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2726),
.Y(n_3344)
);

OR2x2_ASAP7_75t_L g3345 ( 
.A(n_2987),
.B(n_2851),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_2987),
.B(n_2928),
.Y(n_3346)
);

BUFx6f_ASAP7_75t_L g3347 ( 
.A(n_2640),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_SL g3348 ( 
.A1(n_2681),
.A2(n_2848),
.B(n_2932),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2737),
.B(n_2825),
.Y(n_3349)
);

AND2x4_ASAP7_75t_SL g3350 ( 
.A(n_2730),
.B(n_2750),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3170),
.Y(n_3351)
);

NAND2xp5_ASAP7_75t_L g3352 ( 
.A(n_3122),
.B(n_2823),
.Y(n_3352)
);

AOI22xp33_ASAP7_75t_L g3353 ( 
.A1(n_3159),
.A2(n_2938),
.B1(n_2839),
.B2(n_2798),
.Y(n_3353)
);

OR2x2_ASAP7_75t_L g3354 ( 
.A(n_3003),
.B(n_2826),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_R g3355 ( 
.A(n_3125),
.B(n_2895),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3219),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3237),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3049),
.B(n_2826),
.Y(n_3358)
);

BUFx2_ASAP7_75t_SL g3359 ( 
.A(n_3005),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_3251),
.Y(n_3360)
);

NOR3xp33_ASAP7_75t_SL g3361 ( 
.A(n_3021),
.B(n_2871),
.C(n_2870),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3132),
.Y(n_3362)
);

AND2x2_ASAP7_75t_L g3363 ( 
.A(n_3239),
.B(n_3226),
.Y(n_3363)
);

INVx2_ASAP7_75t_L g3364 ( 
.A(n_3346),
.Y(n_3364)
);

NAND3xp33_ASAP7_75t_SL g3365 ( 
.A(n_3085),
.B(n_3007),
.C(n_3175),
.Y(n_3365)
);

OR2x2_ASAP7_75t_L g3366 ( 
.A(n_3003),
.B(n_2800),
.Y(n_3366)
);

OR2x2_ASAP7_75t_L g3367 ( 
.A(n_3028),
.B(n_2800),
.Y(n_3367)
);

INVx4_ASAP7_75t_L g3368 ( 
.A(n_3005),
.Y(n_3368)
);

CKINVDCx16_ASAP7_75t_R g3369 ( 
.A(n_3218),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_3132),
.Y(n_3370)
);

CKINVDCx5p33_ASAP7_75t_R g3371 ( 
.A(n_3125),
.Y(n_3371)
);

BUFx3_ASAP7_75t_L g3372 ( 
.A(n_3119),
.Y(n_3372)
);

BUFx2_ASAP7_75t_L g3373 ( 
.A(n_3186),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3150),
.A2(n_2899),
.B1(n_2898),
.B2(n_2901),
.Y(n_3374)
);

AND2x4_ASAP7_75t_L g3375 ( 
.A(n_3234),
.B(n_2681),
.Y(n_3375)
);

BUFx3_ASAP7_75t_L g3376 ( 
.A(n_3119),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_3346),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3239),
.B(n_3226),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_3202),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3102),
.Y(n_3380)
);

AND2x4_ASAP7_75t_L g3381 ( 
.A(n_3234),
.B(n_2781),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_3061),
.Y(n_3382)
);

NAND2xp33_ASAP7_75t_R g3383 ( 
.A(n_3136),
.B(n_2835),
.Y(n_3383)
);

NAND2xp33_ASAP7_75t_R g3384 ( 
.A(n_3136),
.B(n_2835),
.Y(n_3384)
);

INVx3_ASAP7_75t_L g3385 ( 
.A(n_3061),
.Y(n_3385)
);

OR2x2_ASAP7_75t_SL g3386 ( 
.A(n_3218),
.B(n_2901),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_3202),
.Y(n_3387)
);

NAND3xp33_ASAP7_75t_L g3388 ( 
.A(n_3002),
.B(n_2794),
.C(n_2854),
.Y(n_3388)
);

OR2x6_ASAP7_75t_L g3389 ( 
.A(n_3290),
.B(n_2798),
.Y(n_3389)
);

OAI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3154),
.A2(n_2898),
.B1(n_2899),
.B2(n_2901),
.Y(n_3390)
);

OR2x2_ASAP7_75t_L g3391 ( 
.A(n_3028),
.B(n_2795),
.Y(n_3391)
);

INVx3_ASAP7_75t_L g3392 ( 
.A(n_3061),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_3202),
.Y(n_3393)
);

AND2x4_ASAP7_75t_SL g3394 ( 
.A(n_3005),
.B(n_2750),
.Y(n_3394)
);

CKINVDCx5p33_ASAP7_75t_R g3395 ( 
.A(n_3124),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3030),
.B(n_2854),
.Y(n_3396)
);

NOR2x1_ASAP7_75t_L g3397 ( 
.A(n_3290),
.B(n_2795),
.Y(n_3397)
);

CKINVDCx5p33_ASAP7_75t_R g3398 ( 
.A(n_3124),
.Y(n_3398)
);

NOR2xp33_ASAP7_75t_SL g3399 ( 
.A(n_3021),
.B(n_2938),
.Y(n_3399)
);

NOR2xp33_ASAP7_75t_L g3400 ( 
.A(n_3101),
.B(n_3005),
.Y(n_3400)
);

AND2x2_ASAP7_75t_L g3401 ( 
.A(n_3232),
.B(n_2781),
.Y(n_3401)
);

O2A1O1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_3184),
.A2(n_2876),
.B(n_2875),
.C(n_2871),
.Y(n_3402)
);

AND2x2_ASAP7_75t_L g3403 ( 
.A(n_3232),
.B(n_2848),
.Y(n_3403)
);

AOI22xp5_ASAP7_75t_L g3404 ( 
.A1(n_3252),
.A2(n_2839),
.B1(n_2846),
.B2(n_2873),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3156),
.Y(n_3405)
);

INVx2_ASAP7_75t_L g3406 ( 
.A(n_3202),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3156),
.Y(n_3407)
);

AND2x2_ASAP7_75t_SL g3408 ( 
.A(n_2997),
.B(n_2848),
.Y(n_3408)
);

CKINVDCx5p33_ASAP7_75t_R g3409 ( 
.A(n_3101),
.Y(n_3409)
);

AOI22xp33_ASAP7_75t_SL g3410 ( 
.A1(n_3168),
.A2(n_2923),
.B1(n_2899),
.B2(n_2901),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_R g3411 ( 
.A(n_3119),
.B(n_3005),
.Y(n_3411)
);

HB1xp67_ASAP7_75t_L g3412 ( 
.A(n_3017),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3169),
.Y(n_3413)
);

AND2x2_ASAP7_75t_L g3414 ( 
.A(n_3006),
.B(n_2848),
.Y(n_3414)
);

CKINVDCx5p33_ASAP7_75t_R g3415 ( 
.A(n_3119),
.Y(n_3415)
);

CKINVDCx16_ASAP7_75t_R g3416 ( 
.A(n_3278),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_L g3417 ( 
.A(n_3031),
.B(n_2806),
.Y(n_3417)
);

HB1xp67_ASAP7_75t_L g3418 ( 
.A(n_3052),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3016),
.B(n_2752),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_R g3420 ( 
.A(n_3119),
.B(n_2895),
.Y(n_3420)
);

OAI22xp5_ASAP7_75t_L g3421 ( 
.A1(n_3093),
.A2(n_2898),
.B1(n_2932),
.B2(n_2848),
.Y(n_3421)
);

CKINVDCx16_ASAP7_75t_R g3422 ( 
.A(n_3278),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_3033),
.B(n_2805),
.Y(n_3423)
);

AND2x2_ASAP7_75t_L g3424 ( 
.A(n_3006),
.B(n_2781),
.Y(n_3424)
);

BUFx2_ASAP7_75t_L g3425 ( 
.A(n_3186),
.Y(n_3425)
);

NOR3xp33_ASAP7_75t_SL g3426 ( 
.A(n_3141),
.B(n_2775),
.C(n_2869),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3169),
.Y(n_3427)
);

HB1xp67_ASAP7_75t_L g3428 ( 
.A(n_3166),
.Y(n_3428)
);

HB1xp67_ASAP7_75t_L g3429 ( 
.A(n_3166),
.Y(n_3429)
);

NOR3xp33_ASAP7_75t_SL g3430 ( 
.A(n_3141),
.B(n_2775),
.C(n_2840),
.Y(n_3430)
);

CKINVDCx6p67_ASAP7_75t_R g3431 ( 
.A(n_2999),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3171),
.Y(n_3432)
);

INVx2_ASAP7_75t_L g3433 ( 
.A(n_3266),
.Y(n_3433)
);

AO31x2_ASAP7_75t_L g3434 ( 
.A1(n_3072),
.A2(n_3047),
.A3(n_3084),
.B(n_3260),
.Y(n_3434)
);

NAND2xp5_ASAP7_75t_L g3435 ( 
.A(n_3010),
.B(n_2805),
.Y(n_3435)
);

AO31x2_ASAP7_75t_L g3436 ( 
.A1(n_3076),
.A2(n_2819),
.A3(n_2858),
.B(n_2838),
.Y(n_3436)
);

AND2x2_ASAP7_75t_L g3437 ( 
.A(n_3006),
.B(n_2932),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3266),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_L g3439 ( 
.A(n_2999),
.B(n_2873),
.Y(n_3439)
);

BUFx6f_ASAP7_75t_L g3440 ( 
.A(n_3093),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_3115),
.B(n_2792),
.Y(n_3441)
);

OAI22xp5_ASAP7_75t_L g3442 ( 
.A1(n_3093),
.A2(n_2781),
.B1(n_2932),
.B2(n_2848),
.Y(n_3442)
);

OAI21x1_ASAP7_75t_L g3443 ( 
.A1(n_3137),
.A2(n_2811),
.B(n_2858),
.Y(n_3443)
);

INVx6_ASAP7_75t_SL g3444 ( 
.A(n_3257),
.Y(n_3444)
);

INVx1_ASAP7_75t_L g3445 ( 
.A(n_3171),
.Y(n_3445)
);

CKINVDCx16_ASAP7_75t_R g3446 ( 
.A(n_3144),
.Y(n_3446)
);

HB1xp67_ASAP7_75t_L g3447 ( 
.A(n_3313),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3006),
.B(n_2932),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_3062),
.B(n_2792),
.Y(n_3449)
);

AND2x2_ASAP7_75t_L g3450 ( 
.A(n_3054),
.B(n_3158),
.Y(n_3450)
);

CKINVDCx5p33_ASAP7_75t_R g3451 ( 
.A(n_3112),
.Y(n_3451)
);

AND2x4_ASAP7_75t_L g3452 ( 
.A(n_3234),
.B(n_2742),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_R g3453 ( 
.A(n_3155),
.B(n_2895),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3054),
.B(n_2742),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3181),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3158),
.B(n_2742),
.Y(n_3456)
);

OR2x6_ASAP7_75t_L g3457 ( 
.A(n_3043),
.B(n_2846),
.Y(n_3457)
);

AND2x2_ASAP7_75t_L g3458 ( 
.A(n_3160),
.B(n_2742),
.Y(n_3458)
);

NOR2xp33_ASAP7_75t_R g3459 ( 
.A(n_3096),
.B(n_2873),
.Y(n_3459)
);

NOR3xp33_ASAP7_75t_SL g3460 ( 
.A(n_3151),
.B(n_2751),
.C(n_2840),
.Y(n_3460)
);

AOI221xp5_ASAP7_75t_L g3461 ( 
.A1(n_3051),
.A2(n_2770),
.B1(n_2870),
.B2(n_2779),
.C(n_2752),
.Y(n_3461)
);

BUFx3_ASAP7_75t_L g3462 ( 
.A(n_3018),
.Y(n_3462)
);

NAND2xp33_ASAP7_75t_R g3463 ( 
.A(n_3293),
.B(n_2779),
.Y(n_3463)
);

BUFx2_ASAP7_75t_L g3464 ( 
.A(n_3186),
.Y(n_3464)
);

NAND2xp33_ASAP7_75t_R g3465 ( 
.A(n_3293),
.B(n_3332),
.Y(n_3465)
);

BUFx8_ASAP7_75t_SL g3466 ( 
.A(n_3018),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_3057),
.B(n_2751),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3160),
.B(n_2742),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3149),
.B(n_2928),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_3181),
.Y(n_3470)
);

AOI22xp33_ASAP7_75t_SL g3471 ( 
.A1(n_3182),
.A2(n_3223),
.B1(n_3188),
.B2(n_3245),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3190),
.Y(n_3472)
);

AND2x2_ASAP7_75t_L g3473 ( 
.A(n_3149),
.B(n_2750),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3266),
.Y(n_3474)
);

BUFx3_ASAP7_75t_L g3475 ( 
.A(n_3144),
.Y(n_3475)
);

CKINVDCx5p33_ASAP7_75t_R g3476 ( 
.A(n_3229),
.Y(n_3476)
);

AND2x2_ASAP7_75t_L g3477 ( 
.A(n_3149),
.B(n_2750),
.Y(n_3477)
);

AOI22xp33_ASAP7_75t_L g3478 ( 
.A1(n_3185),
.A2(n_2846),
.B1(n_2839),
.B2(n_2923),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3149),
.B(n_2730),
.Y(n_3479)
);

AND2x4_ASAP7_75t_L g3480 ( 
.A(n_3234),
.B(n_2807),
.Y(n_3480)
);

CKINVDCx5p33_ASAP7_75t_R g3481 ( 
.A(n_3280),
.Y(n_3481)
);

INVx3_ASAP7_75t_L g3482 ( 
.A(n_3061),
.Y(n_3482)
);

AO21x2_ASAP7_75t_L g3483 ( 
.A1(n_3107),
.A2(n_2811),
.B(n_2884),
.Y(n_3483)
);

HB1xp67_ASAP7_75t_L g3484 ( 
.A(n_3339),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3094),
.B(n_2730),
.Y(n_3485)
);

NOR3xp33_ASAP7_75t_SL g3486 ( 
.A(n_3204),
.B(n_2746),
.C(n_2748),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3157),
.Y(n_3487)
);

AOI22xp33_ASAP7_75t_L g3488 ( 
.A1(n_3011),
.A2(n_2923),
.B1(n_2646),
.B2(n_2659),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_R g3489 ( 
.A(n_3280),
.B(n_2646),
.Y(n_3489)
);

BUFx2_ASAP7_75t_L g3490 ( 
.A(n_3227),
.Y(n_3490)
);

AND2x4_ASAP7_75t_L g3491 ( 
.A(n_3148),
.B(n_2811),
.Y(n_3491)
);

CKINVDCx16_ASAP7_75t_R g3492 ( 
.A(n_3333),
.Y(n_3492)
);

NAND2xp33_ASAP7_75t_R g3493 ( 
.A(n_3332),
.B(n_2770),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3190),
.Y(n_3494)
);

CKINVDCx5p33_ASAP7_75t_R g3495 ( 
.A(n_3231),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3195),
.Y(n_3496)
);

OR2x6_ASAP7_75t_L g3497 ( 
.A(n_3324),
.B(n_2984),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3195),
.Y(n_3498)
);

AND2x2_ASAP7_75t_L g3499 ( 
.A(n_3094),
.B(n_2730),
.Y(n_3499)
);

OAI22xp5_ASAP7_75t_L g3500 ( 
.A1(n_3060),
.A2(n_2984),
.B1(n_2748),
.B2(n_2746),
.Y(n_3500)
);

OAI22xp5_ASAP7_75t_L g3501 ( 
.A1(n_3133),
.A2(n_2819),
.B1(n_2858),
.B2(n_2884),
.Y(n_3501)
);

AND2x2_ASAP7_75t_L g3502 ( 
.A(n_3099),
.B(n_2819),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3206),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3099),
.B(n_2884),
.Y(n_3504)
);

AND2x4_ASAP7_75t_SL g3505 ( 
.A(n_3257),
.B(n_2646),
.Y(n_3505)
);

CKINVDCx20_ASAP7_75t_R g3506 ( 
.A(n_3248),
.Y(n_3506)
);

NAND2xp5_ASAP7_75t_L g3507 ( 
.A(n_3075),
.B(n_3090),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3037),
.A2(n_2923),
.B1(n_2646),
.B2(n_2659),
.Y(n_3508)
);

AND2x2_ASAP7_75t_L g3509 ( 
.A(n_3022),
.B(n_2659),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3022),
.B(n_2659),
.Y(n_3510)
);

AND2x4_ASAP7_75t_L g3511 ( 
.A(n_3148),
.B(n_3048),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3206),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3241),
.Y(n_3513)
);

OR2x6_ASAP7_75t_L g3514 ( 
.A(n_3043),
.B(n_3187),
.Y(n_3514)
);

AND2x2_ASAP7_75t_L g3515 ( 
.A(n_3022),
.B(n_3308),
.Y(n_3515)
);

INVxp67_ASAP7_75t_SL g3516 ( 
.A(n_3083),
.Y(n_3516)
);

BUFx12f_ASAP7_75t_L g3517 ( 
.A(n_3248),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3200),
.A2(n_3009),
.B1(n_3189),
.B2(n_3318),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3022),
.B(n_3308),
.Y(n_3519)
);

BUFx3_ASAP7_75t_L g3520 ( 
.A(n_3205),
.Y(n_3520)
);

AND2x2_ASAP7_75t_L g3521 ( 
.A(n_3284),
.B(n_3311),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3241),
.Y(n_3522)
);

CKINVDCx5p33_ASAP7_75t_R g3523 ( 
.A(n_3205),
.Y(n_3523)
);

AOI22xp33_ASAP7_75t_L g3524 ( 
.A1(n_3294),
.A2(n_3249),
.B1(n_3117),
.B2(n_3091),
.Y(n_3524)
);

NOR2xp33_ASAP7_75t_R g3525 ( 
.A(n_3333),
.B(n_3095),
.Y(n_3525)
);

NAND3xp33_ASAP7_75t_SL g3526 ( 
.A(n_3164),
.B(n_3147),
.C(n_3152),
.Y(n_3526)
);

OR2x6_ASAP7_75t_L g3527 ( 
.A(n_3187),
.B(n_3191),
.Y(n_3527)
);

CKINVDCx16_ASAP7_75t_R g3528 ( 
.A(n_3129),
.Y(n_3528)
);

CKINVDCx20_ASAP7_75t_R g3529 ( 
.A(n_3183),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3284),
.B(n_3311),
.Y(n_3530)
);

INVx3_ASAP7_75t_L g3531 ( 
.A(n_3061),
.Y(n_3531)
);

BUFx2_ASAP7_75t_L g3532 ( 
.A(n_3227),
.Y(n_3532)
);

OR2x6_ASAP7_75t_L g3533 ( 
.A(n_3191),
.B(n_3036),
.Y(n_3533)
);

CKINVDCx20_ASAP7_75t_R g3534 ( 
.A(n_3257),
.Y(n_3534)
);

OAI22xp5_ASAP7_75t_L g3535 ( 
.A1(n_3032),
.A2(n_3036),
.B1(n_3215),
.B2(n_3246),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_R g3536 ( 
.A(n_3253),
.B(n_3193),
.Y(n_3536)
);

AND2x2_ASAP7_75t_L g3537 ( 
.A(n_3120),
.B(n_3121),
.Y(n_3537)
);

NOR3xp33_ASAP7_75t_SL g3538 ( 
.A(n_3259),
.B(n_3298),
.C(n_3265),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3254),
.Y(n_3539)
);

AND2x2_ASAP7_75t_L g3540 ( 
.A(n_3120),
.B(n_3121),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3254),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3266),
.Y(n_3542)
);

INVx2_ASAP7_75t_L g3543 ( 
.A(n_3269),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3269),
.Y(n_3544)
);

INVx3_ASAP7_75t_L g3545 ( 
.A(n_3061),
.Y(n_3545)
);

OR2x2_ASAP7_75t_L g3546 ( 
.A(n_3055),
.B(n_3142),
.Y(n_3546)
);

CKINVDCx8_ASAP7_75t_R g3547 ( 
.A(n_3347),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3269),
.Y(n_3548)
);

INVx2_ASAP7_75t_SL g3549 ( 
.A(n_3034),
.Y(n_3549)
);

AO31x2_ASAP7_75t_L g3550 ( 
.A1(n_3321),
.A2(n_3100),
.A3(n_3069),
.B(n_3143),
.Y(n_3550)
);

INVx2_ASAP7_75t_L g3551 ( 
.A(n_3269),
.Y(n_3551)
);

BUFx3_ASAP7_75t_L g3552 ( 
.A(n_3253),
.Y(n_3552)
);

BUFx12f_ASAP7_75t_L g3553 ( 
.A(n_3347),
.Y(n_3553)
);

NOR2xp33_ASAP7_75t_R g3554 ( 
.A(n_3193),
.B(n_3212),
.Y(n_3554)
);

NOR2x1_ASAP7_75t_SL g3555 ( 
.A(n_3292),
.B(n_3257),
.Y(n_3555)
);

AND2x2_ASAP7_75t_L g3556 ( 
.A(n_3126),
.B(n_3040),
.Y(n_3556)
);

NAND2xp5_ASAP7_75t_L g3557 ( 
.A(n_3008),
.B(n_3161),
.Y(n_3557)
);

INVx1_ASAP7_75t_SL g3558 ( 
.A(n_3162),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_3255),
.Y(n_3559)
);

OR2x6_ASAP7_75t_L g3560 ( 
.A(n_3045),
.B(n_3079),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_3296),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3255),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3300),
.Y(n_3563)
);

INVx2_ASAP7_75t_L g3564 ( 
.A(n_3314),
.Y(n_3564)
);

AND2x4_ASAP7_75t_L g3565 ( 
.A(n_3048),
.B(n_3064),
.Y(n_3565)
);

OAI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3130),
.A2(n_3227),
.B(n_3319),
.Y(n_3566)
);

HB1xp67_ASAP7_75t_L g3567 ( 
.A(n_3165),
.Y(n_3567)
);

AOI22xp33_ASAP7_75t_L g3568 ( 
.A1(n_3117),
.A2(n_3078),
.B1(n_3222),
.B2(n_3063),
.Y(n_3568)
);

OR2x6_ASAP7_75t_L g3569 ( 
.A(n_3045),
.B(n_3079),
.Y(n_3569)
);

AOI222xp33_ASAP7_75t_L g3570 ( 
.A1(n_3129),
.A2(n_3098),
.B1(n_3106),
.B2(n_2998),
.C1(n_3013),
.C2(n_3118),
.Y(n_3570)
);

HB1xp67_ASAP7_75t_L g3571 ( 
.A(n_3055),
.Y(n_3571)
);

BUFx3_ASAP7_75t_L g3572 ( 
.A(n_3296),
.Y(n_3572)
);

OR2x2_ASAP7_75t_L g3573 ( 
.A(n_3117),
.B(n_3103),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_L g3574 ( 
.A(n_3176),
.B(n_3177),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3097),
.B(n_3178),
.Y(n_3575)
);

CKINVDCx16_ASAP7_75t_R g3576 ( 
.A(n_3292),
.Y(n_3576)
);

AOI22xp33_ASAP7_75t_L g3577 ( 
.A1(n_3117),
.A2(n_3213),
.B1(n_3309),
.B2(n_3026),
.Y(n_3577)
);

A2O1A1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_3224),
.A2(n_3077),
.B(n_3267),
.C(n_3210),
.Y(n_3578)
);

CKINVDCx20_ASAP7_75t_R g3579 ( 
.A(n_3329),
.Y(n_3579)
);

NAND2xp33_ASAP7_75t_SL g3580 ( 
.A(n_3347),
.B(n_3035),
.Y(n_3580)
);

NAND2xp33_ASAP7_75t_R g3581 ( 
.A(n_3256),
.B(n_3035),
.Y(n_3581)
);

NAND2xp33_ASAP7_75t_R g3582 ( 
.A(n_3256),
.B(n_3073),
.Y(n_3582)
);

INVx2_ASAP7_75t_L g3583 ( 
.A(n_3314),
.Y(n_3583)
);

INVx2_ASAP7_75t_L g3584 ( 
.A(n_3314),
.Y(n_3584)
);

AO31x2_ASAP7_75t_L g3585 ( 
.A1(n_3301),
.A2(n_3081),
.A3(n_3317),
.B(n_3325),
.Y(n_3585)
);

HB1xp67_ASAP7_75t_L g3586 ( 
.A(n_3340),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3110),
.B(n_3113),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3314),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_3300),
.Y(n_3589)
);

OAI21x1_ASAP7_75t_L g3590 ( 
.A1(n_3130),
.A2(n_3320),
.B(n_3262),
.Y(n_3590)
);

AO31x2_ASAP7_75t_L g3591 ( 
.A1(n_3326),
.A2(n_3338),
.A3(n_3302),
.B(n_3330),
.Y(n_3591)
);

AO31x2_ASAP7_75t_L g3592 ( 
.A1(n_3131),
.A2(n_3331),
.A3(n_3073),
.B(n_3128),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_R g3593 ( 
.A(n_3193),
.B(n_3212),
.Y(n_3593)
);

CKINVDCx16_ASAP7_75t_R g3594 ( 
.A(n_3292),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3305),
.Y(n_3595)
);

OAI22xp5_ASAP7_75t_L g3596 ( 
.A1(n_3216),
.A2(n_3261),
.B1(n_3342),
.B2(n_3287),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3126),
.B(n_3040),
.Y(n_3597)
);

INVx1_ASAP7_75t_L g3598 ( 
.A(n_3305),
.Y(n_3598)
);

CKINVDCx20_ASAP7_75t_R g3599 ( 
.A(n_3088),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3110),
.B(n_3113),
.Y(n_3600)
);

NOR2x1_ASAP7_75t_SL g3601 ( 
.A(n_3292),
.B(n_3038),
.Y(n_3601)
);

CKINVDCx5p33_ASAP7_75t_R g3602 ( 
.A(n_3312),
.Y(n_3602)
);

HB1xp67_ASAP7_75t_L g3603 ( 
.A(n_3340),
.Y(n_3603)
);

NOR2x1p5_ASAP7_75t_L g3604 ( 
.A(n_3212),
.B(n_3174),
.Y(n_3604)
);

INVx1_ASAP7_75t_L g3605 ( 
.A(n_3344),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_L g3606 ( 
.A(n_3068),
.B(n_3070),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3068),
.B(n_3070),
.Y(n_3607)
);

AND2x2_ASAP7_75t_L g3608 ( 
.A(n_3042),
.B(n_3244),
.Y(n_3608)
);

OR2x2_ASAP7_75t_L g3609 ( 
.A(n_3103),
.B(n_3174),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3315),
.B(n_3316),
.Y(n_3610)
);

NAND2xp33_ASAP7_75t_R g3611 ( 
.A(n_3244),
.B(n_3263),
.Y(n_3611)
);

CKINVDCx5p33_ASAP7_75t_R g3612 ( 
.A(n_3312),
.Y(n_3612)
);

INVx5_ASAP7_75t_L g3613 ( 
.A(n_3061),
.Y(n_3613)
);

HB1xp67_ASAP7_75t_L g3614 ( 
.A(n_3343),
.Y(n_3614)
);

NOR2xp33_ASAP7_75t_R g3615 ( 
.A(n_3179),
.B(n_3287),
.Y(n_3615)
);

NAND2xp33_ASAP7_75t_R g3616 ( 
.A(n_3244),
.B(n_3263),
.Y(n_3616)
);

BUFx3_ASAP7_75t_L g3617 ( 
.A(n_3244),
.Y(n_3617)
);

INVx5_ASAP7_75t_L g3618 ( 
.A(n_3347),
.Y(n_3618)
);

AND2x2_ASAP7_75t_L g3619 ( 
.A(n_3042),
.B(n_3263),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_R g3620 ( 
.A(n_3347),
.B(n_3038),
.Y(n_3620)
);

OA21x2_ASAP7_75t_L g3621 ( 
.A1(n_3116),
.A2(n_3087),
.B(n_3273),
.Y(n_3621)
);

AND2x2_ASAP7_75t_L g3622 ( 
.A(n_3263),
.B(n_3056),
.Y(n_3622)
);

NAND2xp33_ASAP7_75t_R g3623 ( 
.A(n_3235),
.B(n_3328),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3056),
.B(n_3315),
.Y(n_3624)
);

NOR2x1p5_ASAP7_75t_L g3625 ( 
.A(n_3173),
.B(n_3211),
.Y(n_3625)
);

OR2x2_ASAP7_75t_L g3626 ( 
.A(n_3138),
.B(n_3140),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_L g3627 ( 
.A(n_3316),
.B(n_3001),
.Y(n_3627)
);

INVx3_ASAP7_75t_L g3628 ( 
.A(n_3196),
.Y(n_3628)
);

BUFx2_ASAP7_75t_L g3629 ( 
.A(n_3235),
.Y(n_3629)
);

AND2x2_ASAP7_75t_L g3630 ( 
.A(n_3235),
.B(n_3025),
.Y(n_3630)
);

INVx2_ASAP7_75t_L g3631 ( 
.A(n_3341),
.Y(n_3631)
);

NOR2xp33_ASAP7_75t_R g3632 ( 
.A(n_3240),
.B(n_3258),
.Y(n_3632)
);

NOR2x1_ASAP7_75t_SL g3633 ( 
.A(n_3211),
.B(n_3146),
.Y(n_3633)
);

AND2x2_ASAP7_75t_L g3634 ( 
.A(n_3235),
.B(n_3025),
.Y(n_3634)
);

INVx2_ASAP7_75t_L g3635 ( 
.A(n_3341),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3344),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3343),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_L g3638 ( 
.A1(n_3288),
.A2(n_3173),
.B1(n_3058),
.B2(n_3109),
.Y(n_3638)
);

AND2x2_ASAP7_75t_L g3639 ( 
.A(n_3173),
.B(n_3196),
.Y(n_3639)
);

HB1xp67_ASAP7_75t_L g3640 ( 
.A(n_3334),
.Y(n_3640)
);

NAND2xp33_ASAP7_75t_R g3641 ( 
.A(n_3328),
.B(n_3240),
.Y(n_3641)
);

HB1xp67_ASAP7_75t_L g3642 ( 
.A(n_3334),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3306),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3019),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3258),
.B(n_3275),
.Y(n_3645)
);

CKINVDCx16_ASAP7_75t_R g3646 ( 
.A(n_3034),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3341),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3196),
.B(n_3041),
.Y(n_3648)
);

INVx1_ASAP7_75t_L g3649 ( 
.A(n_3019),
.Y(n_3649)
);

AND2x2_ASAP7_75t_L g3650 ( 
.A(n_3196),
.B(n_3041),
.Y(n_3650)
);

AND2x2_ASAP7_75t_L g3651 ( 
.A(n_3041),
.B(n_3058),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3001),
.B(n_3015),
.Y(n_3652)
);

INVx2_ASAP7_75t_L g3653 ( 
.A(n_3341),
.Y(n_3653)
);

INVxp67_ASAP7_75t_SL g3654 ( 
.A(n_3281),
.Y(n_3654)
);

AO31x2_ASAP7_75t_L g3655 ( 
.A1(n_3027),
.A2(n_3080),
.A3(n_3067),
.B(n_3065),
.Y(n_3655)
);

INVx3_ASAP7_75t_L g3656 ( 
.A(n_3111),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3015),
.B(n_3349),
.Y(n_3657)
);

AND2x4_ASAP7_75t_L g3658 ( 
.A(n_3064),
.B(n_3071),
.Y(n_3658)
);

NAND2xp33_ASAP7_75t_SL g3659 ( 
.A(n_3167),
.B(n_3153),
.Y(n_3659)
);

AOI22xp33_ASAP7_75t_L g3660 ( 
.A1(n_3058),
.A2(n_3109),
.B1(n_3279),
.B2(n_3275),
.Y(n_3660)
);

CKINVDCx11_ASAP7_75t_R g3661 ( 
.A(n_3034),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3027),
.Y(n_3662)
);

OR2x2_ASAP7_75t_L g3663 ( 
.A(n_3138),
.B(n_3140),
.Y(n_3663)
);

AOI22xp33_ASAP7_75t_L g3664 ( 
.A1(n_3109),
.A2(n_3279),
.B1(n_3276),
.B2(n_3328),
.Y(n_3664)
);

OR2x2_ASAP7_75t_L g3665 ( 
.A(n_3297),
.B(n_3303),
.Y(n_3665)
);

CKINVDCx9p33_ASAP7_75t_R g3666 ( 
.A(n_3172),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3197),
.Y(n_3667)
);

BUFx6f_ASAP7_75t_L g3668 ( 
.A(n_3372),
.Y(n_3668)
);

BUFx2_ASAP7_75t_L g3669 ( 
.A(n_3444),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3379),
.Y(n_3670)
);

AOI21xp5_ASAP7_75t_SL g3671 ( 
.A1(n_3365),
.A2(n_3283),
.B(n_3024),
.Y(n_3671)
);

OR2x2_ASAP7_75t_L g3672 ( 
.A(n_3643),
.B(n_3180),
.Y(n_3672)
);

AO21x2_ASAP7_75t_L g3673 ( 
.A1(n_3526),
.A2(n_3324),
.B(n_3348),
.Y(n_3673)
);

OR2x2_ASAP7_75t_L g3674 ( 
.A(n_3643),
.B(n_3194),
.Y(n_3674)
);

OA21x2_ASAP7_75t_L g3675 ( 
.A1(n_3590),
.A2(n_3012),
.B(n_3221),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3557),
.B(n_3146),
.Y(n_3676)
);

AO21x2_ASAP7_75t_L g3677 ( 
.A1(n_3578),
.A2(n_3348),
.B(n_3012),
.Y(n_3677)
);

NAND3xp33_ASAP7_75t_L g3678 ( 
.A(n_3471),
.B(n_3024),
.C(n_3014),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3362),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3362),
.Y(n_3680)
);

OA21x2_ASAP7_75t_L g3681 ( 
.A1(n_3590),
.A2(n_3243),
.B(n_3199),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3370),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3370),
.Y(n_3683)
);

AND2x4_ASAP7_75t_L g3684 ( 
.A(n_3613),
.B(n_3071),
.Y(n_3684)
);

AND2x4_ASAP7_75t_L g3685 ( 
.A(n_3613),
.B(n_3074),
.Y(n_3685)
);

OA21x2_ASAP7_75t_L g3686 ( 
.A1(n_3566),
.A2(n_3230),
.B(n_3053),
.Y(n_3686)
);

OA21x2_ASAP7_75t_L g3687 ( 
.A1(n_3566),
.A2(n_3029),
.B(n_3074),
.Y(n_3687)
);

OAI21x1_ASAP7_75t_L g3688 ( 
.A1(n_3397),
.A2(n_3286),
.B(n_3274),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3379),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3387),
.Y(n_3690)
);

OA21x2_ASAP7_75t_L g3691 ( 
.A1(n_3524),
.A2(n_3105),
.B(n_3044),
.Y(n_3691)
);

INVx1_ASAP7_75t_L g3692 ( 
.A(n_3405),
.Y(n_3692)
);

HB1xp67_ASAP7_75t_L g3693 ( 
.A(n_3412),
.Y(n_3693)
);

BUFx3_ASAP7_75t_L g3694 ( 
.A(n_3372),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3405),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3387),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3407),
.Y(n_3697)
);

OAI222xp33_ASAP7_75t_L g3698 ( 
.A1(n_3518),
.A2(n_3139),
.B1(n_3123),
.B2(n_3134),
.C1(n_3276),
.C2(n_3209),
.Y(n_3698)
);

INVx2_ASAP7_75t_L g3699 ( 
.A(n_3393),
.Y(n_3699)
);

BUFx2_ASAP7_75t_L g3700 ( 
.A(n_3444),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3402),
.A2(n_3024),
.B(n_3014),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3393),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3407),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3413),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3406),
.Y(n_3705)
);

OA21x2_ASAP7_75t_L g3706 ( 
.A1(n_3577),
.A2(n_3271),
.B(n_3277),
.Y(n_3706)
);

INVx1_ASAP7_75t_L g3707 ( 
.A(n_3413),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3406),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3433),
.Y(n_3709)
);

AND2x2_ASAP7_75t_L g3710 ( 
.A(n_3490),
.B(n_3209),
.Y(n_3710)
);

NOR2xp33_ASAP7_75t_L g3711 ( 
.A(n_3416),
.B(n_3328),
.Y(n_3711)
);

AND2x4_ASAP7_75t_L g3712 ( 
.A(n_3613),
.B(n_3163),
.Y(n_3712)
);

BUFx2_ASAP7_75t_L g3713 ( 
.A(n_3444),
.Y(n_3713)
);

INVx2_ASAP7_75t_L g3714 ( 
.A(n_3433),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3490),
.B(n_3163),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_3390),
.A2(n_3024),
.B(n_3014),
.Y(n_3716)
);

AO21x2_ASAP7_75t_L g3717 ( 
.A1(n_3667),
.A2(n_3104),
.B(n_3065),
.Y(n_3717)
);

AND2x4_ASAP7_75t_L g3718 ( 
.A(n_3613),
.B(n_3192),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3427),
.Y(n_3719)
);

OR2x6_ASAP7_75t_L g3720 ( 
.A(n_3533),
.B(n_3560),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3427),
.Y(n_3721)
);

OR2x2_ASAP7_75t_L g3722 ( 
.A(n_3352),
.B(n_3201),
.Y(n_3722)
);

AND2x4_ASAP7_75t_L g3723 ( 
.A(n_3613),
.B(n_3192),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3438),
.Y(n_3724)
);

BUFx2_ASAP7_75t_L g3725 ( 
.A(n_3444),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3432),
.Y(n_3726)
);

BUFx2_ASAP7_75t_L g3727 ( 
.A(n_3386),
.Y(n_3727)
);

AO21x2_ASAP7_75t_L g3728 ( 
.A1(n_3667),
.A2(n_3104),
.B(n_3080),
.Y(n_3728)
);

AO21x2_ASAP7_75t_L g3729 ( 
.A1(n_3601),
.A2(n_3067),
.B(n_3039),
.Y(n_3729)
);

CKINVDCx20_ASAP7_75t_R g3730 ( 
.A(n_3395),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3532),
.B(n_3208),
.Y(n_3731)
);

BUFx3_ASAP7_75t_L g3732 ( 
.A(n_3376),
.Y(n_3732)
);

AOI22xp5_ASAP7_75t_L g3733 ( 
.A1(n_3374),
.A2(n_3014),
.B1(n_3350),
.B2(n_3111),
.Y(n_3733)
);

AOI22xp5_ASAP7_75t_L g3734 ( 
.A1(n_3529),
.A2(n_3350),
.B1(n_3111),
.B2(n_3089),
.Y(n_3734)
);

OA21x2_ASAP7_75t_L g3735 ( 
.A1(n_3443),
.A2(n_3271),
.B(n_3277),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3432),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3461),
.B(n_3336),
.Y(n_3737)
);

INVx2_ASAP7_75t_L g3738 ( 
.A(n_3438),
.Y(n_3738)
);

INVx2_ASAP7_75t_L g3739 ( 
.A(n_3474),
.Y(n_3739)
);

INVx1_ASAP7_75t_L g3740 ( 
.A(n_3445),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3575),
.B(n_3336),
.Y(n_3741)
);

OA21x2_ASAP7_75t_L g3742 ( 
.A1(n_3443),
.A2(n_3285),
.B(n_3039),
.Y(n_3742)
);

OR2x2_ASAP7_75t_L g3743 ( 
.A(n_3571),
.B(n_3228),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3532),
.B(n_3208),
.Y(n_3744)
);

AND2x2_ASAP7_75t_L g3745 ( 
.A(n_3555),
.B(n_3203),
.Y(n_3745)
);

INVx2_ASAP7_75t_SL g3746 ( 
.A(n_3376),
.Y(n_3746)
);

AO21x2_ASAP7_75t_L g3747 ( 
.A1(n_3601),
.A2(n_3633),
.B(n_3483),
.Y(n_3747)
);

AND2x2_ASAP7_75t_L g3748 ( 
.A(n_3555),
.B(n_3203),
.Y(n_3748)
);

HB1xp67_ASAP7_75t_L g3749 ( 
.A(n_3418),
.Y(n_3749)
);

AO21x2_ASAP7_75t_L g3750 ( 
.A1(n_3633),
.A2(n_3285),
.B(n_3217),
.Y(n_3750)
);

AND2x2_ASAP7_75t_L g3751 ( 
.A(n_3373),
.B(n_3111),
.Y(n_3751)
);

INVx1_ASAP7_75t_L g3752 ( 
.A(n_3445),
.Y(n_3752)
);

BUFx6f_ASAP7_75t_SL g3753 ( 
.A(n_3368),
.Y(n_3753)
);

AND4x1_ASAP7_75t_L g3754 ( 
.A(n_3400),
.B(n_3247),
.C(n_3250),
.D(n_3127),
.Y(n_3754)
);

AOI22xp5_ASAP7_75t_L g3755 ( 
.A1(n_3369),
.A2(n_3359),
.B1(n_3404),
.B2(n_3388),
.Y(n_3755)
);

OR2x2_ASAP7_75t_L g3756 ( 
.A(n_3428),
.B(n_3207),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3373),
.B(n_3082),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3429),
.B(n_3307),
.Y(n_3758)
);

AND2x2_ASAP7_75t_L g3759 ( 
.A(n_3425),
.B(n_3082),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_3455),
.Y(n_3760)
);

INVx1_ASAP7_75t_L g3761 ( 
.A(n_3455),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3470),
.Y(n_3762)
);

AND2x2_ASAP7_75t_L g3763 ( 
.A(n_3425),
.B(n_3082),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3470),
.Y(n_3764)
);

HB1xp67_ASAP7_75t_L g3765 ( 
.A(n_3380),
.Y(n_3765)
);

AND2x2_ASAP7_75t_L g3766 ( 
.A(n_3464),
.B(n_3533),
.Y(n_3766)
);

BUFx6f_ASAP7_75t_L g3767 ( 
.A(n_3440),
.Y(n_3767)
);

AOI221xp5_ASAP7_75t_L g3768 ( 
.A1(n_3568),
.A2(n_3225),
.B1(n_3214),
.B2(n_3310),
.C(n_3220),
.Y(n_3768)
);

AO21x2_ASAP7_75t_L g3769 ( 
.A1(n_3483),
.A2(n_3268),
.B(n_3335),
.Y(n_3769)
);

NOR2xp33_ASAP7_75t_L g3770 ( 
.A(n_3416),
.B(n_3066),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3472),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3464),
.B(n_3082),
.Y(n_3772)
);

INVx2_ASAP7_75t_L g3773 ( 
.A(n_3474),
.Y(n_3773)
);

AOI22xp33_ASAP7_75t_L g3774 ( 
.A1(n_3659),
.A2(n_3066),
.B1(n_3059),
.B2(n_3089),
.Y(n_3774)
);

AND2x4_ASAP7_75t_L g3775 ( 
.A(n_3613),
.B(n_3066),
.Y(n_3775)
);

INVx2_ASAP7_75t_L g3776 ( 
.A(n_3542),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3472),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3542),
.Y(n_3778)
);

BUFx3_ASAP7_75t_L g3779 ( 
.A(n_3466),
.Y(n_3779)
);

OAI221xp5_ASAP7_75t_L g3780 ( 
.A1(n_3538),
.A2(n_3345),
.B1(n_3291),
.B2(n_3323),
.C(n_3322),
.Y(n_3780)
);

AOI322xp5_ASAP7_75t_L g3781 ( 
.A1(n_3528),
.A2(n_3092),
.A3(n_3004),
.B1(n_3023),
.B2(n_3046),
.C1(n_3108),
.C2(n_3114),
.Y(n_3781)
);

OR2x6_ASAP7_75t_L g3782 ( 
.A(n_3533),
.B(n_3145),
.Y(n_3782)
);

INVx2_ASAP7_75t_L g3783 ( 
.A(n_3543),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3543),
.Y(n_3784)
);

BUFx6f_ASAP7_75t_L g3785 ( 
.A(n_3440),
.Y(n_3785)
);

BUFx4f_ASAP7_75t_SL g3786 ( 
.A(n_3431),
.Y(n_3786)
);

NOR2xp33_ASAP7_75t_L g3787 ( 
.A(n_3422),
.B(n_3066),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3494),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3544),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3494),
.Y(n_3790)
);

OA21x2_ASAP7_75t_L g3791 ( 
.A1(n_3544),
.A2(n_3238),
.B(n_3198),
.Y(n_3791)
);

HB1xp67_ASAP7_75t_L g3792 ( 
.A(n_3447),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3496),
.Y(n_3793)
);

INVxp67_ASAP7_75t_L g3794 ( 
.A(n_3359),
.Y(n_3794)
);

INVxp67_ASAP7_75t_SL g3795 ( 
.A(n_3463),
.Y(n_3795)
);

AOI21x1_ASAP7_75t_L g3796 ( 
.A1(n_3527),
.A2(n_3299),
.B(n_3337),
.Y(n_3796)
);

HB1xp67_ASAP7_75t_L g3797 ( 
.A(n_3484),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3496),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3498),
.Y(n_3799)
);

AOI322xp5_ASAP7_75t_L g3800 ( 
.A1(n_3528),
.A2(n_3114),
.A3(n_3004),
.B1(n_3108),
.B2(n_3023),
.C1(n_3046),
.C2(n_3050),
.Y(n_3800)
);

AOI21xp5_ASAP7_75t_L g3801 ( 
.A1(n_3535),
.A2(n_3059),
.B(n_3197),
.Y(n_3801)
);

BUFx2_ASAP7_75t_L g3802 ( 
.A(n_3386),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3548),
.Y(n_3803)
);

AND2x4_ASAP7_75t_L g3804 ( 
.A(n_3625),
.B(n_3059),
.Y(n_3804)
);

INVxp67_ASAP7_75t_L g3805 ( 
.A(n_3465),
.Y(n_3805)
);

AND2x2_ASAP7_75t_L g3806 ( 
.A(n_3533),
.B(n_3059),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3397),
.A2(n_3135),
.B(n_3000),
.Y(n_3807)
);

INVx1_ASAP7_75t_L g3808 ( 
.A(n_3498),
.Y(n_3808)
);

OR2x2_ASAP7_75t_L g3809 ( 
.A(n_3573),
.B(n_3303),
.Y(n_3809)
);

INVx2_ASAP7_75t_L g3810 ( 
.A(n_3548),
.Y(n_3810)
);

OA21x2_ASAP7_75t_L g3811 ( 
.A1(n_3551),
.A2(n_3272),
.B(n_3264),
.Y(n_3811)
);

OAI221xp5_ASAP7_75t_L g3812 ( 
.A1(n_3478),
.A2(n_3345),
.B1(n_3323),
.B2(n_3322),
.C(n_3304),
.Y(n_3812)
);

INVxp67_ASAP7_75t_L g3813 ( 
.A(n_3654),
.Y(n_3813)
);

OR2x2_ASAP7_75t_L g3814 ( 
.A(n_3573),
.B(n_3304),
.Y(n_3814)
);

OA21x2_ASAP7_75t_L g3815 ( 
.A1(n_3551),
.A2(n_3264),
.B(n_3295),
.Y(n_3815)
);

INVx2_ASAP7_75t_L g3816 ( 
.A(n_3564),
.Y(n_3816)
);

BUFx3_ASAP7_75t_L g3817 ( 
.A(n_3431),
.Y(n_3817)
);

AOI22xp33_ASAP7_75t_L g3818 ( 
.A1(n_3408),
.A2(n_3089),
.B1(n_3197),
.B2(n_3337),
.Y(n_3818)
);

OR2x2_ASAP7_75t_L g3819 ( 
.A(n_3423),
.B(n_3297),
.Y(n_3819)
);

AND2x2_ASAP7_75t_L g3820 ( 
.A(n_3533),
.B(n_3327),
.Y(n_3820)
);

AOI21xp5_ASAP7_75t_SL g3821 ( 
.A1(n_3560),
.A2(n_3145),
.B(n_3197),
.Y(n_3821)
);

INVx1_ASAP7_75t_L g3822 ( 
.A(n_3503),
.Y(n_3822)
);

INVx3_ASAP7_75t_L g3823 ( 
.A(n_3382),
.Y(n_3823)
);

INVx2_ASAP7_75t_L g3824 ( 
.A(n_3564),
.Y(n_3824)
);

OA21x2_ASAP7_75t_L g3825 ( 
.A1(n_3583),
.A2(n_3233),
.B(n_3270),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_3583),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3584),
.Y(n_3827)
);

AO21x1_ASAP7_75t_SL g3828 ( 
.A1(n_3353),
.A2(n_3242),
.B(n_3289),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3574),
.B(n_3327),
.Y(n_3829)
);

AOI31xp33_ASAP7_75t_L g3830 ( 
.A1(n_3409),
.A2(n_3020),
.A3(n_3289),
.B(n_3282),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3576),
.B(n_3299),
.Y(n_3831)
);

OA21x2_ASAP7_75t_L g3832 ( 
.A1(n_3584),
.A2(n_3238),
.B(n_3272),
.Y(n_3832)
);

OR2x2_ASAP7_75t_L g3833 ( 
.A(n_3546),
.B(n_3282),
.Y(n_3833)
);

OA21x2_ASAP7_75t_L g3834 ( 
.A1(n_3588),
.A2(n_3295),
.B(n_3233),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3588),
.Y(n_3835)
);

AND2x2_ASAP7_75t_L g3836 ( 
.A(n_3576),
.B(n_3198),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_L g3837 ( 
.A(n_3516),
.B(n_3236),
.Y(n_3837)
);

INVx1_ASAP7_75t_L g3838 ( 
.A(n_3503),
.Y(n_3838)
);

OAI21x1_ASAP7_75t_L g3839 ( 
.A1(n_3382),
.A2(n_3392),
.B(n_3385),
.Y(n_3839)
);

OR2x6_ASAP7_75t_L g3840 ( 
.A(n_3560),
.B(n_3145),
.Y(n_3840)
);

HB1xp67_ASAP7_75t_L g3841 ( 
.A(n_3351),
.Y(n_3841)
);

AO21x2_ASAP7_75t_L g3842 ( 
.A1(n_3483),
.A2(n_3460),
.B(n_3620),
.Y(n_3842)
);

OAI22xp33_ASAP7_75t_L g3843 ( 
.A1(n_3383),
.A2(n_3242),
.B1(n_3145),
.B2(n_3086),
.Y(n_3843)
);

INVx3_ASAP7_75t_L g3844 ( 
.A(n_3382),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3512),
.Y(n_3845)
);

INVx2_ASAP7_75t_L g3846 ( 
.A(n_3631),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3512),
.Y(n_3847)
);

OAI33xp33_ASAP7_75t_L g3848 ( 
.A1(n_3351),
.A2(n_3089),
.A3(n_3236),
.B1(n_3270),
.B2(n_3357),
.B3(n_3356),
.Y(n_3848)
);

INVx1_ASAP7_75t_L g3849 ( 
.A(n_3513),
.Y(n_3849)
);

INVxp67_ASAP7_75t_L g3850 ( 
.A(n_3384),
.Y(n_3850)
);

AO21x2_ASAP7_75t_L g3851 ( 
.A1(n_3554),
.A2(n_3593),
.B(n_3631),
.Y(n_3851)
);

AOI21x1_ASAP7_75t_L g3852 ( 
.A1(n_3527),
.A2(n_3514),
.B(n_3560),
.Y(n_3852)
);

OA21x2_ASAP7_75t_L g3853 ( 
.A1(n_3635),
.A2(n_3653),
.B(n_3647),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3594),
.B(n_3651),
.Y(n_3854)
);

NAND2x1_ASAP7_75t_L g3855 ( 
.A(n_3527),
.B(n_3514),
.Y(n_3855)
);

OR2x6_ASAP7_75t_L g3856 ( 
.A(n_3560),
.B(n_3569),
.Y(n_3856)
);

OR2x6_ASAP7_75t_L g3857 ( 
.A(n_3569),
.B(n_3514),
.Y(n_3857)
);

AOI22xp33_ASAP7_75t_L g3858 ( 
.A1(n_3408),
.A2(n_3570),
.B1(n_3579),
.B2(n_3440),
.Y(n_3858)
);

AND2x2_ASAP7_75t_L g3859 ( 
.A(n_3594),
.B(n_3651),
.Y(n_3859)
);

OA21x2_ASAP7_75t_L g3860 ( 
.A1(n_3635),
.A2(n_3653),
.B(n_3647),
.Y(n_3860)
);

INVx1_ASAP7_75t_L g3861 ( 
.A(n_3513),
.Y(n_3861)
);

AO21x2_ASAP7_75t_L g3862 ( 
.A1(n_3536),
.A2(n_3442),
.B(n_3615),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3522),
.Y(n_3863)
);

INVx2_ASAP7_75t_SL g3864 ( 
.A(n_3625),
.Y(n_3864)
);

AO21x2_ASAP7_75t_L g3865 ( 
.A1(n_3511),
.A2(n_3632),
.B(n_3565),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3522),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3655),
.Y(n_3867)
);

INVx2_ASAP7_75t_L g3868 ( 
.A(n_3655),
.Y(n_3868)
);

AOI33xp33_ASAP7_75t_L g3869 ( 
.A1(n_3363),
.A2(n_3378),
.A3(n_3410),
.B1(n_3488),
.B2(n_3664),
.B3(n_3558),
.Y(n_3869)
);

BUFx3_ASAP7_75t_L g3870 ( 
.A(n_3517),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_3408),
.A2(n_3569),
.B(n_3514),
.Y(n_3871)
);

NAND2xp5_ASAP7_75t_L g3872 ( 
.A(n_3487),
.B(n_3567),
.Y(n_3872)
);

INVx3_ASAP7_75t_L g3873 ( 
.A(n_3385),
.Y(n_3873)
);

AOI22xp5_ASAP7_75t_L g3874 ( 
.A1(n_3369),
.A2(n_3492),
.B1(n_3368),
.B2(n_3422),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3539),
.Y(n_3875)
);

BUFx2_ASAP7_75t_L g3876 ( 
.A(n_3527),
.Y(n_3876)
);

AO21x1_ASAP7_75t_SL g3877 ( 
.A1(n_3508),
.A2(n_3638),
.B(n_3660),
.Y(n_3877)
);

AO21x2_ASAP7_75t_L g3878 ( 
.A1(n_3511),
.A2(n_3658),
.B(n_3565),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3546),
.B(n_3665),
.Y(n_3879)
);

HB1xp67_ASAP7_75t_L g3880 ( 
.A(n_3356),
.Y(n_3880)
);

AND2x2_ASAP7_75t_L g3881 ( 
.A(n_3646),
.B(n_3385),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3539),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3541),
.Y(n_3883)
);

AND2x2_ASAP7_75t_L g3884 ( 
.A(n_3646),
.B(n_3392),
.Y(n_3884)
);

AOI22xp5_ASAP7_75t_L g3885 ( 
.A1(n_3492),
.A2(n_3368),
.B1(n_3415),
.B2(n_3409),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3541),
.Y(n_3886)
);

AO21x2_ASAP7_75t_L g3887 ( 
.A1(n_3511),
.A2(n_3658),
.B(n_3565),
.Y(n_3887)
);

INVx2_ASAP7_75t_L g3888 ( 
.A(n_3655),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3665),
.B(n_3609),
.Y(n_3889)
);

INVx1_ASAP7_75t_L g3890 ( 
.A(n_3559),
.Y(n_3890)
);

OR2x2_ASAP7_75t_L g3891 ( 
.A(n_3609),
.B(n_3637),
.Y(n_3891)
);

INVx1_ASAP7_75t_L g3892 ( 
.A(n_3559),
.Y(n_3892)
);

INVxp67_ASAP7_75t_L g3893 ( 
.A(n_3645),
.Y(n_3893)
);

INVxp67_ASAP7_75t_SL g3894 ( 
.A(n_3493),
.Y(n_3894)
);

AND2x2_ASAP7_75t_L g3895 ( 
.A(n_3392),
.B(n_3482),
.Y(n_3895)
);

AO21x2_ASAP7_75t_L g3896 ( 
.A1(n_3511),
.A2(n_3658),
.B(n_3565),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3655),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3357),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_3562),
.Y(n_3899)
);

OR2x2_ASAP7_75t_L g3900 ( 
.A(n_3637),
.B(n_3360),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3562),
.Y(n_3901)
);

AO21x2_ASAP7_75t_L g3902 ( 
.A1(n_3658),
.A2(n_3649),
.B(n_3644),
.Y(n_3902)
);

AND2x4_ASAP7_75t_SL g3903 ( 
.A(n_3440),
.B(n_3527),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3563),
.Y(n_3904)
);

HB1xp67_ASAP7_75t_L g3905 ( 
.A(n_3360),
.Y(n_3905)
);

BUFx2_ASAP7_75t_L g3906 ( 
.A(n_3569),
.Y(n_3906)
);

INVx1_ASAP7_75t_L g3907 ( 
.A(n_3563),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_L g3908 ( 
.A(n_3507),
.B(n_3441),
.Y(n_3908)
);

AND2x4_ASAP7_75t_SL g3909 ( 
.A(n_3440),
.B(n_3534),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3589),
.Y(n_3910)
);

OR2x6_ASAP7_75t_L g3911 ( 
.A(n_3569),
.B(n_3514),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3589),
.Y(n_3912)
);

OA21x2_ASAP7_75t_L g3913 ( 
.A1(n_3629),
.A2(n_3649),
.B(n_3644),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3595),
.Y(n_3914)
);

OR2x6_ASAP7_75t_L g3915 ( 
.A(n_3457),
.B(n_3389),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3482),
.Y(n_3916)
);

AND2x2_ASAP7_75t_L g3917 ( 
.A(n_3482),
.B(n_3531),
.Y(n_3917)
);

HB1xp67_ASAP7_75t_L g3918 ( 
.A(n_3586),
.Y(n_3918)
);

OAI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_3361),
.A2(n_3430),
.B(n_3426),
.Y(n_3919)
);

HB1xp67_ASAP7_75t_L g3920 ( 
.A(n_3603),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_3595),
.Y(n_3921)
);

INVx2_ASAP7_75t_L g3922 ( 
.A(n_3655),
.Y(n_3922)
);

AND2x2_ASAP7_75t_L g3923 ( 
.A(n_3531),
.B(n_3545),
.Y(n_3923)
);

INVx1_ASAP7_75t_SL g3924 ( 
.A(n_3411),
.Y(n_3924)
);

INVx1_ASAP7_75t_L g3925 ( 
.A(n_3598),
.Y(n_3925)
);

INVx2_ASAP7_75t_SL g3926 ( 
.A(n_3618),
.Y(n_3926)
);

HB1xp67_ASAP7_75t_L g3927 ( 
.A(n_3614),
.Y(n_3927)
);

AOI22xp33_ASAP7_75t_L g3928 ( 
.A1(n_3363),
.A2(n_3378),
.B1(n_3599),
.B2(n_3475),
.Y(n_3928)
);

INVxp67_ASAP7_75t_L g3929 ( 
.A(n_3449),
.Y(n_3929)
);

INVx1_ASAP7_75t_L g3930 ( 
.A(n_3598),
.Y(n_3930)
);

INVx1_ASAP7_75t_L g3931 ( 
.A(n_3605),
.Y(n_3931)
);

INVxp67_ASAP7_75t_SL g3932 ( 
.A(n_3581),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3605),
.Y(n_3933)
);

OAI21xp5_ASAP7_75t_L g3934 ( 
.A1(n_3500),
.A2(n_3486),
.B(n_3596),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3436),
.Y(n_3935)
);

OAI211xp5_ASAP7_75t_L g3936 ( 
.A1(n_3621),
.A2(n_3525),
.B(n_3580),
.C(n_3547),
.Y(n_3936)
);

BUFx6f_ASAP7_75t_L g3937 ( 
.A(n_3475),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3358),
.B(n_3435),
.Y(n_3938)
);

AOI22xp33_ASAP7_75t_L g3939 ( 
.A1(n_3858),
.A2(n_3457),
.B1(n_3517),
.B2(n_3617),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3679),
.Y(n_3940)
);

INVx3_ASAP7_75t_L g3941 ( 
.A(n_3747),
.Y(n_3941)
);

INVx1_ASAP7_75t_L g3942 ( 
.A(n_3679),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3813),
.B(n_3929),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_3779),
.B(n_3446),
.Y(n_3944)
);

AND2x2_ASAP7_75t_L g3945 ( 
.A(n_3862),
.B(n_3629),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3862),
.B(n_3727),
.Y(n_3946)
);

AND2x2_ASAP7_75t_L g3947 ( 
.A(n_3862),
.B(n_3604),
.Y(n_3947)
);

INVx2_ASAP7_75t_L g3948 ( 
.A(n_3717),
.Y(n_3948)
);

HB1xp67_ASAP7_75t_L g3949 ( 
.A(n_3765),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3717),
.Y(n_3950)
);

INVx2_ASAP7_75t_L g3951 ( 
.A(n_3717),
.Y(n_3951)
);

AND2x4_ASAP7_75t_SL g3952 ( 
.A(n_3668),
.B(n_3389),
.Y(n_3952)
);

INVx2_ASAP7_75t_L g3953 ( 
.A(n_3728),
.Y(n_3953)
);

AND2x2_ASAP7_75t_L g3954 ( 
.A(n_3727),
.B(n_3604),
.Y(n_3954)
);

AND2x2_ASAP7_75t_L g3955 ( 
.A(n_3802),
.B(n_3865),
.Y(n_3955)
);

INVx2_ASAP7_75t_L g3956 ( 
.A(n_3728),
.Y(n_3956)
);

AND2x2_ASAP7_75t_L g3957 ( 
.A(n_3802),
.B(n_3648),
.Y(n_3957)
);

AOI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3877),
.A2(n_3457),
.B1(n_3617),
.B2(n_3462),
.Y(n_3958)
);

AND2x2_ASAP7_75t_L g3959 ( 
.A(n_3865),
.B(n_3648),
.Y(n_3959)
);

AOI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3932),
.A2(n_3415),
.B1(n_3446),
.B2(n_3399),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3680),
.Y(n_3961)
);

HB1xp67_ASAP7_75t_L g3962 ( 
.A(n_3693),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_L g3963 ( 
.A(n_3841),
.B(n_3636),
.Y(n_3963)
);

NOR2xp33_ASAP7_75t_L g3964 ( 
.A(n_3779),
.B(n_3481),
.Y(n_3964)
);

BUFx2_ASAP7_75t_L g3965 ( 
.A(n_3817),
.Y(n_3965)
);

AND2x2_ASAP7_75t_L g3966 ( 
.A(n_3865),
.B(n_3650),
.Y(n_3966)
);

AND2x4_ASAP7_75t_L g3967 ( 
.A(n_3881),
.B(n_3531),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3680),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3874),
.B(n_3453),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3682),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3682),
.Y(n_3971)
);

AND2x2_ASAP7_75t_L g3972 ( 
.A(n_3854),
.B(n_3650),
.Y(n_3972)
);

INVx3_ASAP7_75t_L g3973 ( 
.A(n_3747),
.Y(n_3973)
);

AND2x2_ASAP7_75t_SL g3974 ( 
.A(n_3903),
.B(n_3621),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3728),
.Y(n_3975)
);

AOI22xp33_ASAP7_75t_L g3976 ( 
.A1(n_3877),
.A2(n_3457),
.B1(n_3462),
.B2(n_3661),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3817),
.Y(n_3977)
);

INVx1_ASAP7_75t_L g3978 ( 
.A(n_3683),
.Y(n_3978)
);

AND2x4_ASAP7_75t_L g3979 ( 
.A(n_3881),
.B(n_3545),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3854),
.B(n_3639),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3859),
.B(n_3639),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3683),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3880),
.B(n_3636),
.Y(n_3983)
);

AND2x4_ASAP7_75t_SL g3984 ( 
.A(n_3668),
.B(n_3389),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3898),
.B(n_3640),
.Y(n_3985)
);

HB1xp67_ASAP7_75t_L g3986 ( 
.A(n_3749),
.Y(n_3986)
);

AOI22xp33_ASAP7_75t_SL g3987 ( 
.A1(n_3795),
.A2(n_3621),
.B1(n_3457),
.B2(n_3506),
.Y(n_3987)
);

AND2x2_ASAP7_75t_L g3988 ( 
.A(n_3859),
.B(n_3591),
.Y(n_3988)
);

AND2x2_ASAP7_75t_L g3989 ( 
.A(n_3673),
.B(n_3591),
.Y(n_3989)
);

AND2x2_ASAP7_75t_L g3990 ( 
.A(n_3673),
.B(n_3591),
.Y(n_3990)
);

AND2x2_ASAP7_75t_L g3991 ( 
.A(n_3673),
.B(n_3591),
.Y(n_3991)
);

AND2x2_ASAP7_75t_L g3992 ( 
.A(n_3894),
.B(n_3591),
.Y(n_3992)
);

INVx2_ASAP7_75t_L g3993 ( 
.A(n_3791),
.Y(n_3993)
);

INVx2_ASAP7_75t_L g3994 ( 
.A(n_3791),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3678),
.A2(n_3520),
.B1(n_3621),
.B2(n_3403),
.Y(n_3995)
);

INVxp67_ASAP7_75t_SL g3996 ( 
.A(n_3678),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3692),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_3884),
.B(n_3545),
.Y(n_3998)
);

INVx2_ASAP7_75t_L g3999 ( 
.A(n_3791),
.Y(n_3999)
);

INVx3_ASAP7_75t_L g4000 ( 
.A(n_3747),
.Y(n_4000)
);

BUFx3_ASAP7_75t_L g4001 ( 
.A(n_3779),
.Y(n_4001)
);

AND2x2_ASAP7_75t_L g4002 ( 
.A(n_3884),
.B(n_3608),
.Y(n_4002)
);

INVxp67_ASAP7_75t_L g4003 ( 
.A(n_3746),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3720),
.B(n_3608),
.Y(n_4004)
);

INVx1_ASAP7_75t_L g4005 ( 
.A(n_3692),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_3936),
.A2(n_3476),
.B1(n_3582),
.B2(n_3481),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3720),
.B(n_3619),
.Y(n_4007)
);

AND3x1_ASAP7_75t_L g4008 ( 
.A(n_3874),
.B(n_3439),
.C(n_3666),
.Y(n_4008)
);

BUFx2_ASAP7_75t_L g4009 ( 
.A(n_3817),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_3792),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3695),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3720),
.B(n_3619),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_3905),
.B(n_3642),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3720),
.B(n_3622),
.Y(n_4014)
);

INVx3_ASAP7_75t_L g4015 ( 
.A(n_3729),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3791),
.Y(n_4016)
);

INVx2_ASAP7_75t_L g4017 ( 
.A(n_3811),
.Y(n_4017)
);

HB1xp67_ASAP7_75t_L g4018 ( 
.A(n_3797),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3720),
.B(n_3622),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3811),
.Y(n_4020)
);

INVx2_ASAP7_75t_L g4021 ( 
.A(n_3811),
.Y(n_4021)
);

OAI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3830),
.A2(n_3641),
.B1(n_3611),
.B2(n_3616),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_L g4023 ( 
.A(n_3676),
.B(n_3396),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3856),
.B(n_3677),
.Y(n_4024)
);

INVx2_ASAP7_75t_L g4025 ( 
.A(n_3811),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3695),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3697),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3815),
.Y(n_4028)
);

INVx2_ASAP7_75t_L g4029 ( 
.A(n_3815),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_3908),
.B(n_3837),
.Y(n_4030)
);

INVx1_ASAP7_75t_L g4031 ( 
.A(n_3697),
.Y(n_4031)
);

BUFx2_ASAP7_75t_L g4032 ( 
.A(n_3694),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3703),
.Y(n_4033)
);

INVx1_ASAP7_75t_L g4034 ( 
.A(n_3703),
.Y(n_4034)
);

NOR2xp33_ASAP7_75t_L g4035 ( 
.A(n_3786),
.B(n_3371),
.Y(n_4035)
);

INVx4_ASAP7_75t_L g4036 ( 
.A(n_3870),
.Y(n_4036)
);

INVx3_ASAP7_75t_L g4037 ( 
.A(n_3729),
.Y(n_4037)
);

NOR2xp33_ASAP7_75t_L g4038 ( 
.A(n_3870),
.B(n_3371),
.Y(n_4038)
);

NOR2xp33_ASAP7_75t_L g4039 ( 
.A(n_3870),
.B(n_3395),
.Y(n_4039)
);

AOI22xp33_ASAP7_75t_L g4040 ( 
.A1(n_3934),
.A2(n_3520),
.B1(n_3401),
.B2(n_3403),
.Y(n_4040)
);

INVx1_ASAP7_75t_L g4041 ( 
.A(n_3704),
.Y(n_4041)
);

INVx2_ASAP7_75t_L g4042 ( 
.A(n_3815),
.Y(n_4042)
);

INVx2_ASAP7_75t_L g4043 ( 
.A(n_3815),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3704),
.Y(n_4044)
);

OR2x2_ASAP7_75t_L g4045 ( 
.A(n_3672),
.B(n_3434),
.Y(n_4045)
);

NOR2x1_ASAP7_75t_L g4046 ( 
.A(n_3671),
.B(n_3389),
.Y(n_4046)
);

AND2x2_ASAP7_75t_L g4047 ( 
.A(n_3856),
.B(n_3630),
.Y(n_4047)
);

AND2x4_ASAP7_75t_L g4048 ( 
.A(n_3804),
.B(n_3434),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_3804),
.B(n_3434),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_3825),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3768),
.B(n_3417),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3707),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3856),
.B(n_3630),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_L g4054 ( 
.A(n_3672),
.B(n_3674),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3856),
.B(n_3634),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3707),
.Y(n_4056)
);

NOR2xp67_ASAP7_75t_L g4057 ( 
.A(n_3871),
.B(n_3618),
.Y(n_4057)
);

OR2x2_ASAP7_75t_L g4058 ( 
.A(n_3674),
.B(n_3434),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3719),
.Y(n_4059)
);

INVxp67_ASAP7_75t_L g4060 ( 
.A(n_3746),
.Y(n_4060)
);

NOR2xp33_ASAP7_75t_L g4061 ( 
.A(n_3937),
.B(n_3398),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3719),
.Y(n_4062)
);

BUFx6f_ASAP7_75t_L g4063 ( 
.A(n_3937),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_3721),
.Y(n_4064)
);

OR2x2_ASAP7_75t_L g4065 ( 
.A(n_3722),
.B(n_3434),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_3721),
.Y(n_4066)
);

HB1xp67_ASAP7_75t_L g4067 ( 
.A(n_3913),
.Y(n_4067)
);

HB1xp67_ASAP7_75t_L g4068 ( 
.A(n_3913),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3726),
.Y(n_4069)
);

INVx2_ASAP7_75t_L g4070 ( 
.A(n_3825),
.Y(n_4070)
);

INVx2_ASAP7_75t_SL g4071 ( 
.A(n_3729),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3913),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3856),
.B(n_3634),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3804),
.B(n_3375),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3825),
.Y(n_4075)
);

INVx2_ASAP7_75t_SL g4076 ( 
.A(n_3684),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3726),
.Y(n_4077)
);

BUFx3_ASAP7_75t_L g4078 ( 
.A(n_3694),
.Y(n_4078)
);

INVx2_ASAP7_75t_L g4079 ( 
.A(n_3825),
.Y(n_4079)
);

AND2x4_ASAP7_75t_L g4080 ( 
.A(n_3804),
.B(n_3375),
.Y(n_4080)
);

AND2x2_ASAP7_75t_L g4081 ( 
.A(n_3677),
.B(n_3515),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3736),
.Y(n_4082)
);

HB1xp67_ASAP7_75t_L g4083 ( 
.A(n_3918),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3677),
.B(n_3515),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_3832),
.Y(n_4085)
);

INVx1_ASAP7_75t_L g4086 ( 
.A(n_3736),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3740),
.Y(n_4087)
);

AND2x2_ASAP7_75t_L g4088 ( 
.A(n_3857),
.B(n_3519),
.Y(n_4088)
);

AND2x2_ASAP7_75t_L g4089 ( 
.A(n_3857),
.B(n_3519),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3857),
.B(n_3656),
.Y(n_4090)
);

AND2x4_ASAP7_75t_L g4091 ( 
.A(n_3864),
.B(n_3375),
.Y(n_4091)
);

BUFx6f_ASAP7_75t_L g4092 ( 
.A(n_3937),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_3737),
.B(n_3419),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3857),
.B(n_3656),
.Y(n_4094)
);

AND2x2_ASAP7_75t_L g4095 ( 
.A(n_3857),
.B(n_3656),
.Y(n_4095)
);

INVx1_ASAP7_75t_L g4096 ( 
.A(n_3740),
.Y(n_4096)
);

INVx1_ASAP7_75t_SL g4097 ( 
.A(n_3924),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3741),
.B(n_3662),
.Y(n_4098)
);

INVx3_ASAP7_75t_L g4099 ( 
.A(n_3684),
.Y(n_4099)
);

AND2x4_ASAP7_75t_L g4100 ( 
.A(n_3864),
.B(n_3375),
.Y(n_4100)
);

NOR2x1_ASAP7_75t_L g4101 ( 
.A(n_3671),
.B(n_3389),
.Y(n_4101)
);

BUFx2_ASAP7_75t_L g4102 ( 
.A(n_3694),
.Y(n_4102)
);

AND2x2_ASAP7_75t_L g4103 ( 
.A(n_3911),
.B(n_3521),
.Y(n_4103)
);

INVx2_ASAP7_75t_SL g4104 ( 
.A(n_3684),
.Y(n_4104)
);

AOI22xp33_ASAP7_75t_L g4105 ( 
.A1(n_3850),
.A2(n_3401),
.B1(n_3549),
.B2(n_3505),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_3920),
.Y(n_4106)
);

OAI22xp33_ASAP7_75t_L g4107 ( 
.A1(n_3830),
.A2(n_3623),
.B1(n_3549),
.B2(n_3547),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_3913),
.Y(n_4108)
);

INVx8_ASAP7_75t_L g4109 ( 
.A(n_3937),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_3911),
.B(n_3521),
.Y(n_4110)
);

INVx1_ASAP7_75t_L g4111 ( 
.A(n_3752),
.Y(n_4111)
);

INVx2_ASAP7_75t_L g4112 ( 
.A(n_3832),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_3752),
.Y(n_4113)
);

INVx3_ASAP7_75t_L g4114 ( 
.A(n_3684),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3722),
.B(n_3662),
.Y(n_4115)
);

AND2x2_ASAP7_75t_L g4116 ( 
.A(n_3911),
.B(n_3530),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_3760),
.Y(n_4117)
);

CKINVDCx20_ASAP7_75t_R g4118 ( 
.A(n_3730),
.Y(n_4118)
);

AOI22xp33_ASAP7_75t_L g4119 ( 
.A1(n_3919),
.A2(n_3505),
.B1(n_3530),
.B2(n_3421),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_3760),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_3761),
.Y(n_4121)
);

BUFx6f_ASAP7_75t_L g4122 ( 
.A(n_3937),
.Y(n_4122)
);

INVx2_ASAP7_75t_L g4123 ( 
.A(n_3832),
.Y(n_4123)
);

INVx2_ASAP7_75t_L g4124 ( 
.A(n_3832),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_3761),
.Y(n_4125)
);

INVx3_ASAP7_75t_L g4126 ( 
.A(n_3685),
.Y(n_4126)
);

INVx1_ASAP7_75t_L g4127 ( 
.A(n_3762),
.Y(n_4127)
);

INVx2_ASAP7_75t_L g4128 ( 
.A(n_3834),
.Y(n_4128)
);

AND2x4_ASAP7_75t_SL g4129 ( 
.A(n_3668),
.B(n_3497),
.Y(n_4129)
);

AND2x2_ASAP7_75t_L g4130 ( 
.A(n_3911),
.B(n_3585),
.Y(n_4130)
);

INVx1_ASAP7_75t_L g4131 ( 
.A(n_3762),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_3911),
.B(n_3585),
.Y(n_4132)
);

AND2x2_ASAP7_75t_L g4133 ( 
.A(n_3805),
.B(n_3585),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3764),
.Y(n_4134)
);

CKINVDCx5p33_ASAP7_75t_R g4135 ( 
.A(n_3753),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_3764),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3771),
.Y(n_4137)
);

OR2x2_ASAP7_75t_L g4138 ( 
.A(n_3819),
.B(n_3354),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3938),
.B(n_3467),
.Y(n_4139)
);

INVx1_ASAP7_75t_L g4140 ( 
.A(n_3771),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3777),
.Y(n_4141)
);

AND2x4_ASAP7_75t_L g4142 ( 
.A(n_3851),
.B(n_3618),
.Y(n_4142)
);

INVxp67_ASAP7_75t_SL g4143 ( 
.A(n_3701),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_3777),
.Y(n_4144)
);

INVx3_ASAP7_75t_L g4145 ( 
.A(n_3685),
.Y(n_4145)
);

NAND2xp5_ASAP7_75t_SL g4146 ( 
.A(n_3885),
.B(n_3420),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_3834),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_3834),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_3819),
.B(n_3354),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_3669),
.B(n_3585),
.Y(n_4150)
);

OAI22xp5_ASAP7_75t_L g4151 ( 
.A1(n_3755),
.A2(n_3612),
.B1(n_3602),
.B2(n_3394),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3893),
.B(n_3927),
.Y(n_4152)
);

AND2x2_ASAP7_75t_L g4153 ( 
.A(n_3669),
.B(n_3585),
.Y(n_4153)
);

NAND2xp5_ASAP7_75t_L g4154 ( 
.A(n_3829),
.B(n_3366),
.Y(n_4154)
);

NOR2x1_ASAP7_75t_L g4155 ( 
.A(n_3732),
.B(n_3552),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3788),
.Y(n_4156)
);

AND2x4_ASAP7_75t_L g4157 ( 
.A(n_3851),
.B(n_3618),
.Y(n_4157)
);

INVx3_ASAP7_75t_L g4158 ( 
.A(n_3685),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_3834),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_3788),
.Y(n_4160)
);

AND2x2_ASAP7_75t_L g4161 ( 
.A(n_3700),
.B(n_3592),
.Y(n_4161)
);

OAI21xp33_ASAP7_75t_L g4162 ( 
.A1(n_3869),
.A2(n_3459),
.B(n_3355),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_3700),
.B(n_3592),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_3790),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_3853),
.Y(n_4165)
);

AND2x2_ASAP7_75t_L g4166 ( 
.A(n_3713),
.B(n_3592),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4078),
.Y(n_4167)
);

OAI21xp33_ASAP7_75t_L g4168 ( 
.A1(n_3996),
.A2(n_3755),
.B(n_3885),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_3962),
.Y(n_4169)
);

OAI22xp5_ASAP7_75t_L g4170 ( 
.A1(n_4006),
.A2(n_3928),
.B1(n_3924),
.B2(n_3774),
.Y(n_4170)
);

AND2x4_ASAP7_75t_L g4171 ( 
.A(n_4155),
.B(n_3909),
.Y(n_4171)
);

INVx2_ASAP7_75t_SL g4172 ( 
.A(n_4001),
.Y(n_4172)
);

AOI22xp5_ASAP7_75t_L g4173 ( 
.A1(n_4008),
.A2(n_3909),
.B1(n_3711),
.B2(n_3725),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_3962),
.Y(n_4174)
);

OR2x6_ASAP7_75t_L g4175 ( 
.A(n_4109),
.B(n_3937),
.Y(n_4175)
);

INVx3_ASAP7_75t_L g4176 ( 
.A(n_4001),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4078),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4002),
.B(n_3972),
.Y(n_4178)
);

BUFx3_ASAP7_75t_L g4179 ( 
.A(n_4001),
.Y(n_4179)
);

AND2x4_ASAP7_75t_L g4180 ( 
.A(n_4155),
.B(n_4078),
.Y(n_4180)
);

INVx3_ASAP7_75t_L g4181 ( 
.A(n_4142),
.Y(n_4181)
);

AOI222xp33_ASAP7_75t_L g4182 ( 
.A1(n_3996),
.A2(n_3780),
.B1(n_3848),
.B2(n_3766),
.C1(n_3716),
.C2(n_3698),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_4063),
.Y(n_4183)
);

INVx2_ASAP7_75t_L g4184 ( 
.A(n_4063),
.Y(n_4184)
);

NAND3xp33_ASAP7_75t_L g4185 ( 
.A(n_3987),
.B(n_3995),
.C(n_4006),
.Y(n_4185)
);

OAI22xp5_ASAP7_75t_L g4186 ( 
.A1(n_4008),
.A2(n_3976),
.B1(n_3958),
.B2(n_4040),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_SL g4187 ( 
.A(n_3964),
.B(n_3398),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3986),
.Y(n_4188)
);

AOI31xp33_ASAP7_75t_L g4189 ( 
.A1(n_4146),
.A2(n_3794),
.A3(n_3770),
.B(n_3787),
.Y(n_4189)
);

OAI211xp5_ASAP7_75t_L g4190 ( 
.A1(n_3987),
.A2(n_4143),
.B(n_3946),
.C(n_4101),
.Y(n_4190)
);

BUFx3_ASAP7_75t_L g4191 ( 
.A(n_4118),
.Y(n_4191)
);

AND2x4_ASAP7_75t_SL g4192 ( 
.A(n_4074),
.B(n_4080),
.Y(n_4192)
);

AO221x2_ASAP7_75t_L g4193 ( 
.A1(n_4151),
.A2(n_3843),
.B1(n_3753),
.B2(n_3852),
.C(n_3903),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3986),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_4097),
.B(n_3732),
.Y(n_4195)
);

OAI221xp5_ASAP7_75t_SL g4196 ( 
.A1(n_4107),
.A2(n_3781),
.B1(n_3800),
.B2(n_3766),
.C(n_3733),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4010),
.Y(n_4197)
);

INVxp67_ASAP7_75t_SL g4198 ( 
.A(n_3947),
.Y(n_4198)
);

OAI22xp33_ASAP7_75t_L g4199 ( 
.A1(n_4143),
.A2(n_3733),
.B1(n_3691),
.B2(n_3734),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4010),
.Y(n_4200)
);

HB1xp67_ASAP7_75t_L g4201 ( 
.A(n_4067),
.Y(n_4201)
);

BUFx2_ASAP7_75t_L g4202 ( 
.A(n_3965),
.Y(n_4202)
);

INVx1_ASAP7_75t_L g4203 ( 
.A(n_4018),
.Y(n_4203)
);

INVx1_ASAP7_75t_L g4204 ( 
.A(n_4018),
.Y(n_4204)
);

OAI211xp5_ASAP7_75t_SL g4205 ( 
.A1(n_4162),
.A2(n_3821),
.B(n_3781),
.C(n_3800),
.Y(n_4205)
);

OAI22xp5_ASAP7_75t_L g4206 ( 
.A1(n_3960),
.A2(n_3909),
.B1(n_3734),
.B2(n_3725),
.Y(n_4206)
);

HB1xp67_ASAP7_75t_L g4207 ( 
.A(n_4067),
.Y(n_4207)
);

INVx1_ASAP7_75t_SL g4208 ( 
.A(n_4097),
.Y(n_4208)
);

OA21x2_ASAP7_75t_L g4209 ( 
.A1(n_4068),
.A2(n_3839),
.B(n_3713),
.Y(n_4209)
);

AND2x2_ASAP7_75t_L g4210 ( 
.A(n_4002),
.B(n_3751),
.Y(n_4210)
);

BUFx3_ASAP7_75t_L g4211 ( 
.A(n_3965),
.Y(n_4211)
);

AOI22xp33_ASAP7_75t_SL g4212 ( 
.A1(n_4151),
.A2(n_3706),
.B1(n_3906),
.B2(n_3691),
.Y(n_4212)
);

OAI221xp5_ASAP7_75t_L g4213 ( 
.A1(n_3960),
.A2(n_4162),
.B1(n_3939),
.B2(n_3969),
.C(n_4119),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3940),
.Y(n_4214)
);

NOR2xp33_ASAP7_75t_R g4215 ( 
.A(n_4135),
.B(n_3476),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3940),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_4063),
.Y(n_4217)
);

NOR2xp33_ASAP7_75t_L g4218 ( 
.A(n_3944),
.B(n_4036),
.Y(n_4218)
);

INVx4_ASAP7_75t_L g4219 ( 
.A(n_4036),
.Y(n_4219)
);

AOI221xp5_ASAP7_75t_L g4220 ( 
.A1(n_4022),
.A2(n_3821),
.B1(n_3818),
.B2(n_3906),
.C(n_3801),
.Y(n_4220)
);

OA211x2_ASAP7_75t_L g4221 ( 
.A1(n_4061),
.A2(n_3855),
.B(n_3872),
.C(n_3753),
.Y(n_4221)
);

AOI22xp33_ASAP7_75t_L g4222 ( 
.A1(n_4051),
.A2(n_3706),
.B1(n_3691),
.B2(n_3842),
.Y(n_4222)
);

OAI221xp5_ASAP7_75t_L g4223 ( 
.A1(n_4051),
.A2(n_3855),
.B1(n_3915),
.B2(n_3876),
.C(n_3754),
.Y(n_4223)
);

OAI211xp5_ASAP7_75t_L g4224 ( 
.A1(n_3946),
.A2(n_3876),
.B(n_3706),
.C(n_3852),
.Y(n_4224)
);

NOR2xp33_ASAP7_75t_R g4225 ( 
.A(n_4036),
.B(n_3495),
.Y(n_4225)
);

OAI22xp5_ASAP7_75t_L g4226 ( 
.A1(n_4046),
.A2(n_3732),
.B1(n_3691),
.B2(n_3915),
.Y(n_4226)
);

AND2x2_ASAP7_75t_L g4227 ( 
.A(n_3972),
.B(n_3751),
.Y(n_4227)
);

OAI221xp5_ASAP7_75t_L g4228 ( 
.A1(n_4046),
.A2(n_3915),
.B1(n_3754),
.B2(n_3812),
.C(n_3706),
.Y(n_4228)
);

AOI33xp33_ASAP7_75t_L g4229 ( 
.A1(n_3992),
.A2(n_3903),
.A3(n_3731),
.B1(n_3744),
.B2(n_3710),
.B3(n_3715),
.Y(n_4229)
);

NAND3xp33_ASAP7_75t_L g4230 ( 
.A(n_4101),
.B(n_3668),
.C(n_3767),
.Y(n_4230)
);

BUFx3_ASAP7_75t_L g4231 ( 
.A(n_3977),
.Y(n_4231)
);

AND2x4_ASAP7_75t_L g4232 ( 
.A(n_4032),
.B(n_3668),
.Y(n_4232)
);

NAND3xp33_ASAP7_75t_L g4233 ( 
.A(n_3949),
.B(n_3668),
.C(n_3767),
.Y(n_4233)
);

NAND2xp5_ASAP7_75t_L g4234 ( 
.A(n_3977),
.B(n_3767),
.Y(n_4234)
);

HB1xp67_ASAP7_75t_L g4235 ( 
.A(n_4068),
.Y(n_4235)
);

AOI221xp5_ASAP7_75t_L g4236 ( 
.A1(n_3943),
.A2(n_3842),
.B1(n_3753),
.B2(n_3731),
.C(n_3744),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_3942),
.Y(n_4237)
);

HB1xp67_ASAP7_75t_L g4238 ( 
.A(n_4072),
.Y(n_4238)
);

OAI211xp5_ASAP7_75t_L g4239 ( 
.A1(n_3947),
.A2(n_3989),
.B(n_3991),
.C(n_3990),
.Y(n_4239)
);

AOI22xp5_ASAP7_75t_L g4240 ( 
.A1(n_3957),
.A2(n_3842),
.B1(n_3785),
.B2(n_3767),
.Y(n_4240)
);

AOI21x1_ASAP7_75t_L g4241 ( 
.A1(n_4009),
.A2(n_3926),
.B(n_3917),
.Y(n_4241)
);

AND2x2_ASAP7_75t_L g4242 ( 
.A(n_3980),
.B(n_3710),
.Y(n_4242)
);

OA21x2_ASAP7_75t_L g4243 ( 
.A1(n_4072),
.A2(n_3839),
.B(n_3688),
.Y(n_4243)
);

NOR2xp67_ASAP7_75t_L g4244 ( 
.A(n_3945),
.B(n_3926),
.Y(n_4244)
);

AOI22xp33_ASAP7_75t_L g4245 ( 
.A1(n_3974),
.A2(n_3828),
.B1(n_3782),
.B2(n_3785),
.Y(n_4245)
);

AOI22xp33_ASAP7_75t_L g4246 ( 
.A1(n_3974),
.A2(n_3828),
.B1(n_3782),
.B2(n_3785),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3942),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_3980),
.B(n_3715),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_4009),
.Y(n_4249)
);

NOR4xp25_ASAP7_75t_L g4250 ( 
.A(n_3955),
.B(n_3757),
.C(n_3772),
.D(n_3763),
.Y(n_4250)
);

AND2x2_ASAP7_75t_L g4251 ( 
.A(n_3981),
.B(n_3757),
.Y(n_4251)
);

OAI211xp5_ASAP7_75t_L g4252 ( 
.A1(n_3989),
.A2(n_3681),
.B(n_3686),
.C(n_3785),
.Y(n_4252)
);

HB1xp67_ASAP7_75t_L g4253 ( 
.A(n_4108),
.Y(n_4253)
);

NOR3xp33_ASAP7_75t_L g4254 ( 
.A(n_4036),
.B(n_3844),
.C(n_3823),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_3961),
.Y(n_4255)
);

OR2x6_ASAP7_75t_L g4256 ( 
.A(n_4109),
.B(n_3767),
.Y(n_4256)
);

OR2x2_ASAP7_75t_L g4257 ( 
.A(n_4152),
.B(n_3889),
.Y(n_4257)
);

OAI332xp33_ASAP7_75t_L g4258 ( 
.A1(n_4045),
.A2(n_3879),
.A3(n_3690),
.B1(n_3696),
.B2(n_3699),
.B3(n_3702),
.C1(n_3705),
.C2(n_3708),
.Y(n_4258)
);

AND2x2_ASAP7_75t_L g4259 ( 
.A(n_3981),
.B(n_3957),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3961),
.Y(n_4260)
);

NOR2xp33_ASAP7_75t_L g4261 ( 
.A(n_4038),
.B(n_3451),
.Y(n_4261)
);

AOI22xp5_ASAP7_75t_L g4262 ( 
.A1(n_3988),
.A2(n_3785),
.B1(n_3767),
.B2(n_3915),
.Y(n_4262)
);

OAI22xp5_ASAP7_75t_L g4263 ( 
.A1(n_4105),
.A2(n_3915),
.B1(n_3523),
.B2(n_3602),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_3954),
.B(n_4074),
.Y(n_4264)
);

AOI22xp5_ASAP7_75t_L g4265 ( 
.A1(n_3988),
.A2(n_3785),
.B1(n_3806),
.B2(n_3759),
.Y(n_4265)
);

NAND3xp33_ASAP7_75t_L g4266 ( 
.A(n_3990),
.B(n_3782),
.C(n_3840),
.Y(n_4266)
);

OR2x2_ASAP7_75t_L g4267 ( 
.A(n_4152),
.B(n_3889),
.Y(n_4267)
);

OAI211xp5_ASAP7_75t_L g4268 ( 
.A1(n_3991),
.A2(n_3681),
.B(n_3686),
.C(n_3675),
.Y(n_4268)
);

AND2x2_ASAP7_75t_L g4269 ( 
.A(n_3954),
.B(n_3759),
.Y(n_4269)
);

AOI21xp5_ASAP7_75t_L g4270 ( 
.A1(n_3974),
.A2(n_3840),
.B(n_3782),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4063),
.Y(n_4271)
);

OR2x2_ASAP7_75t_L g4272 ( 
.A(n_3943),
.B(n_3879),
.Y(n_4272)
);

OAI221xp5_ASAP7_75t_L g4273 ( 
.A1(n_4093),
.A2(n_3840),
.B1(n_3782),
.B2(n_3806),
.C(n_3748),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4030),
.B(n_3756),
.Y(n_4274)
);

OAI332xp33_ASAP7_75t_L g4275 ( 
.A1(n_4045),
.A2(n_3702),
.A3(n_3699),
.B1(n_3696),
.B2(n_3690),
.B3(n_3689),
.C1(n_3705),
.C2(n_3708),
.Y(n_4275)
);

INVx1_ASAP7_75t_L g4276 ( 
.A(n_3968),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4063),
.Y(n_4277)
);

BUFx3_ASAP7_75t_L g4278 ( 
.A(n_4032),
.Y(n_4278)
);

INVx1_ASAP7_75t_L g4279 ( 
.A(n_3968),
.Y(n_4279)
);

NOR3xp33_ASAP7_75t_SL g4280 ( 
.A(n_4039),
.B(n_3495),
.C(n_3451),
.Y(n_4280)
);

BUFx2_ASAP7_75t_L g4281 ( 
.A(n_4102),
.Y(n_4281)
);

OR2x2_ASAP7_75t_L g4282 ( 
.A(n_4030),
.B(n_3756),
.Y(n_4282)
);

INVx1_ASAP7_75t_L g4283 ( 
.A(n_3970),
.Y(n_4283)
);

NOR2x1_ASAP7_75t_SL g4284 ( 
.A(n_3945),
.B(n_3851),
.Y(n_4284)
);

AND2x2_ASAP7_75t_L g4285 ( 
.A(n_4074),
.B(n_3763),
.Y(n_4285)
);

AOI221xp5_ASAP7_75t_L g4286 ( 
.A1(n_4093),
.A2(n_3772),
.B1(n_3750),
.B2(n_3748),
.C(n_3745),
.Y(n_4286)
);

AND2x4_ASAP7_75t_SL g4287 ( 
.A(n_4074),
.B(n_4080),
.Y(n_4287)
);

INVx1_ASAP7_75t_L g4288 ( 
.A(n_3970),
.Y(n_4288)
);

NOR3xp33_ASAP7_75t_L g4289 ( 
.A(n_4102),
.B(n_3844),
.C(n_3823),
.Y(n_4289)
);

INVx2_ASAP7_75t_L g4290 ( 
.A(n_4063),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3971),
.Y(n_4291)
);

INVx1_ASAP7_75t_L g4292 ( 
.A(n_3971),
.Y(n_4292)
);

NAND3xp33_ASAP7_75t_L g4293 ( 
.A(n_4083),
.B(n_3840),
.C(n_3681),
.Y(n_4293)
);

OR2x2_ASAP7_75t_L g4294 ( 
.A(n_4054),
.B(n_3758),
.Y(n_4294)
);

OAI21xp5_ASAP7_75t_L g4295 ( 
.A1(n_4057),
.A2(n_3688),
.B(n_3807),
.Y(n_4295)
);

NAND2xp33_ASAP7_75t_R g4296 ( 
.A(n_3955),
.B(n_3489),
.Y(n_4296)
);

NOR4xp25_ASAP7_75t_SL g4297 ( 
.A(n_3978),
.B(n_3523),
.C(n_3612),
.D(n_3931),
.Y(n_4297)
);

BUFx3_ASAP7_75t_L g4298 ( 
.A(n_4109),
.Y(n_4298)
);

NAND2xp5_ASAP7_75t_L g4299 ( 
.A(n_4106),
.B(n_3836),
.Y(n_4299)
);

OAI22xp5_ASAP7_75t_L g4300 ( 
.A1(n_4058),
.A2(n_3840),
.B1(n_3497),
.B2(n_3394),
.Y(n_4300)
);

BUFx3_ASAP7_75t_L g4301 ( 
.A(n_4109),
.Y(n_4301)
);

BUFx3_ASAP7_75t_L g4302 ( 
.A(n_4109),
.Y(n_4302)
);

AND2x4_ASAP7_75t_L g4303 ( 
.A(n_4080),
.B(n_3878),
.Y(n_4303)
);

NAND2xp5_ASAP7_75t_L g4304 ( 
.A(n_4003),
.B(n_3836),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_4080),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4092),
.Y(n_4306)
);

AOI222xp33_ASAP7_75t_L g4307 ( 
.A1(n_3992),
.A2(n_3820),
.B1(n_3831),
.B2(n_3745),
.C1(n_3917),
.C2(n_3895),
.Y(n_4307)
);

AOI22xp33_ASAP7_75t_L g4308 ( 
.A1(n_4133),
.A2(n_3681),
.B1(n_3686),
.B2(n_3750),
.Y(n_4308)
);

INVx2_ASAP7_75t_L g4309 ( 
.A(n_4092),
.Y(n_4309)
);

AOI33xp33_ASAP7_75t_L g4310 ( 
.A1(n_4133),
.A2(n_3820),
.A3(n_3933),
.B1(n_3931),
.B2(n_3930),
.B3(n_3790),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_R g4311 ( 
.A(n_4035),
.B(n_3553),
.Y(n_4311)
);

INVxp67_ASAP7_75t_SL g4312 ( 
.A(n_4099),
.Y(n_4312)
);

OAI211xp5_ASAP7_75t_SL g4313 ( 
.A1(n_4058),
.A2(n_3823),
.B(n_3844),
.C(n_3873),
.Y(n_4313)
);

NOR2xp33_ASAP7_75t_R g4314 ( 
.A(n_4092),
.B(n_3553),
.Y(n_4314)
);

NAND3xp33_ASAP7_75t_L g4315 ( 
.A(n_4003),
.B(n_3686),
.C(n_3900),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_4108),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_L g4317 ( 
.A(n_4060),
.B(n_3831),
.Y(n_4317)
);

NAND4xp25_ASAP7_75t_L g4318 ( 
.A(n_4057),
.B(n_3895),
.C(n_3923),
.D(n_3823),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_3978),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_4092),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4091),
.B(n_3923),
.Y(n_4321)
);

OAI33xp33_ASAP7_75t_L g4322 ( 
.A1(n_4060),
.A2(n_3900),
.A3(n_3933),
.B1(n_3930),
.B2(n_3925),
.B3(n_3808),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3982),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4091),
.B(n_3473),
.Y(n_4324)
);

CKINVDCx16_ASAP7_75t_R g4325 ( 
.A(n_4091),
.Y(n_4325)
);

HB1xp67_ASAP7_75t_L g4326 ( 
.A(n_4092),
.Y(n_4326)
);

OR2x2_ASAP7_75t_L g4327 ( 
.A(n_4054),
.B(n_3758),
.Y(n_4327)
);

AOI22xp33_ASAP7_75t_L g4328 ( 
.A1(n_4065),
.A2(n_3750),
.B1(n_3675),
.B2(n_3687),
.Y(n_4328)
);

INVx2_ASAP7_75t_L g4329 ( 
.A(n_4092),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4122),
.Y(n_4330)
);

OAI22xp5_ASAP7_75t_L g4331 ( 
.A1(n_4065),
.A2(n_3497),
.B1(n_3452),
.B2(n_3381),
.Y(n_4331)
);

OAI22xp33_ASAP7_75t_L g4332 ( 
.A1(n_4122),
.A2(n_3497),
.B1(n_3618),
.B2(n_3687),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_3982),
.Y(n_4333)
);

AOI21xp5_ASAP7_75t_L g4334 ( 
.A1(n_4024),
.A2(n_3807),
.B(n_3685),
.Y(n_4334)
);

OR2x6_ASAP7_75t_L g4335 ( 
.A(n_4122),
.B(n_3844),
.Y(n_4335)
);

INVx1_ASAP7_75t_L g4336 ( 
.A(n_3997),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_3997),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_4005),
.Y(n_4338)
);

OR2x6_ASAP7_75t_L g4339 ( 
.A(n_4122),
.B(n_3873),
.Y(n_4339)
);

INVx1_ASAP7_75t_L g4340 ( 
.A(n_4005),
.Y(n_4340)
);

AND2x4_ASAP7_75t_L g4341 ( 
.A(n_4091),
.B(n_3878),
.Y(n_4341)
);

INVx2_ASAP7_75t_SL g4342 ( 
.A(n_4122),
.Y(n_4342)
);

OR2x2_ASAP7_75t_L g4343 ( 
.A(n_4023),
.B(n_3743),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4122),
.Y(n_4344)
);

NOR3xp33_ASAP7_75t_L g4345 ( 
.A(n_4024),
.B(n_3916),
.C(n_3873),
.Y(n_4345)
);

OAI33xp33_ASAP7_75t_L g4346 ( 
.A1(n_3985),
.A2(n_3883),
.A3(n_3925),
.B1(n_3838),
.B2(n_3921),
.B3(n_3914),
.Y(n_4346)
);

OAI221xp5_ASAP7_75t_L g4347 ( 
.A1(n_4081),
.A2(n_3916),
.B1(n_3873),
.B2(n_3675),
.C(n_3687),
.Y(n_4347)
);

NOR2x1_ASAP7_75t_SL g4348 ( 
.A(n_3959),
.B(n_3878),
.Y(n_4348)
);

OR2x2_ASAP7_75t_L g4349 ( 
.A(n_4023),
.B(n_3743),
.Y(n_4349)
);

NOR2xp33_ASAP7_75t_L g4350 ( 
.A(n_4100),
.B(n_3916),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4011),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_L g4352 ( 
.A(n_4100),
.B(n_3450),
.Y(n_4352)
);

AO21x2_ASAP7_75t_L g4353 ( 
.A1(n_4165),
.A2(n_3896),
.B(n_3887),
.Y(n_4353)
);

AOI22xp33_ASAP7_75t_L g4354 ( 
.A1(n_4130),
.A2(n_3675),
.B1(n_3687),
.B2(n_3769),
.Y(n_4354)
);

AO21x1_ASAP7_75t_SL g4355 ( 
.A1(n_3985),
.A2(n_4013),
.B(n_3983),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4011),
.Y(n_4356)
);

INVx1_ASAP7_75t_L g4357 ( 
.A(n_4026),
.Y(n_4357)
);

BUFx6f_ASAP7_75t_L g4358 ( 
.A(n_4142),
.Y(n_4358)
);

OR2x2_ASAP7_75t_L g4359 ( 
.A(n_4139),
.B(n_3891),
.Y(n_4359)
);

AOI221x1_ASAP7_75t_SL g4360 ( 
.A1(n_4013),
.A2(n_3793),
.B1(n_3798),
.B2(n_3921),
.C(n_3914),
.Y(n_4360)
);

AO21x2_ASAP7_75t_L g4361 ( 
.A1(n_4165),
.A2(n_3950),
.B(n_3948),
.Y(n_4361)
);

INVx2_ASAP7_75t_L g4362 ( 
.A(n_4165),
.Y(n_4362)
);

INVx2_ASAP7_75t_L g4363 ( 
.A(n_3959),
.Y(n_4363)
);

AOI22xp33_ASAP7_75t_L g4364 ( 
.A1(n_4130),
.A2(n_3769),
.B1(n_3916),
.B2(n_3902),
.Y(n_4364)
);

NAND2xp5_ASAP7_75t_L g4365 ( 
.A(n_4100),
.B(n_3450),
.Y(n_4365)
);

HB1xp67_ASAP7_75t_L g4366 ( 
.A(n_4026),
.Y(n_4366)
);

AND2x2_ASAP7_75t_L g4367 ( 
.A(n_4100),
.B(n_3473),
.Y(n_4367)
);

OAI22xp33_ASAP7_75t_L g4368 ( 
.A1(n_3941),
.A2(n_3618),
.B1(n_3572),
.B2(n_3552),
.Y(n_4368)
);

AOI21xp33_ASAP7_75t_L g4369 ( 
.A1(n_4132),
.A2(n_3887),
.B(n_3896),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4027),
.Y(n_4370)
);

NOR5xp2_ASAP7_75t_SL g4371 ( 
.A(n_4129),
.B(n_3501),
.C(n_3550),
.D(n_3592),
.E(n_3796),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4103),
.B(n_3477),
.Y(n_4372)
);

INVxp67_ASAP7_75t_L g4373 ( 
.A(n_3966),
.Y(n_4373)
);

OR2x2_ASAP7_75t_L g4374 ( 
.A(n_4139),
.B(n_3891),
.Y(n_4374)
);

OAI22xp5_ASAP7_75t_L g4375 ( 
.A1(n_4129),
.A2(n_3452),
.B1(n_3381),
.B2(n_3775),
.Y(n_4375)
);

AND2x6_ASAP7_75t_SL g4376 ( 
.A(n_4088),
.B(n_3381),
.Y(n_4376)
);

AOI22xp33_ASAP7_75t_L g4377 ( 
.A1(n_4132),
.A2(n_3769),
.B1(n_3902),
.B2(n_3910),
.Y(n_4377)
);

AOI222xp33_ASAP7_75t_L g4378 ( 
.A1(n_4150),
.A2(n_3775),
.B1(n_3712),
.B2(n_3718),
.C1(n_3723),
.C2(n_3904),
.Y(n_4378)
);

NOR2xp33_ASAP7_75t_L g4379 ( 
.A(n_4088),
.B(n_3887),
.Y(n_4379)
);

INVxp67_ASAP7_75t_L g4380 ( 
.A(n_4355),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4211),
.Y(n_4381)
);

AND2x2_ASAP7_75t_L g4382 ( 
.A(n_4192),
.B(n_4004),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_4208),
.B(n_4150),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4211),
.Y(n_4384)
);

OR2x2_ASAP7_75t_L g4385 ( 
.A(n_4281),
.B(n_4138),
.Y(n_4385)
);

INVx2_ASAP7_75t_L g4386 ( 
.A(n_4231),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4201),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_4172),
.B(n_4153),
.Y(n_4388)
);

NOR2xp33_ASAP7_75t_L g4389 ( 
.A(n_4187),
.B(n_4089),
.Y(n_4389)
);

OR2x2_ASAP7_75t_L g4390 ( 
.A(n_4363),
.B(n_4138),
.Y(n_4390)
);

INVx2_ASAP7_75t_L g4391 ( 
.A(n_4231),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_4278),
.Y(n_4392)
);

INVx1_ASAP7_75t_L g4393 ( 
.A(n_4201),
.Y(n_4393)
);

NAND2x1_ASAP7_75t_L g4394 ( 
.A(n_4171),
.B(n_3966),
.Y(n_4394)
);

HB1xp67_ASAP7_75t_L g4395 ( 
.A(n_4202),
.Y(n_4395)
);

OR2x2_ASAP7_75t_L g4396 ( 
.A(n_4363),
.B(n_4149),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4192),
.B(n_4004),
.Y(n_4397)
);

HB1xp67_ASAP7_75t_L g4398 ( 
.A(n_4249),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4207),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4287),
.B(n_4007),
.Y(n_4400)
);

OR2x2_ASAP7_75t_L g4401 ( 
.A(n_4257),
.B(n_4149),
.Y(n_4401)
);

AND2x2_ASAP7_75t_L g4402 ( 
.A(n_4287),
.B(n_4007),
.Y(n_4402)
);

AND2x4_ASAP7_75t_L g4403 ( 
.A(n_4171),
.B(n_4076),
.Y(n_4403)
);

AND2x2_ASAP7_75t_L g4404 ( 
.A(n_4259),
.B(n_4012),
.Y(n_4404)
);

NOR2xp67_ASAP7_75t_L g4405 ( 
.A(n_4190),
.B(n_4076),
.Y(n_4405)
);

AND2x2_ASAP7_75t_L g4406 ( 
.A(n_4178),
.B(n_4012),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4278),
.Y(n_4407)
);

AND2x2_ASAP7_75t_SL g4408 ( 
.A(n_4171),
.B(n_3952),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4207),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4235),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4341),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4235),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_4176),
.B(n_4153),
.Y(n_4413)
);

AND2x2_ASAP7_75t_L g4414 ( 
.A(n_4264),
.B(n_4014),
.Y(n_4414)
);

INVx1_ASAP7_75t_L g4415 ( 
.A(n_4238),
.Y(n_4415)
);

AND2x2_ASAP7_75t_L g4416 ( 
.A(n_4227),
.B(n_4014),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_4353),
.Y(n_4417)
);

OAI31xp33_ASAP7_75t_L g4418 ( 
.A1(n_4185),
.A2(n_3952),
.A3(n_3984),
.B(n_4129),
.Y(n_4418)
);

INVx2_ASAP7_75t_SL g4419 ( 
.A(n_4341),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4238),
.Y(n_4420)
);

HB1xp67_ASAP7_75t_L g4421 ( 
.A(n_4244),
.Y(n_4421)
);

INVx3_ASAP7_75t_L g4422 ( 
.A(n_4353),
.Y(n_4422)
);

AND2x2_ASAP7_75t_L g4423 ( 
.A(n_4269),
.B(n_4019),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4242),
.B(n_4019),
.Y(n_4424)
);

AND2x2_ASAP7_75t_L g4425 ( 
.A(n_4248),
.B(n_4089),
.Y(n_4425)
);

AND2x2_ASAP7_75t_L g4426 ( 
.A(n_4210),
.B(n_4103),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4253),
.Y(n_4427)
);

OR2x2_ASAP7_75t_L g4428 ( 
.A(n_4267),
.B(n_3963),
.Y(n_4428)
);

OR2x2_ASAP7_75t_L g4429 ( 
.A(n_4169),
.B(n_4174),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4251),
.B(n_4321),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4253),
.Y(n_4431)
);

OR2x2_ASAP7_75t_L g4432 ( 
.A(n_4188),
.B(n_3963),
.Y(n_4432)
);

NAND2x1p5_ASAP7_75t_L g4433 ( 
.A(n_4219),
.B(n_4142),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_4325),
.B(n_4110),
.Y(n_4434)
);

OR2x2_ASAP7_75t_L g4435 ( 
.A(n_4194),
.B(n_3983),
.Y(n_4435)
);

AND2x2_ASAP7_75t_L g4436 ( 
.A(n_4285),
.B(n_4110),
.Y(n_4436)
);

INVx2_ASAP7_75t_L g4437 ( 
.A(n_4316),
.Y(n_4437)
);

AND2x4_ASAP7_75t_L g4438 ( 
.A(n_4180),
.B(n_4076),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4316),
.Y(n_4439)
);

INVx2_ASAP7_75t_L g4440 ( 
.A(n_4284),
.Y(n_4440)
);

AND2x4_ASAP7_75t_L g4441 ( 
.A(n_4180),
.B(n_4104),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4366),
.Y(n_4442)
);

INVx2_ASAP7_75t_L g4443 ( 
.A(n_4243),
.Y(n_4443)
);

NAND2xp5_ASAP7_75t_L g4444 ( 
.A(n_4176),
.B(n_4161),
.Y(n_4444)
);

OR2x2_ASAP7_75t_L g4445 ( 
.A(n_4197),
.B(n_4115),
.Y(n_4445)
);

NAND2xp5_ASAP7_75t_L g4446 ( 
.A(n_4179),
.B(n_4161),
.Y(n_4446)
);

INVx2_ASAP7_75t_L g4447 ( 
.A(n_4243),
.Y(n_4447)
);

INVx1_ASAP7_75t_L g4448 ( 
.A(n_4366),
.Y(n_4448)
);

INVx2_ASAP7_75t_L g4449 ( 
.A(n_4243),
.Y(n_4449)
);

BUFx2_ASAP7_75t_L g4450 ( 
.A(n_4215),
.Y(n_4450)
);

AND2x2_ASAP7_75t_L g4451 ( 
.A(n_4305),
.B(n_4116),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4179),
.B(n_4163),
.Y(n_4452)
);

INVx1_ASAP7_75t_SL g4453 ( 
.A(n_4215),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_4167),
.B(n_4163),
.Y(n_4454)
);

INVx1_ASAP7_75t_L g4455 ( 
.A(n_4200),
.Y(n_4455)
);

NAND2xp5_ASAP7_75t_L g4456 ( 
.A(n_4167),
.B(n_4166),
.Y(n_4456)
);

NAND2xp5_ASAP7_75t_SL g4457 ( 
.A(n_4173),
.B(n_4199),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4324),
.B(n_4116),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4203),
.Y(n_4459)
);

AND2x2_ASAP7_75t_L g4460 ( 
.A(n_4367),
.B(n_4047),
.Y(n_4460)
);

INVx2_ASAP7_75t_L g4461 ( 
.A(n_4341),
.Y(n_4461)
);

HB1xp67_ASAP7_75t_L g4462 ( 
.A(n_4326),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4180),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_4177),
.B(n_4166),
.Y(n_4464)
);

INVx2_ASAP7_75t_L g4465 ( 
.A(n_4303),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_4177),
.B(n_4104),
.Y(n_4466)
);

OR2x2_ASAP7_75t_L g4467 ( 
.A(n_4204),
.B(n_4115),
.Y(n_4467)
);

AND2x2_ASAP7_75t_L g4468 ( 
.A(n_4372),
.B(n_4047),
.Y(n_4468)
);

AND2x2_ASAP7_75t_L g4469 ( 
.A(n_4280),
.B(n_4053),
.Y(n_4469)
);

INVx1_ASAP7_75t_L g4470 ( 
.A(n_4312),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_4280),
.B(n_4053),
.Y(n_4471)
);

AND2x2_ASAP7_75t_L g4472 ( 
.A(n_4232),
.B(n_4055),
.Y(n_4472)
);

HB1xp67_ASAP7_75t_L g4473 ( 
.A(n_4326),
.Y(n_4473)
);

INVx3_ASAP7_75t_L g4474 ( 
.A(n_4303),
.Y(n_4474)
);

INVxp67_ASAP7_75t_SL g4475 ( 
.A(n_4348),
.Y(n_4475)
);

AND2x2_ASAP7_75t_L g4476 ( 
.A(n_4232),
.B(n_4055),
.Y(n_4476)
);

AND2x2_ASAP7_75t_SL g4477 ( 
.A(n_4222),
.B(n_3952),
.Y(n_4477)
);

BUFx3_ASAP7_75t_L g4478 ( 
.A(n_4191),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_4362),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_4303),
.B(n_4104),
.Y(n_4480)
);

INVx1_ASAP7_75t_L g4481 ( 
.A(n_4362),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_4361),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4195),
.B(n_4073),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4361),
.Y(n_4484)
);

AND2x2_ASAP7_75t_L g4485 ( 
.A(n_4350),
.B(n_4073),
.Y(n_4485)
);

AND2x4_ASAP7_75t_L g4486 ( 
.A(n_4181),
.B(n_4142),
.Y(n_4486)
);

INVx1_ASAP7_75t_L g4487 ( 
.A(n_4214),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4216),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4209),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_L g4490 ( 
.A(n_4229),
.B(n_3998),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_L g4491 ( 
.A(n_4229),
.B(n_3998),
.Y(n_4491)
);

INVxp67_ASAP7_75t_SL g4492 ( 
.A(n_4191),
.Y(n_4492)
);

HB1xp67_ASAP7_75t_L g4493 ( 
.A(n_4335),
.Y(n_4493)
);

AND2x2_ASAP7_75t_L g4494 ( 
.A(n_4350),
.B(n_3967),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4237),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4218),
.B(n_3967),
.Y(n_4496)
);

BUFx2_ASAP7_75t_L g4497 ( 
.A(n_4376),
.Y(n_4497)
);

AND2x2_ASAP7_75t_L g4498 ( 
.A(n_4218),
.B(n_3967),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_4168),
.B(n_4081),
.Y(n_4499)
);

BUFx2_ASAP7_75t_L g4500 ( 
.A(n_4225),
.Y(n_4500)
);

INVx2_ASAP7_75t_L g4501 ( 
.A(n_4358),
.Y(n_4501)
);

AND2x2_ASAP7_75t_L g4502 ( 
.A(n_4298),
.B(n_3967),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4358),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4247),
.Y(n_4504)
);

INVx1_ASAP7_75t_L g4505 ( 
.A(n_4255),
.Y(n_4505)
);

AND2x2_ASAP7_75t_L g4506 ( 
.A(n_4298),
.B(n_3979),
.Y(n_4506)
);

AND2x2_ASAP7_75t_L g4507 ( 
.A(n_4301),
.B(n_3979),
.Y(n_4507)
);

AND2x2_ASAP7_75t_L g4508 ( 
.A(n_4301),
.B(n_3979),
.Y(n_4508)
);

OR2x2_ASAP7_75t_L g4509 ( 
.A(n_4272),
.B(n_4154),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4260),
.Y(n_4510)
);

AND2x2_ASAP7_75t_L g4511 ( 
.A(n_4302),
.B(n_3979),
.Y(n_4511)
);

BUFx2_ASAP7_75t_L g4512 ( 
.A(n_4225),
.Y(n_4512)
);

INVx1_ASAP7_75t_L g4513 ( 
.A(n_4276),
.Y(n_4513)
);

OR2x2_ASAP7_75t_L g4514 ( 
.A(n_4250),
.B(n_4154),
.Y(n_4514)
);

INVx2_ASAP7_75t_L g4515 ( 
.A(n_4358),
.Y(n_4515)
);

AND2x2_ASAP7_75t_L g4516 ( 
.A(n_4302),
.B(n_3984),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4279),
.Y(n_4517)
);

OR2x2_ASAP7_75t_L g4518 ( 
.A(n_4373),
.B(n_4098),
.Y(n_4518)
);

AND2x2_ASAP7_75t_L g4519 ( 
.A(n_4307),
.B(n_3984),
.Y(n_4519)
);

AND2x2_ASAP7_75t_L g4520 ( 
.A(n_4175),
.B(n_4084),
.Y(n_4520)
);

NAND2x1_ASAP7_75t_L g4521 ( 
.A(n_4335),
.B(n_4157),
.Y(n_4521)
);

NOR2x1_ASAP7_75t_L g4522 ( 
.A(n_4219),
.B(n_3941),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_4234),
.B(n_4084),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_4189),
.B(n_4098),
.Y(n_4524)
);

OR2x2_ASAP7_75t_L g4525 ( 
.A(n_4359),
.B(n_4027),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4283),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4360),
.B(n_4048),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4175),
.B(n_4099),
.Y(n_4528)
);

INVx2_ASAP7_75t_L g4529 ( 
.A(n_4209),
.Y(n_4529)
);

AND2x4_ASAP7_75t_SL g4530 ( 
.A(n_4175),
.B(n_4256),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_L g4531 ( 
.A(n_4299),
.B(n_4048),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4261),
.B(n_4099),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4209),
.Y(n_4533)
);

AND2x2_ASAP7_75t_L g4534 ( 
.A(n_4261),
.B(n_4099),
.Y(n_4534)
);

INVx2_ASAP7_75t_L g4535 ( 
.A(n_4358),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4304),
.B(n_4048),
.Y(n_4536)
);

AND2x2_ASAP7_75t_L g4537 ( 
.A(n_4193),
.B(n_4114),
.Y(n_4537)
);

INVx2_ASAP7_75t_L g4538 ( 
.A(n_4241),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_4317),
.B(n_4048),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4193),
.B(n_4114),
.Y(n_4540)
);

AND2x2_ASAP7_75t_L g4541 ( 
.A(n_4193),
.B(n_4256),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4288),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_4291),
.Y(n_4543)
);

INVx5_ASAP7_75t_L g4544 ( 
.A(n_4256),
.Y(n_4544)
);

BUFx2_ASAP7_75t_L g4545 ( 
.A(n_4181),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4292),
.Y(n_4546)
);

OAI21xp5_ASAP7_75t_SL g4547 ( 
.A1(n_4213),
.A2(n_4049),
.B(n_4157),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4319),
.Y(n_4548)
);

INVx1_ASAP7_75t_L g4549 ( 
.A(n_4323),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4265),
.B(n_4114),
.Y(n_4550)
);

OR2x2_ASAP7_75t_L g4551 ( 
.A(n_4374),
.B(n_4031),
.Y(n_4551)
);

OR2x2_ASAP7_75t_L g4552 ( 
.A(n_4294),
.B(n_4031),
.Y(n_4552)
);

AND2x2_ASAP7_75t_L g4553 ( 
.A(n_4378),
.B(n_4114),
.Y(n_4553)
);

AND2x4_ASAP7_75t_L g4554 ( 
.A(n_4335),
.B(n_4157),
.Y(n_4554)
);

INVx1_ASAP7_75t_L g4555 ( 
.A(n_4333),
.Y(n_4555)
);

AND2x2_ASAP7_75t_L g4556 ( 
.A(n_4297),
.B(n_4126),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4186),
.B(n_4049),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4379),
.B(n_4126),
.Y(n_4558)
);

BUFx2_ASAP7_75t_L g4559 ( 
.A(n_4339),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_4198),
.B(n_4049),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4339),
.B(n_4157),
.Y(n_4561)
);

NOR2xp33_ASAP7_75t_L g4562 ( 
.A(n_4223),
.B(n_4126),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_4339),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4379),
.B(n_4126),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4352),
.B(n_4049),
.Y(n_4565)
);

INVx1_ASAP7_75t_L g4566 ( 
.A(n_4431),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_4492),
.B(n_4342),
.Y(n_4567)
);

AND2x2_ASAP7_75t_L g4568 ( 
.A(n_4434),
.B(n_4450),
.Y(n_4568)
);

INVxp67_ASAP7_75t_L g4569 ( 
.A(n_4450),
.Y(n_4569)
);

INVx1_ASAP7_75t_L g4570 ( 
.A(n_4431),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_4478),
.B(n_4233),
.Y(n_4571)
);

INVx1_ASAP7_75t_L g4572 ( 
.A(n_4431),
.Y(n_4572)
);

OR2x2_ASAP7_75t_L g4573 ( 
.A(n_4385),
.B(n_4490),
.Y(n_4573)
);

AND2x4_ASAP7_75t_L g4574 ( 
.A(n_4438),
.B(n_4183),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4437),
.Y(n_4575)
);

AND2x4_ASAP7_75t_L g4576 ( 
.A(n_4438),
.B(n_4183),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_L g4577 ( 
.A(n_4478),
.B(n_4365),
.Y(n_4577)
);

NAND2x1p5_ASAP7_75t_L g4578 ( 
.A(n_4544),
.B(n_4184),
.Y(n_4578)
);

INVx1_ASAP7_75t_L g4579 ( 
.A(n_4437),
.Y(n_4579)
);

OR2x2_ASAP7_75t_L g4580 ( 
.A(n_4385),
.B(n_4327),
.Y(n_4580)
);

INVx1_ASAP7_75t_L g4581 ( 
.A(n_4437),
.Y(n_4581)
);

AND2x2_ASAP7_75t_L g4582 ( 
.A(n_4434),
.B(n_4478),
.Y(n_4582)
);

INVx3_ASAP7_75t_SL g4583 ( 
.A(n_4408),
.Y(n_4583)
);

CKINVDCx16_ASAP7_75t_R g4584 ( 
.A(n_4453),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_4489),
.Y(n_4585)
);

OR2x2_ASAP7_75t_L g4586 ( 
.A(n_4491),
.B(n_4274),
.Y(n_4586)
);

OR2x2_ASAP7_75t_L g4587 ( 
.A(n_4395),
.B(n_4282),
.Y(n_4587)
);

AOI21x1_ASAP7_75t_SL g4588 ( 
.A1(n_4556),
.A2(n_4094),
.B(n_4090),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4414),
.B(n_4289),
.Y(n_4589)
);

INVx2_ASAP7_75t_L g4590 ( 
.A(n_4545),
.Y(n_4590)
);

INVx1_ASAP7_75t_L g4591 ( 
.A(n_4439),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4414),
.B(n_4262),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_4398),
.B(n_4310),
.Y(n_4593)
);

AND2x2_ASAP7_75t_L g4594 ( 
.A(n_4423),
.B(n_4254),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4439),
.Y(n_4595)
);

INVx1_ASAP7_75t_L g4596 ( 
.A(n_4439),
.Y(n_4596)
);

INVx2_ASAP7_75t_L g4597 ( 
.A(n_4545),
.Y(n_4597)
);

AND2x2_ASAP7_75t_L g4598 ( 
.A(n_4423),
.B(n_4404),
.Y(n_4598)
);

OR2x2_ASAP7_75t_L g4599 ( 
.A(n_4401),
.B(n_4343),
.Y(n_4599)
);

OR2x2_ASAP7_75t_L g4600 ( 
.A(n_4401),
.B(n_4349),
.Y(n_4600)
);

AND2x2_ASAP7_75t_L g4601 ( 
.A(n_4404),
.B(n_4311),
.Y(n_4601)
);

BUFx2_ASAP7_75t_L g4602 ( 
.A(n_4403),
.Y(n_4602)
);

INVx2_ASAP7_75t_L g4603 ( 
.A(n_4438),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4509),
.B(n_4170),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4381),
.B(n_4310),
.Y(n_4605)
);

OR2x2_ASAP7_75t_L g4606 ( 
.A(n_4509),
.B(n_4206),
.Y(n_4606)
);

OR2x2_ASAP7_75t_L g4607 ( 
.A(n_4381),
.B(n_4384),
.Y(n_4607)
);

AND2x4_ASAP7_75t_L g4608 ( 
.A(n_4438),
.B(n_4184),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4451),
.B(n_4311),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4462),
.Y(n_4610)
);

INVxp67_ASAP7_75t_SL g4611 ( 
.A(n_4394),
.Y(n_4611)
);

OAI21xp33_ASAP7_75t_L g4612 ( 
.A1(n_4499),
.A2(n_4205),
.B(n_4196),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4384),
.B(n_4182),
.Y(n_4613)
);

AND2x2_ASAP7_75t_L g4614 ( 
.A(n_4451),
.B(n_4145),
.Y(n_4614)
);

AND2x4_ASAP7_75t_SL g4615 ( 
.A(n_4403),
.B(n_4145),
.Y(n_4615)
);

BUFx3_ASAP7_75t_L g4616 ( 
.A(n_4386),
.Y(n_4616)
);

AND2x2_ASAP7_75t_L g4617 ( 
.A(n_4382),
.B(n_4145),
.Y(n_4617)
);

OR2x2_ASAP7_75t_L g4618 ( 
.A(n_4386),
.B(n_4318),
.Y(n_4618)
);

BUFx2_ASAP7_75t_L g4619 ( 
.A(n_4403),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4473),
.Y(n_4620)
);

OR2x2_ASAP7_75t_L g4621 ( 
.A(n_4470),
.B(n_4429),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4382),
.B(n_4145),
.Y(n_4622)
);

INVx2_ASAP7_75t_L g4623 ( 
.A(n_4441),
.Y(n_4623)
);

NAND2xp67_ASAP7_75t_L g4624 ( 
.A(n_4391),
.B(n_4217),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4397),
.B(n_4158),
.Y(n_4625)
);

INVx2_ASAP7_75t_L g4626 ( 
.A(n_4441),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_4387),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4387),
.Y(n_4628)
);

NAND2xp5_ASAP7_75t_L g4629 ( 
.A(n_4391),
.B(n_4258),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4392),
.B(n_4236),
.Y(n_4630)
);

AND2x2_ASAP7_75t_L g4631 ( 
.A(n_4397),
.B(n_4158),
.Y(n_4631)
);

OR2x2_ASAP7_75t_L g4632 ( 
.A(n_4470),
.B(n_4217),
.Y(n_4632)
);

NAND2xp5_ASAP7_75t_L g4633 ( 
.A(n_4392),
.B(n_4271),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4400),
.B(n_4158),
.Y(n_4634)
);

INVx2_ASAP7_75t_L g4635 ( 
.A(n_4441),
.Y(n_4635)
);

AND2x2_ASAP7_75t_L g4636 ( 
.A(n_4400),
.B(n_4402),
.Y(n_4636)
);

OR2x2_ASAP7_75t_L g4637 ( 
.A(n_4407),
.B(n_4263),
.Y(n_4637)
);

NAND2xp5_ASAP7_75t_L g4638 ( 
.A(n_4407),
.B(n_4271),
.Y(n_4638)
);

AND2x2_ASAP7_75t_L g4639 ( 
.A(n_4402),
.B(n_4158),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4472),
.B(n_4314),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4393),
.Y(n_4641)
);

INVx1_ASAP7_75t_SL g4642 ( 
.A(n_4408),
.Y(n_4642)
);

AND2x2_ASAP7_75t_L g4643 ( 
.A(n_4472),
.B(n_4314),
.Y(n_4643)
);

AND2x2_ASAP7_75t_L g4644 ( 
.A(n_4476),
.B(n_4375),
.Y(n_4644)
);

INVx1_ASAP7_75t_L g4645 ( 
.A(n_4393),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4399),
.Y(n_4646)
);

INVx1_ASAP7_75t_L g4647 ( 
.A(n_4399),
.Y(n_4647)
);

AND2x2_ASAP7_75t_SL g4648 ( 
.A(n_4477),
.B(n_4222),
.Y(n_4648)
);

NAND2xp5_ASAP7_75t_L g4649 ( 
.A(n_4405),
.B(n_4430),
.Y(n_4649)
);

INVx1_ASAP7_75t_L g4650 ( 
.A(n_4409),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4409),
.Y(n_4651)
);

OR2x2_ASAP7_75t_L g4652 ( 
.A(n_4514),
.B(n_4277),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4405),
.B(n_4277),
.Y(n_4653)
);

NOR2xp67_ASAP7_75t_L g4654 ( 
.A(n_4544),
.B(n_4230),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_4430),
.B(n_4290),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4476),
.B(n_4090),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4410),
.Y(n_4657)
);

INVx1_ASAP7_75t_L g4658 ( 
.A(n_4410),
.Y(n_4658)
);

OR2x2_ASAP7_75t_L g4659 ( 
.A(n_4429),
.B(n_4290),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4408),
.B(n_4094),
.Y(n_4660)
);

OR2x2_ASAP7_75t_L g4661 ( 
.A(n_4514),
.B(n_4306),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4441),
.Y(n_4662)
);

INVx2_ASAP7_75t_L g4663 ( 
.A(n_4403),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_L g4664 ( 
.A(n_4477),
.B(n_4306),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4433),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4477),
.B(n_4309),
.Y(n_4666)
);

HB1xp67_ASAP7_75t_L g4667 ( 
.A(n_4489),
.Y(n_4667)
);

NOR2xp33_ASAP7_75t_L g4668 ( 
.A(n_4500),
.B(n_4275),
.Y(n_4668)
);

INVxp67_ASAP7_75t_SL g4669 ( 
.A(n_4394),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4412),
.Y(n_4670)
);

AND2x4_ASAP7_75t_L g4671 ( 
.A(n_4544),
.B(n_4309),
.Y(n_4671)
);

AND2x2_ASAP7_75t_L g4672 ( 
.A(n_4406),
.B(n_4095),
.Y(n_4672)
);

OR2x2_ASAP7_75t_L g4673 ( 
.A(n_4523),
.B(n_4320),
.Y(n_4673)
);

AND2x4_ASAP7_75t_SL g4674 ( 
.A(n_4496),
.B(n_4320),
.Y(n_4674)
);

NOR2xp67_ASAP7_75t_L g4675 ( 
.A(n_4544),
.B(n_4224),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4497),
.B(n_4329),
.Y(n_4676)
);

OR2x2_ASAP7_75t_L g4677 ( 
.A(n_4390),
.B(n_4329),
.Y(n_4677)
);

INVx3_ASAP7_75t_L g4678 ( 
.A(n_4480),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_4406),
.B(n_4095),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4433),
.Y(n_4680)
);

INVx1_ASAP7_75t_L g4681 ( 
.A(n_4412),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4497),
.B(n_4330),
.Y(n_4682)
);

HB1xp67_ASAP7_75t_L g4683 ( 
.A(n_4489),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4436),
.B(n_4330),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4415),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_4519),
.B(n_4344),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4519),
.B(n_4344),
.Y(n_4687)
);

INVxp67_ASAP7_75t_L g4688 ( 
.A(n_4389),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4390),
.B(n_4239),
.Y(n_4689)
);

AND2x2_ASAP7_75t_L g4690 ( 
.A(n_4436),
.B(n_4345),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_4500),
.B(n_4212),
.Y(n_4691)
);

INVx1_ASAP7_75t_L g4692 ( 
.A(n_4415),
.Y(n_4692)
);

OR2x2_ASAP7_75t_L g4693 ( 
.A(n_4428),
.B(n_4228),
.Y(n_4693)
);

OR2x2_ASAP7_75t_L g4694 ( 
.A(n_4396),
.B(n_4336),
.Y(n_4694)
);

INVx1_ASAP7_75t_L g4695 ( 
.A(n_4420),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4420),
.Y(n_4696)
);

OR2x2_ASAP7_75t_L g4697 ( 
.A(n_4428),
.B(n_4226),
.Y(n_4697)
);

NOR2xp67_ASAP7_75t_L g4698 ( 
.A(n_4544),
.B(n_4295),
.Y(n_4698)
);

NOR2xp33_ASAP7_75t_L g4699 ( 
.A(n_4512),
.B(n_4322),
.Y(n_4699)
);

BUFx2_ASAP7_75t_L g4700 ( 
.A(n_4480),
.Y(n_4700)
);

INVx1_ASAP7_75t_SL g4701 ( 
.A(n_4512),
.Y(n_4701)
);

OR2x2_ASAP7_75t_L g4702 ( 
.A(n_4383),
.B(n_4240),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4427),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4380),
.B(n_4337),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4416),
.B(n_4245),
.Y(n_4705)
);

BUFx2_ASAP7_75t_L g4706 ( 
.A(n_4480),
.Y(n_4706)
);

AND2x2_ASAP7_75t_L g4707 ( 
.A(n_4416),
.B(n_4245),
.Y(n_4707)
);

OR2x2_ASAP7_75t_L g4708 ( 
.A(n_4396),
.B(n_4338),
.Y(n_4708)
);

INVx1_ASAP7_75t_L g4709 ( 
.A(n_4427),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4442),
.Y(n_4710)
);

INVx2_ASAP7_75t_L g4711 ( 
.A(n_4433),
.Y(n_4711)
);

AND2x2_ASAP7_75t_L g4712 ( 
.A(n_4426),
.B(n_4246),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4529),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4529),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_4418),
.B(n_4340),
.Y(n_4715)
);

OR2x2_ASAP7_75t_L g4716 ( 
.A(n_4483),
.B(n_4266),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4442),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4426),
.B(n_4246),
.Y(n_4718)
);

NAND2x1_ASAP7_75t_L g4719 ( 
.A(n_4554),
.B(n_4334),
.Y(n_4719)
);

AND2x2_ASAP7_75t_L g4720 ( 
.A(n_4424),
.B(n_4220),
.Y(n_4720)
);

INVx1_ASAP7_75t_L g4721 ( 
.A(n_4448),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4448),
.Y(n_4722)
);

INVx2_ASAP7_75t_L g4723 ( 
.A(n_4529),
.Y(n_4723)
);

INVx4_ASAP7_75t_L g4724 ( 
.A(n_4544),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4482),
.Y(n_4725)
);

INVx3_ASAP7_75t_L g4726 ( 
.A(n_4480),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4582),
.B(n_4501),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4585),
.Y(n_4728)
);

NOR2xp67_ASAP7_75t_SL g4729 ( 
.A(n_4584),
.B(n_4493),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_L g4730 ( 
.A(n_4582),
.B(n_4501),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4585),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4678),
.Y(n_4732)
);

INVx1_ASAP7_75t_L g4733 ( 
.A(n_4667),
.Y(n_4733)
);

OR2x2_ASAP7_75t_L g4734 ( 
.A(n_4701),
.B(n_4466),
.Y(n_4734)
);

INVx1_ASAP7_75t_L g4735 ( 
.A(n_4667),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4678),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4568),
.B(n_4460),
.Y(n_4737)
);

INVx2_ASAP7_75t_L g4738 ( 
.A(n_4678),
.Y(n_4738)
);

AND2x2_ASAP7_75t_L g4739 ( 
.A(n_4568),
.B(n_4496),
.Y(n_4739)
);

OAI21xp33_ASAP7_75t_L g4740 ( 
.A1(n_4612),
.A2(n_4457),
.B(n_4547),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4598),
.B(n_4503),
.Y(n_4741)
);

INVx1_ASAP7_75t_L g4742 ( 
.A(n_4683),
.Y(n_4742)
);

INVx2_ASAP7_75t_L g4743 ( 
.A(n_4726),
.Y(n_4743)
);

INVx1_ASAP7_75t_L g4744 ( 
.A(n_4683),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4598),
.B(n_4503),
.Y(n_4745)
);

AND2x4_ASAP7_75t_L g4746 ( 
.A(n_4726),
.B(n_4463),
.Y(n_4746)
);

OR2x2_ASAP7_75t_L g4747 ( 
.A(n_4587),
.B(n_4524),
.Y(n_4747)
);

NOR2xp67_ASAP7_75t_L g4748 ( 
.A(n_4726),
.B(n_4421),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4590),
.Y(n_4749)
);

OR2x2_ASAP7_75t_L g4750 ( 
.A(n_4587),
.B(n_4580),
.Y(n_4750)
);

INVx1_ASAP7_75t_L g4751 ( 
.A(n_4590),
.Y(n_4751)
);

NAND2x1p5_ASAP7_75t_L g4752 ( 
.A(n_4724),
.B(n_4521),
.Y(n_4752)
);

OAI21xp33_ASAP7_75t_SL g4753 ( 
.A1(n_4648),
.A2(n_4418),
.B(n_4556),
.Y(n_4753)
);

BUFx3_ASAP7_75t_L g4754 ( 
.A(n_4602),
.Y(n_4754)
);

INVx2_ASAP7_75t_L g4755 ( 
.A(n_4619),
.Y(n_4755)
);

NAND2xp5_ASAP7_75t_L g4756 ( 
.A(n_4648),
.B(n_4515),
.Y(n_4756)
);

AND2x2_ASAP7_75t_L g4757 ( 
.A(n_4636),
.B(n_4460),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_L g4758 ( 
.A(n_4616),
.B(n_4515),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4597),
.Y(n_4759)
);

NOR2xp33_ASAP7_75t_L g4760 ( 
.A(n_4583),
.B(n_4547),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4615),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4636),
.B(n_4458),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4609),
.B(n_4458),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4597),
.Y(n_4764)
);

INVx1_ASAP7_75t_L g4765 ( 
.A(n_4700),
.Y(n_4765)
);

AND2x4_ASAP7_75t_L g4766 ( 
.A(n_4706),
.B(n_4463),
.Y(n_4766)
);

AND2x2_ASAP7_75t_L g4767 ( 
.A(n_4609),
.B(n_4424),
.Y(n_4767)
);

NAND2xp5_ASAP7_75t_L g4768 ( 
.A(n_4616),
.B(n_4684),
.Y(n_4768)
);

HB1xp67_ASAP7_75t_L g4769 ( 
.A(n_4624),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4615),
.Y(n_4770)
);

OA21x2_ASAP7_75t_L g4771 ( 
.A1(n_4691),
.A2(n_4533),
.B(n_4447),
.Y(n_4771)
);

OAI21xp33_ASAP7_75t_L g4772 ( 
.A1(n_4668),
.A2(n_4562),
.B(n_4557),
.Y(n_4772)
);

INVx1_ASAP7_75t_SL g4773 ( 
.A(n_4583),
.Y(n_4773)
);

INVx1_ASAP7_75t_L g4774 ( 
.A(n_4621),
.Y(n_4774)
);

INVx2_ASAP7_75t_SL g4775 ( 
.A(n_4674),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4621),
.Y(n_4776)
);

INVx2_ASAP7_75t_L g4777 ( 
.A(n_4578),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4677),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4644),
.B(n_4498),
.Y(n_4779)
);

OR2x2_ASAP7_75t_L g4780 ( 
.A(n_4607),
.B(n_4445),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4677),
.Y(n_4781)
);

OR2x2_ASAP7_75t_L g4782 ( 
.A(n_4689),
.B(n_4445),
.Y(n_4782)
);

AND2x2_ASAP7_75t_L g4783 ( 
.A(n_4614),
.B(n_4425),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4684),
.B(n_4535),
.Y(n_4784)
);

AND2x2_ASAP7_75t_L g4785 ( 
.A(n_4614),
.B(n_4425),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4663),
.B(n_4535),
.Y(n_4786)
);

INVx1_ASAP7_75t_L g4787 ( 
.A(n_4713),
.Y(n_4787)
);

NAND2xp5_ASAP7_75t_L g4788 ( 
.A(n_4663),
.B(n_4532),
.Y(n_4788)
);

NAND2x1p5_ASAP7_75t_L g4789 ( 
.A(n_4724),
.B(n_4521),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4713),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4714),
.Y(n_4791)
);

INVx1_ASAP7_75t_SL g4792 ( 
.A(n_4674),
.Y(n_4792)
);

NAND2xp5_ASAP7_75t_L g4793 ( 
.A(n_4569),
.B(n_4532),
.Y(n_4793)
);

INVx1_ASAP7_75t_SL g4794 ( 
.A(n_4599),
.Y(n_4794)
);

AND2x2_ASAP7_75t_L g4795 ( 
.A(n_4644),
.B(n_4468),
.Y(n_4795)
);

OR2x2_ASAP7_75t_L g4796 ( 
.A(n_4689),
.B(n_4467),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4714),
.Y(n_4797)
);

HB1xp67_ASAP7_75t_L g4798 ( 
.A(n_4603),
.Y(n_4798)
);

INVx1_ASAP7_75t_L g4799 ( 
.A(n_4723),
.Y(n_4799)
);

INVx1_ASAP7_75t_L g4800 ( 
.A(n_4723),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4672),
.B(n_4468),
.Y(n_4801)
);

OR2x2_ASAP7_75t_L g4802 ( 
.A(n_4686),
.B(n_4687),
.Y(n_4802)
);

NOR2x1_ASAP7_75t_L g4803 ( 
.A(n_4724),
.B(n_4559),
.Y(n_4803)
);

AND2x4_ASAP7_75t_L g4804 ( 
.A(n_4574),
.B(n_4486),
.Y(n_4804)
);

AND2x2_ASAP7_75t_L g4805 ( 
.A(n_4672),
.B(n_4498),
.Y(n_4805)
);

AND2x2_ASAP7_75t_L g4806 ( 
.A(n_4679),
.B(n_4534),
.Y(n_4806)
);

NAND2x1_ASAP7_75t_L g4807 ( 
.A(n_4574),
.B(n_4559),
.Y(n_4807)
);

OR2x2_ASAP7_75t_L g4808 ( 
.A(n_4652),
.B(n_4467),
.Y(n_4808)
);

OAI22xp5_ASAP7_75t_L g4809 ( 
.A1(n_4613),
.A2(n_4199),
.B1(n_4221),
.B2(n_4293),
.Y(n_4809)
);

AND2x2_ASAP7_75t_L g4810 ( 
.A(n_4679),
.B(n_4494),
.Y(n_4810)
);

INVxp67_ASAP7_75t_L g4811 ( 
.A(n_4611),
.Y(n_4811)
);

AND2x2_ASAP7_75t_L g4812 ( 
.A(n_4656),
.B(n_4494),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4656),
.B(n_4485),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_L g4814 ( 
.A(n_4642),
.B(n_4534),
.Y(n_4814)
);

OR2x2_ASAP7_75t_L g4815 ( 
.A(n_4661),
.B(n_4432),
.Y(n_4815)
);

NAND2x1p5_ASAP7_75t_L g4816 ( 
.A(n_4654),
.B(n_4541),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4617),
.B(n_4622),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4720),
.B(n_4553),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_4659),
.Y(n_4819)
);

OR2x2_ASAP7_75t_L g4820 ( 
.A(n_4655),
.B(n_4432),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4720),
.B(n_4553),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4659),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4566),
.Y(n_4823)
);

INVx2_ASAP7_75t_L g4824 ( 
.A(n_4578),
.Y(n_4824)
);

HB1xp67_ASAP7_75t_L g4825 ( 
.A(n_4603),
.Y(n_4825)
);

AND2x2_ASAP7_75t_L g4826 ( 
.A(n_4617),
.B(n_4485),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4705),
.B(n_4707),
.Y(n_4827)
);

AOI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_4668),
.A2(n_4296),
.B1(n_4471),
.B2(n_4469),
.Y(n_4828)
);

AND2x2_ASAP7_75t_L g4829 ( 
.A(n_4622),
.B(n_4502),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4570),
.Y(n_4830)
);

OR2x2_ASAP7_75t_L g4831 ( 
.A(n_4600),
.B(n_4435),
.Y(n_4831)
);

INVx1_ASAP7_75t_L g4832 ( 
.A(n_4572),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4575),
.Y(n_4833)
);

HB1xp67_ASAP7_75t_L g4834 ( 
.A(n_4623),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4705),
.B(n_4537),
.Y(n_4835)
);

INVx1_ASAP7_75t_L g4836 ( 
.A(n_4579),
.Y(n_4836)
);

AND2x2_ASAP7_75t_L g4837 ( 
.A(n_4625),
.B(n_4502),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_L g4838 ( 
.A(n_4707),
.B(n_4537),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4577),
.B(n_4567),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4581),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4625),
.B(n_4506),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4631),
.B(n_4506),
.Y(n_4842)
);

NAND2xp5_ASAP7_75t_L g4843 ( 
.A(n_4712),
.B(n_4540),
.Y(n_4843)
);

HB1xp67_ASAP7_75t_L g4844 ( 
.A(n_4623),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4591),
.Y(n_4845)
);

INVx1_ASAP7_75t_SL g4846 ( 
.A(n_4649),
.Y(n_4846)
);

INVx2_ASAP7_75t_SL g4847 ( 
.A(n_4574),
.Y(n_4847)
);

AND2x2_ASAP7_75t_L g4848 ( 
.A(n_4631),
.B(n_4507),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4595),
.Y(n_4849)
);

HB1xp67_ASAP7_75t_L g4850 ( 
.A(n_4626),
.Y(n_4850)
);

OAI21xp5_ASAP7_75t_L g4851 ( 
.A1(n_4699),
.A2(n_4541),
.B(n_4540),
.Y(n_4851)
);

INVx1_ASAP7_75t_L g4852 ( 
.A(n_4596),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4626),
.Y(n_4853)
);

AND2x2_ASAP7_75t_L g4854 ( 
.A(n_4634),
.B(n_4507),
.Y(n_4854)
);

AND2x4_ASAP7_75t_L g4855 ( 
.A(n_4576),
.B(n_4486),
.Y(n_4855)
);

INVx2_ASAP7_75t_L g4856 ( 
.A(n_4576),
.Y(n_4856)
);

AOI22xp5_ASAP7_75t_L g4857 ( 
.A1(n_4699),
.A2(n_4296),
.B1(n_4471),
.B2(n_4469),
.Y(n_4857)
);

NAND2xp5_ASAP7_75t_L g4858 ( 
.A(n_4712),
.B(n_4508),
.Y(n_4858)
);

OR2x2_ASAP7_75t_L g4859 ( 
.A(n_4676),
.B(n_4435),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4635),
.Y(n_4860)
);

NAND4xp25_ASAP7_75t_L g4861 ( 
.A(n_4601),
.B(n_4516),
.C(n_4511),
.D(n_4508),
.Y(n_4861)
);

OAI21xp33_ASAP7_75t_L g4862 ( 
.A1(n_4629),
.A2(n_4516),
.B(n_4511),
.Y(n_4862)
);

INVx1_ASAP7_75t_SL g4863 ( 
.A(n_4634),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4635),
.Y(n_4864)
);

INVx2_ASAP7_75t_L g4865 ( 
.A(n_4576),
.Y(n_4865)
);

AND2x2_ASAP7_75t_L g4866 ( 
.A(n_4639),
.B(n_4520),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4718),
.B(n_4662),
.Y(n_4867)
);

OR2x2_ASAP7_75t_L g4868 ( 
.A(n_4750),
.B(n_4682),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4798),
.Y(n_4869)
);

INVx2_ASAP7_75t_SL g4870 ( 
.A(n_4804),
.Y(n_4870)
);

INVx1_ASAP7_75t_SL g4871 ( 
.A(n_4737),
.Y(n_4871)
);

INVxp67_ASAP7_75t_L g4872 ( 
.A(n_4729),
.Y(n_4872)
);

INVx1_ASAP7_75t_L g4873 ( 
.A(n_4798),
.Y(n_4873)
);

INVx1_ASAP7_75t_L g4874 ( 
.A(n_4825),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_4825),
.Y(n_4875)
);

AOI22xp5_ASAP7_75t_SL g4876 ( 
.A1(n_4809),
.A2(n_4669),
.B1(n_4737),
.B2(n_4754),
.Y(n_4876)
);

INVx1_ASAP7_75t_SL g4877 ( 
.A(n_4739),
.Y(n_4877)
);

OAI33xp33_ASAP7_75t_L g4878 ( 
.A1(n_4740),
.A2(n_4593),
.A3(n_4605),
.B1(n_4630),
.B2(n_4715),
.B3(n_4573),
.Y(n_4878)
);

OAI21xp33_ASAP7_75t_L g4879 ( 
.A1(n_4772),
.A2(n_4857),
.B(n_4827),
.Y(n_4879)
);

OR2x2_ASAP7_75t_L g4880 ( 
.A(n_4858),
.B(n_4604),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4834),
.Y(n_4881)
);

INVx2_ASAP7_75t_L g4882 ( 
.A(n_4804),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4834),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4754),
.B(n_4610),
.Y(n_4884)
);

OAI322xp33_ASAP7_75t_L g4885 ( 
.A1(n_4828),
.A2(n_4693),
.A3(n_4697),
.B1(n_4527),
.B2(n_4606),
.C1(n_4586),
.C2(n_4702),
.Y(n_4885)
);

OR2x2_ASAP7_75t_L g4886 ( 
.A(n_4867),
.B(n_4704),
.Y(n_4886)
);

INVx2_ASAP7_75t_L g4887 ( 
.A(n_4804),
.Y(n_4887)
);

BUFx2_ASAP7_75t_SL g4888 ( 
.A(n_4748),
.Y(n_4888)
);

INVx1_ASAP7_75t_SL g4889 ( 
.A(n_4855),
.Y(n_4889)
);

INVx1_ASAP7_75t_L g4890 ( 
.A(n_4844),
.Y(n_4890)
);

AND2x4_ASAP7_75t_L g4891 ( 
.A(n_4855),
.B(n_4662),
.Y(n_4891)
);

AOI22x1_ASAP7_75t_L g4892 ( 
.A1(n_4816),
.A2(n_4475),
.B1(n_4601),
.B2(n_4640),
.Y(n_4892)
);

AND2x2_ASAP7_75t_L g4893 ( 
.A(n_4795),
.B(n_4640),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4795),
.B(n_4589),
.Y(n_4894)
);

INVx1_ASAP7_75t_SL g4895 ( 
.A(n_4855),
.Y(n_4895)
);

AND2x2_ASAP7_75t_L g4896 ( 
.A(n_4757),
.B(n_4643),
.Y(n_4896)
);

AOI22xp5_ASAP7_75t_L g4897 ( 
.A1(n_4753),
.A2(n_4718),
.B1(n_4643),
.B2(n_4592),
.Y(n_4897)
);

AND2x2_ASAP7_75t_L g4898 ( 
.A(n_4757),
.B(n_4660),
.Y(n_4898)
);

AND2x2_ASAP7_75t_L g4899 ( 
.A(n_4762),
.B(n_4660),
.Y(n_4899)
);

AOI211xp5_ASAP7_75t_L g4900 ( 
.A1(n_4851),
.A2(n_4675),
.B(n_4698),
.C(n_4571),
.Y(n_4900)
);

INVx1_ASAP7_75t_L g4901 ( 
.A(n_4844),
.Y(n_4901)
);

INVx2_ASAP7_75t_L g4902 ( 
.A(n_4752),
.Y(n_4902)
);

INVx1_ASAP7_75t_L g4903 ( 
.A(n_4850),
.Y(n_4903)
);

A2O1A1Ixp33_ASAP7_75t_L g4904 ( 
.A1(n_4760),
.A2(n_4719),
.B(n_4286),
.C(n_4270),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4850),
.Y(n_4905)
);

NAND2xp5_ASAP7_75t_L g4906 ( 
.A(n_4847),
.B(n_4620),
.Y(n_4906)
);

OR2x2_ASAP7_75t_L g4907 ( 
.A(n_4768),
.B(n_4673),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4847),
.Y(n_4908)
);

INVx2_ASAP7_75t_L g4909 ( 
.A(n_4752),
.Y(n_4909)
);

NAND4xp25_ASAP7_75t_L g4910 ( 
.A(n_4818),
.B(n_4688),
.C(n_4637),
.D(n_4618),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4762),
.B(n_4589),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4779),
.B(n_4592),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4728),
.Y(n_4913)
);

OAI22xp5_ASAP7_75t_L g4914 ( 
.A1(n_4821),
.A2(n_4716),
.B1(n_4315),
.B2(n_4653),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4731),
.Y(n_4915)
);

INVx1_ASAP7_75t_L g4916 ( 
.A(n_4733),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4767),
.B(n_4594),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4735),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4767),
.B(n_4763),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4742),
.Y(n_4920)
);

INVx1_ASAP7_75t_SL g4921 ( 
.A(n_4815),
.Y(n_4921)
);

NOR4xp25_ASAP7_75t_L g4922 ( 
.A(n_4744),
.B(n_4628),
.C(n_4641),
.D(n_4627),
.Y(n_4922)
);

INVx3_ASAP7_75t_L g4923 ( 
.A(n_4746),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4732),
.Y(n_4924)
);

AOI32xp33_ASAP7_75t_L g4925 ( 
.A1(n_4760),
.A2(n_4690),
.A3(n_4594),
.B1(n_4530),
.B2(n_4639),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4732),
.Y(n_4926)
);

NOR3xp33_ASAP7_75t_L g4927 ( 
.A(n_4862),
.B(n_4666),
.C(n_4664),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4763),
.B(n_4690),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4801),
.B(n_4608),
.Y(n_4929)
);

OAI32xp33_ASAP7_75t_L g4930 ( 
.A1(n_4816),
.A2(n_4538),
.A3(n_4533),
.B1(n_4449),
.B2(n_4447),
.Y(n_4930)
);

OR2x6_ASAP7_75t_L g4931 ( 
.A(n_4807),
.B(n_4633),
.Y(n_4931)
);

OR2x2_ASAP7_75t_L g4932 ( 
.A(n_4782),
.B(n_4638),
.Y(n_4932)
);

OAI22xp33_ASAP7_75t_SL g4933 ( 
.A1(n_4789),
.A2(n_4694),
.B1(n_4708),
.B2(n_4538),
.Y(n_4933)
);

AND2x2_ASAP7_75t_SL g4934 ( 
.A(n_4831),
.B(n_4796),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_SL g4935 ( 
.A(n_4773),
.B(n_4520),
.Y(n_4935)
);

OAI22xp33_ASAP7_75t_L g4936 ( 
.A1(n_4747),
.A2(n_4273),
.B1(n_4538),
.B2(n_4533),
.Y(n_4936)
);

NAND2x1p5_ASAP7_75t_L g4937 ( 
.A(n_4803),
.B(n_4671),
.Y(n_4937)
);

OR2x2_ASAP7_75t_L g4938 ( 
.A(n_4835),
.B(n_4694),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_4801),
.B(n_4608),
.Y(n_4939)
);

INVx1_ASAP7_75t_L g4940 ( 
.A(n_4736),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4736),
.Y(n_4941)
);

OR2x2_ASAP7_75t_L g4942 ( 
.A(n_4838),
.B(n_4708),
.Y(n_4942)
);

NAND2xp5_ASAP7_75t_SL g4943 ( 
.A(n_4775),
.B(n_4794),
.Y(n_4943)
);

AND2x4_ASAP7_75t_SL g4944 ( 
.A(n_4810),
.B(n_4671),
.Y(n_4944)
);

OAI22xp5_ASAP7_75t_L g4945 ( 
.A1(n_4808),
.A2(n_4843),
.B1(n_4859),
.B2(n_4756),
.Y(n_4945)
);

OAI211xp5_ASAP7_75t_L g4946 ( 
.A1(n_4792),
.A2(n_4369),
.B(n_4680),
.C(n_4665),
.Y(n_4946)
);

A2O1A1Ixp33_ASAP7_75t_L g4947 ( 
.A1(n_4775),
.A2(n_4530),
.B(n_4268),
.C(n_4252),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4789),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4813),
.B(n_4608),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4813),
.B(n_4665),
.Y(n_4950)
);

INVx1_ASAP7_75t_L g4951 ( 
.A(n_4738),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4812),
.B(n_4680),
.Y(n_4952)
);

INVx1_ASAP7_75t_SL g4953 ( 
.A(n_4766),
.Y(n_4953)
);

AND2x2_ASAP7_75t_L g4954 ( 
.A(n_4812),
.B(n_4810),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4766),
.B(n_4645),
.Y(n_4955)
);

NOR2xp33_ASAP7_75t_L g4956 ( 
.A(n_4861),
.B(n_4455),
.Y(n_4956)
);

INVx2_ASAP7_75t_SL g4957 ( 
.A(n_4766),
.Y(n_4957)
);

NAND2xp33_ASAP7_75t_L g4958 ( 
.A(n_4826),
.B(n_4780),
.Y(n_4958)
);

OAI22xp5_ASAP7_75t_L g4959 ( 
.A1(n_4774),
.A2(n_4377),
.B1(n_4308),
.B2(n_4364),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4738),
.Y(n_4960)
);

INVx1_ASAP7_75t_L g4961 ( 
.A(n_4743),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4743),
.Y(n_4962)
);

AOI21xp5_ASAP7_75t_L g4963 ( 
.A1(n_4769),
.A2(n_4440),
.B(n_4711),
.Y(n_4963)
);

INVx2_ASAP7_75t_L g4964 ( 
.A(n_4746),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4776),
.A2(n_4769),
.B1(n_4802),
.B2(n_4811),
.Y(n_4965)
);

AOI22xp5_ASAP7_75t_L g4966 ( 
.A1(n_4806),
.A2(n_4550),
.B1(n_4331),
.B2(n_4528),
.Y(n_4966)
);

AND2x2_ASAP7_75t_L g4967 ( 
.A(n_4826),
.B(n_4530),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4811),
.B(n_4646),
.Y(n_4968)
);

INVx3_ASAP7_75t_L g4969 ( 
.A(n_4746),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4856),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4755),
.B(n_4856),
.Y(n_4971)
);

NOR2xp33_ASAP7_75t_L g4972 ( 
.A(n_4814),
.B(n_4455),
.Y(n_4972)
);

OR2x2_ASAP7_75t_L g4973 ( 
.A(n_4727),
.B(n_4632),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4865),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4865),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4817),
.Y(n_4976)
);

AOI322xp5_ASAP7_75t_L g4977 ( 
.A1(n_4846),
.A2(n_4459),
.A3(n_4695),
.B1(n_4692),
.B2(n_4651),
.C1(n_4657),
.C2(n_4658),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4817),
.Y(n_4978)
);

OAI21xp33_ASAP7_75t_L g4979 ( 
.A1(n_4805),
.A2(n_4550),
.B(n_4531),
.Y(n_4979)
);

OAI21xp33_ASAP7_75t_L g4980 ( 
.A1(n_4783),
.A2(n_4785),
.B(n_4793),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4783),
.B(n_4785),
.Y(n_4981)
);

INVx1_ASAP7_75t_L g4982 ( 
.A(n_4755),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4829),
.B(n_4528),
.Y(n_4983)
);

OAI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_4778),
.A2(n_4650),
.B(n_4647),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4741),
.Y(n_4985)
);

AOI32xp33_ASAP7_75t_L g4986 ( 
.A1(n_4863),
.A2(n_4313),
.A3(n_4332),
.B1(n_4440),
.B2(n_4459),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4745),
.Y(n_4987)
);

AND2x2_ASAP7_75t_L g4988 ( 
.A(n_4919),
.B(n_4829),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_4871),
.B(n_4953),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4912),
.B(n_4837),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4937),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4923),
.Y(n_4992)
);

INVx1_ASAP7_75t_L g4993 ( 
.A(n_4923),
.Y(n_4993)
);

OAI22xp33_ASAP7_75t_L g4994 ( 
.A1(n_4897),
.A2(n_4447),
.B1(n_4449),
.B2(n_4443),
.Y(n_4994)
);

OR2x2_ASAP7_75t_L g4995 ( 
.A(n_4953),
.B(n_4969),
.Y(n_4995)
);

INVx1_ASAP7_75t_SL g4996 ( 
.A(n_4934),
.Y(n_4996)
);

AND2x2_ASAP7_75t_L g4997 ( 
.A(n_4954),
.B(n_4837),
.Y(n_4997)
);

INVxp67_ASAP7_75t_L g4998 ( 
.A(n_4888),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4969),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4957),
.B(n_4841),
.Y(n_5000)
);

NOR2xp33_ASAP7_75t_L g5001 ( 
.A(n_4871),
.B(n_4781),
.Y(n_5001)
);

HB1xp67_ASAP7_75t_L g5002 ( 
.A(n_4937),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4964),
.Y(n_5003)
);

BUFx2_ASAP7_75t_L g5004 ( 
.A(n_4931),
.Y(n_5004)
);

INVx1_ASAP7_75t_L g5005 ( 
.A(n_4889),
.Y(n_5005)
);

INVx1_ASAP7_75t_L g5006 ( 
.A(n_4889),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4895),
.Y(n_5007)
);

HB1xp67_ASAP7_75t_L g5008 ( 
.A(n_4931),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4895),
.Y(n_5009)
);

OR2x2_ASAP7_75t_L g5010 ( 
.A(n_4877),
.B(n_4771),
.Y(n_5010)
);

INVx1_ASAP7_75t_SL g5011 ( 
.A(n_4944),
.Y(n_5011)
);

AND2x2_ASAP7_75t_L g5012 ( 
.A(n_4893),
.B(n_4841),
.Y(n_5012)
);

AND2x4_ASAP7_75t_L g5013 ( 
.A(n_4891),
.B(n_4777),
.Y(n_5013)
);

INVx1_ASAP7_75t_SL g5014 ( 
.A(n_4877),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4891),
.Y(n_5015)
);

INVx1_ASAP7_75t_SL g5016 ( 
.A(n_4921),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4869),
.Y(n_5017)
);

INVxp67_ASAP7_75t_L g5018 ( 
.A(n_4931),
.Y(n_5018)
);

AND2x4_ASAP7_75t_L g5019 ( 
.A(n_4870),
.B(n_4777),
.Y(n_5019)
);

INVx1_ASAP7_75t_L g5020 ( 
.A(n_4873),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4898),
.B(n_4842),
.Y(n_5021)
);

INVx1_ASAP7_75t_L g5022 ( 
.A(n_4874),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4899),
.B(n_4842),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4896),
.B(n_4848),
.Y(n_5024)
);

AO21x2_ASAP7_75t_L g5025 ( 
.A1(n_4875),
.A2(n_4484),
.B(n_4482),
.Y(n_5025)
);

INVx3_ASAP7_75t_L g5026 ( 
.A(n_4882),
.Y(n_5026)
);

INVx1_ASAP7_75t_L g5027 ( 
.A(n_4881),
.Y(n_5027)
);

INVx1_ASAP7_75t_L g5028 ( 
.A(n_4883),
.Y(n_5028)
);

INVx2_ASAP7_75t_SL g5029 ( 
.A(n_4890),
.Y(n_5029)
);

INVx2_ASAP7_75t_L g5030 ( 
.A(n_4901),
.Y(n_5030)
);

HB1xp67_ASAP7_75t_L g5031 ( 
.A(n_4903),
.Y(n_5031)
);

OR2x2_ASAP7_75t_L g5032 ( 
.A(n_4921),
.B(n_4771),
.Y(n_5032)
);

AND2x2_ASAP7_75t_L g5033 ( 
.A(n_4928),
.B(n_4911),
.Y(n_5033)
);

INVx1_ASAP7_75t_SL g5034 ( 
.A(n_4868),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_4905),
.Y(n_5035)
);

OR2x2_ASAP7_75t_L g5036 ( 
.A(n_4981),
.B(n_4730),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_SL g5037 ( 
.A(n_4933),
.B(n_4959),
.Y(n_5037)
);

BUFx3_ASAP7_75t_L g5038 ( 
.A(n_4887),
.Y(n_5038)
);

INVxp67_ASAP7_75t_SL g5039 ( 
.A(n_4958),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_4983),
.B(n_4848),
.Y(n_5040)
);

NAND2xp5_ASAP7_75t_L g5041 ( 
.A(n_4976),
.B(n_4854),
.Y(n_5041)
);

CKINVDCx16_ASAP7_75t_R g5042 ( 
.A(n_4880),
.Y(n_5042)
);

INVx1_ASAP7_75t_SL g5043 ( 
.A(n_4967),
.Y(n_5043)
);

OAI22xp5_ASAP7_75t_L g5044 ( 
.A1(n_4872),
.A2(n_4734),
.B1(n_4765),
.B2(n_4839),
.Y(n_5044)
);

INVx1_ASAP7_75t_L g5045 ( 
.A(n_4955),
.Y(n_5045)
);

INVx1_ASAP7_75t_SL g5046 ( 
.A(n_4949),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_4978),
.B(n_4854),
.Y(n_5047)
);

OR2x2_ASAP7_75t_L g5048 ( 
.A(n_4955),
.B(n_4771),
.Y(n_5048)
);

INVx1_ASAP7_75t_SL g5049 ( 
.A(n_4929),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_4939),
.Y(n_5050)
);

AND2x2_ASAP7_75t_L g5051 ( 
.A(n_4908),
.B(n_4866),
.Y(n_5051)
);

OR2x2_ASAP7_75t_L g5052 ( 
.A(n_4973),
.B(n_4819),
.Y(n_5052)
);

INVx4_ASAP7_75t_L g5053 ( 
.A(n_4902),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4927),
.B(n_4866),
.Y(n_5054)
);

BUFx2_ASAP7_75t_L g5055 ( 
.A(n_4909),
.Y(n_5055)
);

INVx1_ASAP7_75t_SL g5056 ( 
.A(n_4932),
.Y(n_5056)
);

INVx1_ASAP7_75t_L g5057 ( 
.A(n_4952),
.Y(n_5057)
);

INVx3_ASAP7_75t_L g5058 ( 
.A(n_4948),
.Y(n_5058)
);

INVx1_ASAP7_75t_SL g5059 ( 
.A(n_4938),
.Y(n_5059)
);

AO21x2_ASAP7_75t_L g5060 ( 
.A1(n_4984),
.A2(n_4484),
.B(n_4725),
.Y(n_5060)
);

INVx1_ASAP7_75t_SL g5061 ( 
.A(n_4942),
.Y(n_5061)
);

INVx1_ASAP7_75t_SL g5062 ( 
.A(n_4894),
.Y(n_5062)
);

INVx1_ASAP7_75t_SL g5063 ( 
.A(n_4917),
.Y(n_5063)
);

HB1xp67_ASAP7_75t_L g5064 ( 
.A(n_4965),
.Y(n_5064)
);

INVx2_ASAP7_75t_SL g5065 ( 
.A(n_4924),
.Y(n_5065)
);

AOI22xp33_ASAP7_75t_L g5066 ( 
.A1(n_4878),
.A2(n_4440),
.B1(n_4822),
.B2(n_4820),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_4925),
.B(n_4761),
.Y(n_5067)
);

INVx2_ASAP7_75t_SL g5068 ( 
.A(n_4926),
.Y(n_5068)
);

OR2x2_ASAP7_75t_L g5069 ( 
.A(n_4922),
.B(n_4632),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_4982),
.B(n_4761),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4950),
.Y(n_5071)
);

INVx4_ASAP7_75t_L g5072 ( 
.A(n_4940),
.Y(n_5072)
);

INVx1_ASAP7_75t_SL g5073 ( 
.A(n_4884),
.Y(n_5073)
);

HB1xp67_ASAP7_75t_L g5074 ( 
.A(n_4965),
.Y(n_5074)
);

AND2x2_ASAP7_75t_L g5075 ( 
.A(n_4966),
.B(n_4770),
.Y(n_5075)
);

HB1xp67_ASAP7_75t_L g5076 ( 
.A(n_4971),
.Y(n_5076)
);

HB1xp67_ASAP7_75t_L g5077 ( 
.A(n_4971),
.Y(n_5077)
);

NAND3xp33_ASAP7_75t_L g5078 ( 
.A(n_4900),
.B(n_4770),
.C(n_4751),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_4970),
.B(n_4749),
.Y(n_5079)
);

INVx1_ASAP7_75t_L g5080 ( 
.A(n_4884),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4906),
.Y(n_5081)
);

OAI22xp5_ASAP7_75t_L g5082 ( 
.A1(n_4904),
.A2(n_4788),
.B1(n_4784),
.B2(n_4565),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_4980),
.B(n_4759),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4906),
.Y(n_5084)
);

BUFx3_ASAP7_75t_L g5085 ( 
.A(n_4941),
.Y(n_5085)
);

INVx1_ASAP7_75t_L g5086 ( 
.A(n_4951),
.Y(n_5086)
);

INVx1_ASAP7_75t_SL g5087 ( 
.A(n_4943),
.Y(n_5087)
);

AOI22xp33_ASAP7_75t_L g5088 ( 
.A1(n_4879),
.A2(n_4764),
.B1(n_4681),
.B2(n_4685),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4960),
.Y(n_5089)
);

OAI22xp5_ASAP7_75t_L g5090 ( 
.A1(n_4947),
.A2(n_4539),
.B1(n_4536),
.B2(n_4388),
.Y(n_5090)
);

AND2x2_ASAP7_75t_L g5091 ( 
.A(n_4974),
.B(n_4853),
.Y(n_5091)
);

OAI221xp5_ASAP7_75t_L g5092 ( 
.A1(n_4986),
.A2(n_4758),
.B1(n_4786),
.B2(n_4824),
.C(n_4864),
.Y(n_5092)
);

AND2x2_ASAP7_75t_L g5093 ( 
.A(n_4975),
.B(n_4860),
.Y(n_5093)
);

OR2x2_ASAP7_75t_L g5094 ( 
.A(n_4922),
.B(n_4787),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_L g5095 ( 
.A(n_4979),
.B(n_4711),
.Y(n_5095)
);

NAND2xp5_ASAP7_75t_L g5096 ( 
.A(n_4956),
.B(n_4824),
.Y(n_5096)
);

HB1xp67_ASAP7_75t_L g5097 ( 
.A(n_4892),
.Y(n_5097)
);

OAI32xp33_ASAP7_75t_L g5098 ( 
.A1(n_5069),
.A2(n_4914),
.A3(n_4959),
.B1(n_4452),
.B2(n_4446),
.Y(n_5098)
);

NAND2xp5_ASAP7_75t_L g5099 ( 
.A(n_5012),
.B(n_4876),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_5012),
.B(n_4972),
.Y(n_5100)
);

AND2x4_ASAP7_75t_L g5101 ( 
.A(n_5019),
.B(n_4961),
.Y(n_5101)
);

NAND2xp5_ASAP7_75t_L g5102 ( 
.A(n_4988),
.B(n_4962),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5010),
.Y(n_5103)
);

AOI22xp33_ASAP7_75t_L g5104 ( 
.A1(n_4996),
.A2(n_4914),
.B1(n_4885),
.B2(n_4910),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_4988),
.B(n_4963),
.Y(n_5105)
);

NAND2xp5_ASAP7_75t_L g5106 ( 
.A(n_4997),
.B(n_4945),
.Y(n_5106)
);

NAND4xp25_ASAP7_75t_SL g5107 ( 
.A(n_5087),
.B(n_4946),
.C(n_4977),
.D(n_4886),
.Y(n_5107)
);

INVx1_ASAP7_75t_SL g5108 ( 
.A(n_5032),
.Y(n_5108)
);

XOR2x2_ASAP7_75t_L g5109 ( 
.A(n_5043),
.B(n_4935),
.Y(n_5109)
);

INVx1_ASAP7_75t_L g5110 ( 
.A(n_5010),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5032),
.Y(n_5111)
);

INVx1_ASAP7_75t_L g5112 ( 
.A(n_4995),
.Y(n_5112)
);

AOI22xp5_ASAP7_75t_L g5113 ( 
.A1(n_5042),
.A2(n_4910),
.B1(n_4936),
.B2(n_4945),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4995),
.Y(n_5114)
);

NOR2x1_ASAP7_75t_L g5115 ( 
.A(n_5069),
.B(n_4790),
.Y(n_5115)
);

OAI22xp5_ASAP7_75t_L g5116 ( 
.A1(n_5064),
.A2(n_4443),
.B1(n_4449),
.B2(n_4907),
.Y(n_5116)
);

OAI21xp33_ASAP7_75t_L g5117 ( 
.A1(n_5067),
.A2(n_4413),
.B(n_4985),
.Y(n_5117)
);

NAND2xp5_ASAP7_75t_L g5118 ( 
.A(n_4997),
.B(n_4913),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_5023),
.B(n_4915),
.Y(n_5119)
);

OAI222xp33_ASAP7_75t_L g5120 ( 
.A1(n_5094),
.A2(n_5037),
.B1(n_5074),
.B2(n_5048),
.C1(n_5016),
.C2(n_5014),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_5023),
.B(n_4987),
.Y(n_5121)
);

AOI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_5033),
.A2(n_5011),
.B1(n_5075),
.B2(n_5039),
.Y(n_5122)
);

INVx2_ASAP7_75t_L g5123 ( 
.A(n_5013),
.Y(n_5123)
);

NOR2xp33_ASAP7_75t_SL g5124 ( 
.A(n_5048),
.B(n_4916),
.Y(n_5124)
);

AOI22xp5_ASAP7_75t_L g5125 ( 
.A1(n_5033),
.A2(n_4486),
.B1(n_4564),
.B2(n_4558),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_SL g5126 ( 
.A(n_5034),
.B(n_4486),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_5019),
.B(n_4918),
.Y(n_5127)
);

INVx1_ASAP7_75t_L g5128 ( 
.A(n_5013),
.Y(n_5128)
);

OAI211xp5_ASAP7_75t_L g5129 ( 
.A1(n_5037),
.A2(n_5066),
.B(n_5094),
.C(n_5088),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_L g5130 ( 
.A(n_5019),
.B(n_4920),
.Y(n_5130)
);

INVx2_ASAP7_75t_L g5131 ( 
.A(n_5013),
.Y(n_5131)
);

OAI211xp5_ASAP7_75t_L g5132 ( 
.A1(n_5066),
.A2(n_5088),
.B(n_5097),
.C(n_5002),
.Y(n_5132)
);

AOI22xp33_ASAP7_75t_L g5133 ( 
.A1(n_5075),
.A2(n_4563),
.B1(n_4300),
.B2(n_4558),
.Y(n_5133)
);

AOI22xp5_ASAP7_75t_L g5134 ( 
.A1(n_5046),
.A2(n_4564),
.B1(n_4563),
.B2(n_4561),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_5008),
.Y(n_5135)
);

AND2x2_ASAP7_75t_L g5136 ( 
.A(n_5051),
.B(n_4670),
.Y(n_5136)
);

AND2x2_ASAP7_75t_L g5137 ( 
.A(n_5051),
.B(n_4696),
.Y(n_5137)
);

INVxp67_ASAP7_75t_L g5138 ( 
.A(n_5004),
.Y(n_5138)
);

AOI221xp5_ASAP7_75t_L g5139 ( 
.A1(n_4994),
.A2(n_4930),
.B1(n_4984),
.B2(n_4709),
.C(n_4703),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_4989),
.Y(n_5140)
);

AOI21xp5_ASAP7_75t_L g5141 ( 
.A1(n_5024),
.A2(n_4968),
.B(n_4443),
.Y(n_5141)
);

OAI21xp5_ASAP7_75t_SL g5142 ( 
.A1(n_4998),
.A2(n_4968),
.B(n_4830),
.Y(n_5142)
);

AOI222xp33_ASAP7_75t_L g5143 ( 
.A1(n_5018),
.A2(n_4710),
.B1(n_4717),
.B2(n_4721),
.C1(n_4722),
.C2(n_4791),
.Y(n_5143)
);

AOI322xp5_ASAP7_75t_L g5144 ( 
.A1(n_5054),
.A2(n_4800),
.A3(n_4797),
.B1(n_4799),
.B2(n_4840),
.C1(n_4836),
.C2(n_4833),
.Y(n_5144)
);

AOI222xp33_ASAP7_75t_L g5145 ( 
.A1(n_5076),
.A2(n_4852),
.B1(n_4849),
.B2(n_4845),
.C1(n_4832),
.C2(n_4823),
.Y(n_5145)
);

INVx1_ASAP7_75t_L g5146 ( 
.A(n_5026),
.Y(n_5146)
);

OAI22xp33_ASAP7_75t_SL g5147 ( 
.A1(n_4991),
.A2(n_4419),
.B1(n_4474),
.B2(n_4461),
.Y(n_5147)
);

AND2x2_ASAP7_75t_L g5148 ( 
.A(n_5047),
.B(n_4671),
.Y(n_5148)
);

AOI211xp5_ASAP7_75t_SL g5149 ( 
.A1(n_5001),
.A2(n_5026),
.B(n_5015),
.C(n_5006),
.Y(n_5149)
);

AND2x2_ASAP7_75t_L g5150 ( 
.A(n_5047),
.B(n_4554),
.Y(n_5150)
);

INVx1_ASAP7_75t_SL g5151 ( 
.A(n_5052),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4990),
.A2(n_4419),
.B(n_4479),
.Y(n_5152)
);

NOR3xp33_ASAP7_75t_SL g5153 ( 
.A(n_5092),
.B(n_4560),
.C(n_4456),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_5026),
.Y(n_5154)
);

HB1xp67_ASAP7_75t_L g5155 ( 
.A(n_4991),
.Y(n_5155)
);

AOI322xp5_ASAP7_75t_L g5156 ( 
.A1(n_5073),
.A2(n_4377),
.A3(n_4364),
.B1(n_4308),
.B2(n_4328),
.C1(n_4354),
.C2(n_4332),
.Y(n_5156)
);

OAI22xp33_ASAP7_75t_L g5157 ( 
.A1(n_5056),
.A2(n_4444),
.B1(n_4422),
.B2(n_4454),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_SL g5158 ( 
.A(n_5059),
.B(n_4554),
.Y(n_5158)
);

O2A1O1Ixp33_ASAP7_75t_L g5159 ( 
.A1(n_5077),
.A2(n_4488),
.B(n_4495),
.C(n_4487),
.Y(n_5159)
);

AOI22xp33_ASAP7_75t_L g5160 ( 
.A1(n_5038),
.A2(n_4561),
.B1(n_4554),
.B2(n_4346),
.Y(n_5160)
);

INVx1_ASAP7_75t_L g5161 ( 
.A(n_5000),
.Y(n_5161)
);

AOI211xp5_ASAP7_75t_L g5162 ( 
.A1(n_5044),
.A2(n_4368),
.B(n_4488),
.C(n_4487),
.Y(n_5162)
);

INVx1_ASAP7_75t_SL g5163 ( 
.A(n_5052),
.Y(n_5163)
);

INVx1_ASAP7_75t_L g5164 ( 
.A(n_5021),
.Y(n_5164)
);

INVx1_ASAP7_75t_L g5165 ( 
.A(n_5040),
.Y(n_5165)
);

NAND3xp33_ASAP7_75t_L g5166 ( 
.A(n_5001),
.B(n_5078),
.C(n_5007),
.Y(n_5166)
);

NAND3xp33_ASAP7_75t_L g5167 ( 
.A(n_5005),
.B(n_4522),
.C(n_4481),
.Y(n_5167)
);

AOI32xp33_ASAP7_75t_L g5168 ( 
.A1(n_5061),
.A2(n_4561),
.A3(n_4368),
.B1(n_4522),
.B2(n_4504),
.Y(n_5168)
);

AOI21xp33_ASAP7_75t_L g5169 ( 
.A1(n_5062),
.A2(n_4561),
.B(n_4461),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_5038),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_5070),
.Y(n_5171)
);

AOI21xp33_ASAP7_75t_L g5172 ( 
.A1(n_5063),
.A2(n_4411),
.B(n_4465),
.Y(n_5172)
);

OR2x2_ASAP7_75t_L g5173 ( 
.A(n_5041),
.B(n_4552),
.Y(n_5173)
);

OAI22xp5_ASAP7_75t_L g5174 ( 
.A1(n_5083),
.A2(n_4328),
.B1(n_4422),
.B2(n_4464),
.Y(n_5174)
);

OAI32xp33_ASAP7_75t_L g5175 ( 
.A1(n_5009),
.A2(n_4422),
.A3(n_4411),
.B1(n_4474),
.B2(n_4465),
.Y(n_5175)
);

AOI22xp5_ASAP7_75t_L g5176 ( 
.A1(n_5049),
.A2(n_5090),
.B1(n_5082),
.B2(n_5050),
.Y(n_5176)
);

INVx2_ASAP7_75t_SL g5177 ( 
.A(n_5070),
.Y(n_5177)
);

AOI211x1_ASAP7_75t_L g5178 ( 
.A1(n_5095),
.A2(n_4495),
.B(n_4505),
.C(n_4504),
.Y(n_5178)
);

AOI21xp5_ASAP7_75t_L g5179 ( 
.A1(n_5096),
.A2(n_4481),
.B(n_4479),
.Y(n_5179)
);

NAND2xp33_ASAP7_75t_SL g5180 ( 
.A(n_5029),
.B(n_5031),
.Y(n_5180)
);

OAI21xp33_ASAP7_75t_L g5181 ( 
.A1(n_5036),
.A2(n_4518),
.B(n_4552),
.Y(n_5181)
);

INVx2_ASAP7_75t_L g5182 ( 
.A(n_5072),
.Y(n_5182)
);

AOI22xp5_ASAP7_75t_L g5183 ( 
.A1(n_5057),
.A2(n_4474),
.B1(n_4510),
.B2(n_4505),
.Y(n_5183)
);

AOI22xp33_ASAP7_75t_L g5184 ( 
.A1(n_5055),
.A2(n_4347),
.B1(n_4474),
.B2(n_4518),
.Y(n_5184)
);

OR2x2_ASAP7_75t_L g5185 ( 
.A(n_5003),
.B(n_4525),
.Y(n_5185)
);

INVx1_ASAP7_75t_L g5186 ( 
.A(n_5091),
.Y(n_5186)
);

OR2x2_ASAP7_75t_L g5187 ( 
.A(n_4992),
.B(n_4525),
.Y(n_5187)
);

INVx1_ASAP7_75t_L g5188 ( 
.A(n_5091),
.Y(n_5188)
);

AND2x2_ASAP7_75t_L g5189 ( 
.A(n_5071),
.B(n_4510),
.Y(n_5189)
);

AOI211xp5_ASAP7_75t_L g5190 ( 
.A1(n_5120),
.A2(n_5080),
.B(n_4999),
.C(n_4993),
.Y(n_5190)
);

INVx1_ASAP7_75t_L g5191 ( 
.A(n_5101),
.Y(n_5191)
);

NOR2xp67_ASAP7_75t_SL g5192 ( 
.A(n_5166),
.B(n_5170),
.Y(n_5192)
);

AND2x2_ASAP7_75t_L g5193 ( 
.A(n_5150),
.B(n_5079),
.Y(n_5193)
);

INVx1_ASAP7_75t_L g5194 ( 
.A(n_5101),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5128),
.Y(n_5195)
);

OAI22xp5_ASAP7_75t_L g5196 ( 
.A1(n_5104),
.A2(n_5029),
.B1(n_5084),
.B2(n_5081),
.Y(n_5196)
);

O2A1O1Ixp33_ASAP7_75t_SL g5197 ( 
.A1(n_5108),
.A2(n_5065),
.B(n_5068),
.C(n_5045),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_L g5198 ( 
.A(n_5148),
.B(n_5058),
.Y(n_5198)
);

AOI21xp33_ASAP7_75t_L g5199 ( 
.A1(n_5151),
.A2(n_5035),
.B(n_5030),
.Y(n_5199)
);

OAI22xp33_ASAP7_75t_L g5200 ( 
.A1(n_5113),
.A2(n_5072),
.B1(n_4422),
.B2(n_5035),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_L g5201 ( 
.A(n_5151),
.B(n_5053),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_5123),
.Y(n_5202)
);

NOR2xp33_ASAP7_75t_L g5203 ( 
.A(n_5163),
.B(n_5053),
.Y(n_5203)
);

INVx1_ASAP7_75t_SL g5204 ( 
.A(n_5163),
.Y(n_5204)
);

AOI22xp5_ASAP7_75t_L g5205 ( 
.A1(n_5129),
.A2(n_5079),
.B1(n_5058),
.B2(n_5093),
.Y(n_5205)
);

HB1xp67_ASAP7_75t_L g5206 ( 
.A(n_5115),
.Y(n_5206)
);

CKINVDCx16_ASAP7_75t_R g5207 ( 
.A(n_5122),
.Y(n_5207)
);

INVx1_ASAP7_75t_L g5208 ( 
.A(n_5131),
.Y(n_5208)
);

INVx1_ASAP7_75t_L g5209 ( 
.A(n_5105),
.Y(n_5209)
);

OAI22xp5_ASAP7_75t_L g5210 ( 
.A1(n_5133),
.A2(n_5058),
.B1(n_5017),
.B2(n_5022),
.Y(n_5210)
);

INVx2_ASAP7_75t_SL g5211 ( 
.A(n_5177),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5136),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_5125),
.B(n_5093),
.Y(n_5213)
);

OAI22xp5_ASAP7_75t_SL g5214 ( 
.A1(n_5106),
.A2(n_5068),
.B1(n_5065),
.B2(n_5053),
.Y(n_5214)
);

INVx1_ASAP7_75t_L g5215 ( 
.A(n_5137),
.Y(n_5215)
);

AOI21xp5_ASAP7_75t_L g5216 ( 
.A1(n_5108),
.A2(n_5060),
.B(n_5030),
.Y(n_5216)
);

AOI211xp5_ASAP7_75t_SL g5217 ( 
.A1(n_5132),
.A2(n_5027),
.B(n_5028),
.C(n_5020),
.Y(n_5217)
);

INVx1_ASAP7_75t_L g5218 ( 
.A(n_5127),
.Y(n_5218)
);

OAI22xp33_ASAP7_75t_L g5219 ( 
.A1(n_5124),
.A2(n_5072),
.B1(n_5085),
.B2(n_4417),
.Y(n_5219)
);

INVx1_ASAP7_75t_L g5220 ( 
.A(n_5130),
.Y(n_5220)
);

AOI222xp33_ASAP7_75t_L g5221 ( 
.A1(n_5139),
.A2(n_5085),
.B1(n_5089),
.B2(n_5086),
.C1(n_4548),
.C2(n_4543),
.Y(n_5221)
);

NOR4xp25_ASAP7_75t_SL g5222 ( 
.A(n_5180),
.B(n_4517),
.C(n_4526),
.D(n_4513),
.Y(n_5222)
);

OAI22xp33_ASAP7_75t_SL g5223 ( 
.A1(n_5124),
.A2(n_4517),
.B1(n_4526),
.B2(n_4513),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_L g5224 ( 
.A(n_5171),
.B(n_4542),
.Y(n_5224)
);

INVx3_ASAP7_75t_L g5225 ( 
.A(n_5182),
.Y(n_5225)
);

AOI222xp33_ASAP7_75t_L g5226 ( 
.A1(n_5111),
.A2(n_4542),
.B1(n_4543),
.B2(n_4546),
.C1(n_4555),
.C2(n_4548),
.Y(n_5226)
);

OAI31xp33_ASAP7_75t_L g5227 ( 
.A1(n_5107),
.A2(n_4546),
.A3(n_4555),
.B(n_4549),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5146),
.Y(n_5228)
);

NOR2xp33_ASAP7_75t_L g5229 ( 
.A(n_5112),
.B(n_5060),
.Y(n_5229)
);

AOI21xp33_ASAP7_75t_L g5230 ( 
.A1(n_5114),
.A2(n_5060),
.B(n_5025),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_5149),
.B(n_4549),
.Y(n_5231)
);

INVx1_ASAP7_75t_L g5232 ( 
.A(n_5154),
.Y(n_5232)
);

NAND2xp33_ASAP7_75t_SL g5233 ( 
.A(n_5185),
.B(n_4551),
.Y(n_5233)
);

AOI21xp33_ASAP7_75t_L g5234 ( 
.A1(n_5138),
.A2(n_5147),
.B(n_5140),
.Y(n_5234)
);

INVx2_ASAP7_75t_L g5235 ( 
.A(n_5187),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5103),
.Y(n_5236)
);

AOI21xp33_ASAP7_75t_SL g5237 ( 
.A1(n_5168),
.A2(n_5025),
.B(n_4551),
.Y(n_5237)
);

NOR2xp33_ASAP7_75t_L g5238 ( 
.A(n_5158),
.B(n_5025),
.Y(n_5238)
);

NAND2xp5_ASAP7_75t_L g5239 ( 
.A(n_5149),
.B(n_4351),
.Y(n_5239)
);

INVx1_ASAP7_75t_L g5240 ( 
.A(n_5110),
.Y(n_5240)
);

INVx1_ASAP7_75t_L g5241 ( 
.A(n_5109),
.Y(n_5241)
);

AOI32xp33_ASAP7_75t_L g5242 ( 
.A1(n_5135),
.A2(n_4417),
.A3(n_4354),
.B1(n_4356),
.B2(n_4370),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5155),
.Y(n_5243)
);

AOI321xp33_ASAP7_75t_L g5244 ( 
.A1(n_5098),
.A2(n_4417),
.A3(n_4588),
.B1(n_4357),
.B2(n_4000),
.C(n_3941),
.Y(n_5244)
);

INVx1_ASAP7_75t_L g5245 ( 
.A(n_5102),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_5134),
.B(n_4033),
.Y(n_5246)
);

INVxp33_ASAP7_75t_L g5247 ( 
.A(n_5126),
.Y(n_5247)
);

NAND4xp25_ASAP7_75t_SL g5248 ( 
.A(n_5160),
.B(n_4371),
.C(n_4164),
.D(n_4160),
.Y(n_5248)
);

AOI22xp33_ASAP7_75t_L g5249 ( 
.A1(n_5174),
.A2(n_4000),
.B1(n_3973),
.B2(n_3941),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5121),
.Y(n_5250)
);

INVx3_ASAP7_75t_L g5251 ( 
.A(n_5186),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_SL g5252 ( 
.A(n_5184),
.B(n_3973),
.Y(n_5252)
);

OAI22xp5_ASAP7_75t_L g5253 ( 
.A1(n_5176),
.A2(n_4034),
.B1(n_4164),
.B2(n_4160),
.Y(n_5253)
);

OAI211xp5_ASAP7_75t_L g5254 ( 
.A1(n_5145),
.A2(n_4000),
.B(n_3973),
.C(n_4371),
.Y(n_5254)
);

NAND2xp5_ASAP7_75t_L g5255 ( 
.A(n_5188),
.B(n_4033),
.Y(n_5255)
);

AND2x2_ASAP7_75t_L g5256 ( 
.A(n_5153),
.B(n_3896),
.Y(n_5256)
);

AND2x2_ASAP7_75t_L g5257 ( 
.A(n_5161),
.B(n_3712),
.Y(n_5257)
);

INVx2_ASAP7_75t_L g5258 ( 
.A(n_5173),
.Y(n_5258)
);

AOI311xp33_ASAP7_75t_L g5259 ( 
.A1(n_5169),
.A2(n_4034),
.A3(n_4156),
.B(n_4069),
.C(n_4066),
.Y(n_5259)
);

NOR2x1_ASAP7_75t_L g5260 ( 
.A(n_5116),
.B(n_3973),
.Y(n_5260)
);

AND2x2_ASAP7_75t_L g5261 ( 
.A(n_5164),
.B(n_3712),
.Y(n_5261)
);

INVx1_ASAP7_75t_L g5262 ( 
.A(n_5118),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_SL g5263 ( 
.A(n_5099),
.B(n_4000),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_5119),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5152),
.B(n_4041),
.Y(n_5265)
);

INVx1_ASAP7_75t_L g5266 ( 
.A(n_5100),
.Y(n_5266)
);

NAND2xp5_ASAP7_75t_L g5267 ( 
.A(n_5144),
.B(n_4041),
.Y(n_5267)
);

OAI322xp33_ASAP7_75t_L g5268 ( 
.A1(n_5174),
.A2(n_4071),
.A3(n_4015),
.B1(n_4037),
.B2(n_3956),
.C1(n_3975),
.C2(n_3951),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_5206),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5206),
.Y(n_5270)
);

OR2x2_ASAP7_75t_L g5271 ( 
.A(n_5191),
.B(n_5165),
.Y(n_5271)
);

OR2x2_ASAP7_75t_L g5272 ( 
.A(n_5194),
.B(n_5142),
.Y(n_5272)
);

NOR2xp33_ASAP7_75t_L g5273 ( 
.A(n_5247),
.B(n_5181),
.Y(n_5273)
);

INVx2_ASAP7_75t_L g5274 ( 
.A(n_5260),
.Y(n_5274)
);

INVx1_ASAP7_75t_SL g5275 ( 
.A(n_5233),
.Y(n_5275)
);

INVx1_ASAP7_75t_SL g5276 ( 
.A(n_5193),
.Y(n_5276)
);

INVx1_ASAP7_75t_L g5277 ( 
.A(n_5198),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_SL g5278 ( 
.A(n_5216),
.B(n_5116),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5201),
.Y(n_5279)
);

AND2x2_ASAP7_75t_L g5280 ( 
.A(n_5207),
.B(n_5117),
.Y(n_5280)
);

AND2x2_ASAP7_75t_L g5281 ( 
.A(n_5261),
.B(n_5189),
.Y(n_5281)
);

INVx1_ASAP7_75t_L g5282 ( 
.A(n_5201),
.Y(n_5282)
);

NAND2xp5_ASAP7_75t_L g5283 ( 
.A(n_5251),
.B(n_5141),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_5251),
.Y(n_5284)
);

OR2x2_ASAP7_75t_L g5285 ( 
.A(n_5204),
.B(n_5167),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_5203),
.B(n_5205),
.Y(n_5286)
);

INVx1_ASAP7_75t_SL g5287 ( 
.A(n_5214),
.Y(n_5287)
);

AND2x2_ASAP7_75t_L g5288 ( 
.A(n_5257),
.B(n_5172),
.Y(n_5288)
);

NAND2x1p5_ASAP7_75t_L g5289 ( 
.A(n_5225),
.B(n_5183),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_5225),
.B(n_5143),
.Y(n_5290)
);

NAND2xp5_ASAP7_75t_SL g5291 ( 
.A(n_5216),
.B(n_5156),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_5238),
.Y(n_5292)
);

NOR2xp33_ASAP7_75t_L g5293 ( 
.A(n_5199),
.B(n_5175),
.Y(n_5293)
);

NAND2xp5_ASAP7_75t_L g5294 ( 
.A(n_5211),
.B(n_5143),
.Y(n_5294)
);

NAND2xp5_ASAP7_75t_L g5295 ( 
.A(n_5250),
.B(n_5162),
.Y(n_5295)
);

AOI22xp33_ASAP7_75t_L g5296 ( 
.A1(n_5248),
.A2(n_5192),
.B1(n_5196),
.B2(n_5256),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_5243),
.B(n_5157),
.Y(n_5297)
);

NOR2x1_ASAP7_75t_L g5298 ( 
.A(n_5219),
.B(n_5159),
.Y(n_5298)
);

AND2x4_ASAP7_75t_L g5299 ( 
.A(n_5235),
.B(n_5179),
.Y(n_5299)
);

NOR2xp33_ASAP7_75t_L g5300 ( 
.A(n_5237),
.B(n_5178),
.Y(n_5300)
);

AOI22xp33_ASAP7_75t_L g5301 ( 
.A1(n_5227),
.A2(n_5145),
.B1(n_4071),
.B2(n_4037),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_5238),
.Y(n_5302)
);

OR2x2_ASAP7_75t_L g5303 ( 
.A(n_5213),
.B(n_4044),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5212),
.B(n_4044),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_L g5305 ( 
.A(n_5215),
.B(n_5202),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_5208),
.B(n_4052),
.Y(n_5306)
);

OR2x2_ASAP7_75t_L g5307 ( 
.A(n_5210),
.B(n_5195),
.Y(n_5307)
);

INVxp67_ASAP7_75t_SL g5308 ( 
.A(n_5219),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_SL g5309 ( 
.A(n_5223),
.B(n_4052),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_5236),
.B(n_4056),
.Y(n_5310)
);

AND2x4_ASAP7_75t_L g5311 ( 
.A(n_5258),
.B(n_4056),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_5240),
.B(n_4059),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5190),
.B(n_5221),
.Y(n_5313)
);

INVx1_ASAP7_75t_L g5314 ( 
.A(n_5231),
.Y(n_5314)
);

INVx1_ASAP7_75t_L g5315 ( 
.A(n_5229),
.Y(n_5315)
);

NOR2xp33_ASAP7_75t_L g5316 ( 
.A(n_5197),
.B(n_4059),
.Y(n_5316)
);

INVx2_ASAP7_75t_L g5317 ( 
.A(n_5228),
.Y(n_5317)
);

INVx1_ASAP7_75t_L g5318 ( 
.A(n_5229),
.Y(n_5318)
);

NAND2xp5_ASAP7_75t_L g5319 ( 
.A(n_5217),
.B(n_5241),
.Y(n_5319)
);

INVx1_ASAP7_75t_L g5320 ( 
.A(n_5239),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5232),
.B(n_5200),
.Y(n_5321)
);

INVx2_ASAP7_75t_L g5322 ( 
.A(n_5218),
.Y(n_5322)
);

NAND2x1_ASAP7_75t_L g5323 ( 
.A(n_5249),
.B(n_4015),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_5220),
.B(n_4062),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_5224),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_5200),
.B(n_4062),
.Y(n_5326)
);

INVx1_ASAP7_75t_L g5327 ( 
.A(n_5246),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_SL g5328 ( 
.A(n_5244),
.B(n_4064),
.Y(n_5328)
);

OR2x2_ASAP7_75t_L g5329 ( 
.A(n_5267),
.B(n_4064),
.Y(n_5329)
);

INVx1_ASAP7_75t_L g5330 ( 
.A(n_5265),
.Y(n_5330)
);

AND2x2_ASAP7_75t_L g5331 ( 
.A(n_5245),
.B(n_3712),
.Y(n_5331)
);

INVx1_ASAP7_75t_L g5332 ( 
.A(n_5255),
.Y(n_5332)
);

INVx1_ASAP7_75t_L g5333 ( 
.A(n_5226),
.Y(n_5333)
);

OR2x2_ASAP7_75t_L g5334 ( 
.A(n_5262),
.B(n_4066),
.Y(n_5334)
);

AND2x2_ASAP7_75t_L g5335 ( 
.A(n_5266),
.B(n_3718),
.Y(n_5335)
);

INVx1_ASAP7_75t_SL g5336 ( 
.A(n_5234),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5276),
.B(n_5242),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_SL g5338 ( 
.A(n_5275),
.B(n_5259),
.Y(n_5338)
);

HB1xp67_ASAP7_75t_L g5339 ( 
.A(n_5289),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_5289),
.Y(n_5340)
);

OAI321xp33_ASAP7_75t_L g5341 ( 
.A1(n_5319),
.A2(n_5253),
.A3(n_5264),
.B1(n_5209),
.B2(n_5252),
.C(n_5263),
.Y(n_5341)
);

AOI211x1_ASAP7_75t_L g5342 ( 
.A1(n_5291),
.A2(n_5328),
.B(n_5254),
.C(n_5278),
.Y(n_5342)
);

INVx1_ASAP7_75t_L g5343 ( 
.A(n_5283),
.Y(n_5343)
);

XOR2x2_ASAP7_75t_L g5344 ( 
.A(n_5273),
.B(n_5222),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_SL g5345 ( 
.A(n_5299),
.B(n_5230),
.Y(n_5345)
);

NAND2xp5_ASAP7_75t_L g5346 ( 
.A(n_5284),
.B(n_5254),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5308),
.Y(n_5347)
);

INVx1_ASAP7_75t_L g5348 ( 
.A(n_5308),
.Y(n_5348)
);

AOI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_5278),
.A2(n_5268),
.B(n_5249),
.Y(n_5349)
);

AOI221xp5_ASAP7_75t_SL g5350 ( 
.A1(n_5291),
.A2(n_4037),
.B1(n_4015),
.B2(n_3951),
.C(n_3953),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5290),
.Y(n_5351)
);

NOR2x1_ASAP7_75t_L g5352 ( 
.A(n_5298),
.B(n_4015),
.Y(n_5352)
);

NOR2xp33_ASAP7_75t_L g5353 ( 
.A(n_5336),
.B(n_4069),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5284),
.B(n_5281),
.Y(n_5354)
);

NOR2xp33_ASAP7_75t_SL g5355 ( 
.A(n_5273),
.B(n_4077),
.Y(n_5355)
);

AOI21xp5_ASAP7_75t_L g5356 ( 
.A1(n_5286),
.A2(n_5300),
.B(n_5309),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5272),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_5288),
.Y(n_5358)
);

AOI221xp5_ASAP7_75t_L g5359 ( 
.A1(n_5300),
.A2(n_4071),
.B1(n_4037),
.B2(n_3951),
.C(n_3953),
.Y(n_5359)
);

AOI221xp5_ASAP7_75t_L g5360 ( 
.A1(n_5293),
.A2(n_3948),
.B1(n_3950),
.B2(n_3953),
.C(n_3956),
.Y(n_5360)
);

NOR3x1_ASAP7_75t_L g5361 ( 
.A(n_5313),
.B(n_4082),
.C(n_4077),
.Y(n_5361)
);

NAND2xp5_ASAP7_75t_L g5362 ( 
.A(n_5331),
.B(n_5335),
.Y(n_5362)
);

AO22x2_ASAP7_75t_L g5363 ( 
.A1(n_5269),
.A2(n_5270),
.B1(n_5333),
.B2(n_5274),
.Y(n_5363)
);

NAND3xp33_ASAP7_75t_SL g5364 ( 
.A(n_5287),
.B(n_4086),
.C(n_4082),
.Y(n_5364)
);

NAND2xp5_ASAP7_75t_L g5365 ( 
.A(n_5299),
.B(n_4086),
.Y(n_5365)
);

NOR2x1_ASAP7_75t_L g5366 ( 
.A(n_5274),
.B(n_4087),
.Y(n_5366)
);

NOR2xp33_ASAP7_75t_L g5367 ( 
.A(n_5307),
.B(n_4087),
.Y(n_5367)
);

INVx1_ASAP7_75t_L g5368 ( 
.A(n_5294),
.Y(n_5368)
);

AOI22xp5_ASAP7_75t_L g5369 ( 
.A1(n_5280),
.A2(n_4111),
.B1(n_4156),
.B2(n_4096),
.Y(n_5369)
);

NAND5xp2_ASAP7_75t_L g5370 ( 
.A(n_5296),
.B(n_4111),
.C(n_4096),
.D(n_4127),
.E(n_4144),
.Y(n_5370)
);

AOI22xp5_ASAP7_75t_L g5371 ( 
.A1(n_5293),
.A2(n_4134),
.B1(n_4120),
.B2(n_4117),
.Y(n_5371)
);

NAND2xp5_ASAP7_75t_L g5372 ( 
.A(n_5316),
.B(n_4113),
.Y(n_5372)
);

NOR3xp33_ASAP7_75t_L g5373 ( 
.A(n_5279),
.B(n_4117),
.C(n_4113),
.Y(n_5373)
);

NOR2xp33_ASAP7_75t_SL g5374 ( 
.A(n_5285),
.B(n_4120),
.Y(n_5374)
);

AND2x2_ASAP7_75t_L g5375 ( 
.A(n_5282),
.B(n_4121),
.Y(n_5375)
);

AOI211xp5_ASAP7_75t_L g5376 ( 
.A1(n_5316),
.A2(n_4137),
.B(n_4125),
.C(n_4121),
.Y(n_5376)
);

NOR3xp33_ASAP7_75t_L g5377 ( 
.A(n_5305),
.B(n_4127),
.C(n_4125),
.Y(n_5377)
);

AOI21xp5_ASAP7_75t_L g5378 ( 
.A1(n_5309),
.A2(n_4134),
.B(n_4131),
.Y(n_5378)
);

AND4x1_ASAP7_75t_L g5379 ( 
.A(n_5296),
.B(n_4136),
.C(n_4144),
.D(n_4141),
.Y(n_5379)
);

AOI221xp5_ASAP7_75t_SL g5380 ( 
.A1(n_5328),
.A2(n_3948),
.B1(n_3950),
.B2(n_3956),
.C(n_3975),
.Y(n_5380)
);

AO21x1_ASAP7_75t_L g5381 ( 
.A1(n_5323),
.A2(n_3975),
.B(n_3993),
.Y(n_5381)
);

NOR4xp25_ASAP7_75t_L g5382 ( 
.A(n_5297),
.B(n_4131),
.C(n_4136),
.D(n_4137),
.Y(n_5382)
);

OAI221xp5_ASAP7_75t_SL g5383 ( 
.A1(n_5271),
.A2(n_4140),
.B1(n_4141),
.B2(n_4147),
.C(n_4148),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_5321),
.Y(n_5384)
);

NAND3xp33_ASAP7_75t_SL g5385 ( 
.A(n_5295),
.B(n_4140),
.C(n_3994),
.Y(n_5385)
);

NAND2xp5_ASAP7_75t_L g5386 ( 
.A(n_5311),
.B(n_3993),
.Y(n_5386)
);

AOI21xp5_ASAP7_75t_L g5387 ( 
.A1(n_5315),
.A2(n_3994),
.B(n_3993),
.Y(n_5387)
);

NOR3x1_ASAP7_75t_L g5388 ( 
.A(n_5277),
.B(n_3814),
.C(n_3809),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_5311),
.Y(n_5389)
);

HB1xp67_ASAP7_75t_L g5390 ( 
.A(n_5324),
.Y(n_5390)
);

AOI221xp5_ASAP7_75t_L g5391 ( 
.A1(n_5301),
.A2(n_4159),
.B1(n_4148),
.B2(n_4147),
.C(n_4128),
.Y(n_5391)
);

NAND2xp5_ASAP7_75t_L g5392 ( 
.A(n_5347),
.B(n_5314),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_5390),
.Y(n_5393)
);

AND3x1_ASAP7_75t_L g5394 ( 
.A(n_5370),
.B(n_5317),
.C(n_5322),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_5339),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_5348),
.B(n_5320),
.Y(n_5396)
);

NAND2xp5_ASAP7_75t_L g5397 ( 
.A(n_5342),
.B(n_5324),
.Y(n_5397)
);

NAND2xp5_ASAP7_75t_L g5398 ( 
.A(n_5340),
.B(n_5330),
.Y(n_5398)
);

AOI22xp5_ASAP7_75t_L g5399 ( 
.A1(n_5357),
.A2(n_5327),
.B1(n_5325),
.B2(n_5302),
.Y(n_5399)
);

HB1xp67_ASAP7_75t_L g5400 ( 
.A(n_5352),
.Y(n_5400)
);

NAND3xp33_ASAP7_75t_L g5401 ( 
.A(n_5379),
.B(n_5301),
.C(n_5292),
.Y(n_5401)
);

NAND3xp33_ASAP7_75t_L g5402 ( 
.A(n_5374),
.B(n_5332),
.C(n_5318),
.Y(n_5402)
);

AND2x2_ASAP7_75t_L g5403 ( 
.A(n_5388),
.B(n_5303),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5349),
.B(n_5306),
.Y(n_5404)
);

OAI321xp33_ASAP7_75t_L g5405 ( 
.A1(n_5337),
.A2(n_5329),
.A3(n_5304),
.B1(n_5312),
.B2(n_5310),
.C(n_5326),
.Y(n_5405)
);

NOR2xp33_ASAP7_75t_L g5406 ( 
.A(n_5354),
.B(n_5334),
.Y(n_5406)
);

NAND3xp33_ASAP7_75t_L g5407 ( 
.A(n_5356),
.B(n_3999),
.C(n_3994),
.Y(n_5407)
);

AND2x2_ASAP7_75t_L g5408 ( 
.A(n_5384),
.B(n_3718),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5363),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5363),
.Y(n_5410)
);

AOI22xp33_ASAP7_75t_L g5411 ( 
.A1(n_5368),
.A2(n_4159),
.B1(n_4148),
.B2(n_4147),
.Y(n_5411)
);

NOR2xp33_ASAP7_75t_L g5412 ( 
.A(n_5341),
.B(n_3718),
.Y(n_5412)
);

NAND3xp33_ASAP7_75t_L g5413 ( 
.A(n_5355),
.B(n_4016),
.C(n_3999),
.Y(n_5413)
);

NAND2xp5_ASAP7_75t_L g5414 ( 
.A(n_5363),
.B(n_3902),
.Y(n_5414)
);

AOI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_5345),
.A2(n_4016),
.B(n_3999),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5362),
.Y(n_5416)
);

HB1xp67_ASAP7_75t_L g5417 ( 
.A(n_5366),
.Y(n_5417)
);

AOI22xp5_ASAP7_75t_L g5418 ( 
.A1(n_5358),
.A2(n_3723),
.B1(n_3775),
.B2(n_4124),
.Y(n_5418)
);

NAND2xp5_ASAP7_75t_L g5419 ( 
.A(n_5375),
.B(n_3793),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_5389),
.Y(n_5420)
);

NAND4xp25_ASAP7_75t_L g5421 ( 
.A(n_5370),
.B(n_5338),
.C(n_5361),
.D(n_5353),
.Y(n_5421)
);

NAND2xp5_ASAP7_75t_L g5422 ( 
.A(n_5367),
.B(n_3798),
.Y(n_5422)
);

INVx1_ASAP7_75t_L g5423 ( 
.A(n_5372),
.Y(n_5423)
);

NAND5xp2_ASAP7_75t_L g5424 ( 
.A(n_5351),
.B(n_3796),
.C(n_3509),
.D(n_3510),
.E(n_3479),
.Y(n_5424)
);

O2A1O1Ixp5_ASAP7_75t_L g5425 ( 
.A1(n_5381),
.A2(n_4029),
.B(n_4128),
.C(n_4124),
.Y(n_5425)
);

NOR2xp33_ASAP7_75t_L g5426 ( 
.A(n_5343),
.B(n_3723),
.Y(n_5426)
);

NOR2xp33_ASAP7_75t_L g5427 ( 
.A(n_5385),
.B(n_4159),
.Y(n_5427)
);

INVx1_ASAP7_75t_L g5428 ( 
.A(n_5372),
.Y(n_5428)
);

AOI211x1_ASAP7_75t_L g5429 ( 
.A1(n_5364),
.A2(n_3904),
.B(n_3901),
.C(n_3899),
.Y(n_5429)
);

INVx1_ASAP7_75t_L g5430 ( 
.A(n_5344),
.Y(n_5430)
);

AOI211xp5_ASAP7_75t_L g5431 ( 
.A1(n_5383),
.A2(n_4128),
.B(n_4124),
.C(n_4123),
.Y(n_5431)
);

NOR2xp33_ASAP7_75t_L g5432 ( 
.A(n_5346),
.B(n_3723),
.Y(n_5432)
);

NAND4xp25_ASAP7_75t_SL g5433 ( 
.A(n_5350),
.B(n_4123),
.C(n_4112),
.D(n_4085),
.Y(n_5433)
);

NOR2xp33_ASAP7_75t_L g5434 ( 
.A(n_5365),
.B(n_3809),
.Y(n_5434)
);

NAND2xp5_ASAP7_75t_L g5435 ( 
.A(n_5371),
.B(n_3799),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_5386),
.Y(n_5436)
);

NOR2xp33_ASAP7_75t_L g5437 ( 
.A(n_5369),
.B(n_3814),
.Y(n_5437)
);

NAND4xp75_ASAP7_75t_L g5438 ( 
.A(n_5380),
.B(n_4123),
.C(n_4112),
.D(n_4085),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5386),
.Y(n_5439)
);

NOR2xp33_ASAP7_75t_L g5440 ( 
.A(n_5393),
.B(n_5378),
.Y(n_5440)
);

NAND2xp5_ASAP7_75t_SL g5441 ( 
.A(n_5394),
.B(n_5382),
.Y(n_5441)
);

NOR3x1_ASAP7_75t_L g5442 ( 
.A(n_5421),
.B(n_5373),
.C(n_5377),
.Y(n_5442)
);

A2O1A1Ixp33_ASAP7_75t_L g5443 ( 
.A1(n_5412),
.A2(n_5387),
.B(n_5376),
.C(n_5359),
.Y(n_5443)
);

OAI211xp5_ASAP7_75t_L g5444 ( 
.A1(n_5399),
.A2(n_5397),
.B(n_5395),
.C(n_5392),
.Y(n_5444)
);

NAND4xp25_ASAP7_75t_SL g5445 ( 
.A(n_5418),
.B(n_5360),
.C(n_5391),
.D(n_4112),
.Y(n_5445)
);

AND4x1_ASAP7_75t_L g5446 ( 
.A(n_5406),
.B(n_3822),
.C(n_3838),
.D(n_3808),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_5408),
.B(n_3799),
.Y(n_5447)
);

CKINVDCx5p33_ASAP7_75t_R g5448 ( 
.A(n_5416),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_5432),
.B(n_3822),
.Y(n_5449)
);

NAND2xp5_ASAP7_75t_L g5450 ( 
.A(n_5426),
.B(n_5403),
.Y(n_5450)
);

NAND4xp25_ASAP7_75t_L g5451 ( 
.A(n_5430),
.B(n_4085),
.C(n_4079),
.D(n_4075),
.Y(n_5451)
);

OAI21xp5_ASAP7_75t_L g5452 ( 
.A1(n_5402),
.A2(n_4079),
.B(n_4075),
.Y(n_5452)
);

NAND4xp25_ASAP7_75t_L g5453 ( 
.A(n_5404),
.B(n_4079),
.C(n_4075),
.D(n_4070),
.Y(n_5453)
);

OAI211xp5_ASAP7_75t_L g5454 ( 
.A1(n_5409),
.A2(n_4070),
.B(n_4050),
.C(n_4043),
.Y(n_5454)
);

NAND2xp5_ASAP7_75t_L g5455 ( 
.A(n_5410),
.B(n_3845),
.Y(n_5455)
);

NOR3x1_ASAP7_75t_L g5456 ( 
.A(n_5401),
.B(n_3882),
.C(n_3849),
.Y(n_5456)
);

NOR3x1_ASAP7_75t_L g5457 ( 
.A(n_5396),
.B(n_3882),
.C(n_3849),
.Y(n_5457)
);

AOI22xp5_ASAP7_75t_L g5458 ( 
.A1(n_5420),
.A2(n_4070),
.B1(n_4050),
.B2(n_4043),
.Y(n_5458)
);

NAND5xp2_ASAP7_75t_L g5459 ( 
.A(n_5405),
.B(n_3509),
.C(n_3510),
.D(n_3469),
.E(n_3479),
.Y(n_5459)
);

AOI211xp5_ASAP7_75t_L g5460 ( 
.A1(n_5407),
.A2(n_4050),
.B(n_4043),
.C(n_4042),
.Y(n_5460)
);

AOI211xp5_ASAP7_75t_L g5461 ( 
.A1(n_5398),
.A2(n_4042),
.B(n_4029),
.C(n_4028),
.Y(n_5461)
);

NAND2xp5_ASAP7_75t_L g5462 ( 
.A(n_5437),
.B(n_3845),
.Y(n_5462)
);

AOI211xp5_ASAP7_75t_L g5463 ( 
.A1(n_5415),
.A2(n_4042),
.B(n_4029),
.C(n_4028),
.Y(n_5463)
);

NAND4xp25_ASAP7_75t_L g5464 ( 
.A(n_5427),
.B(n_4028),
.C(n_4025),
.D(n_4021),
.Y(n_5464)
);

OAI211xp5_ASAP7_75t_L g5465 ( 
.A1(n_5417),
.A2(n_4025),
.B(n_4021),
.C(n_4020),
.Y(n_5465)
);

AOI22xp5_ASAP7_75t_L g5466 ( 
.A1(n_5434),
.A2(n_4025),
.B1(n_4021),
.B2(n_4020),
.Y(n_5466)
);

NAND3xp33_ASAP7_75t_L g5467 ( 
.A(n_5417),
.B(n_4020),
.C(n_4017),
.Y(n_5467)
);

A2O1A1Ixp33_ASAP7_75t_L g5468 ( 
.A1(n_5427),
.A2(n_5413),
.B(n_5414),
.C(n_5400),
.Y(n_5468)
);

OAI22xp5_ASAP7_75t_L g5469 ( 
.A1(n_5411),
.A2(n_4017),
.B1(n_4016),
.B2(n_3702),
.Y(n_5469)
);

NAND4xp75_ASAP7_75t_L g5470 ( 
.A(n_5423),
.B(n_5428),
.C(n_5436),
.D(n_5439),
.Y(n_5470)
);

NOR3xp33_ASAP7_75t_L g5471 ( 
.A(n_5400),
.B(n_4017),
.C(n_3699),
.Y(n_5471)
);

NOR2x1p5_ASAP7_75t_L g5472 ( 
.A(n_5422),
.B(n_3561),
.Y(n_5472)
);

NOR2xp33_ASAP7_75t_L g5473 ( 
.A(n_5419),
.B(n_3561),
.Y(n_5473)
);

NOR2x1_ASAP7_75t_L g5474 ( 
.A(n_5433),
.B(n_3572),
.Y(n_5474)
);

OA211x2_ASAP7_75t_L g5475 ( 
.A1(n_5411),
.A2(n_3610),
.B(n_3607),
.C(n_3606),
.Y(n_5475)
);

NAND3xp33_ASAP7_75t_L g5476 ( 
.A(n_5431),
.B(n_3708),
.C(n_3709),
.Y(n_5476)
);

NOR3xp33_ASAP7_75t_L g5477 ( 
.A(n_5435),
.B(n_3709),
.C(n_3696),
.Y(n_5477)
);

NAND4xp25_ASAP7_75t_SL g5478 ( 
.A(n_5429),
.B(n_3709),
.C(n_3689),
.D(n_3670),
.Y(n_5478)
);

OAI211xp5_ASAP7_75t_SL g5479 ( 
.A1(n_5425),
.A2(n_3714),
.B(n_3670),
.C(n_3689),
.Y(n_5479)
);

NOR3x1_ASAP7_75t_L g5480 ( 
.A(n_5438),
.B(n_3892),
.C(n_3861),
.Y(n_5480)
);

NOR2x1_ASAP7_75t_L g5481 ( 
.A(n_5424),
.B(n_3847),
.Y(n_5481)
);

O2A1O1Ixp33_ASAP7_75t_L g5482 ( 
.A1(n_5443),
.A2(n_5425),
.B(n_3724),
.C(n_3773),
.Y(n_5482)
);

NAND2xp5_ASAP7_75t_SL g5483 ( 
.A(n_5474),
.B(n_3670),
.Y(n_5483)
);

INVx2_ASAP7_75t_L g5484 ( 
.A(n_5480),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_SL g5485 ( 
.A(n_5450),
.B(n_3690),
.Y(n_5485)
);

INVx1_ASAP7_75t_L g5486 ( 
.A(n_5481),
.Y(n_5486)
);

NOR3xp33_ASAP7_75t_L g5487 ( 
.A(n_5444),
.B(n_5441),
.C(n_5440),
.Y(n_5487)
);

NOR2x1_ASAP7_75t_L g5488 ( 
.A(n_5470),
.B(n_3847),
.Y(n_5488)
);

AND4x1_ASAP7_75t_L g5489 ( 
.A(n_5442),
.B(n_3883),
.C(n_3886),
.D(n_3912),
.Y(n_5489)
);

NAND4xp25_ASAP7_75t_L g5490 ( 
.A(n_5459),
.B(n_3775),
.C(n_3705),
.D(n_3846),
.Y(n_5490)
);

NOR2x1p5_ASAP7_75t_L g5491 ( 
.A(n_5448),
.B(n_3714),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5472),
.Y(n_5492)
);

AOI221xp5_ASAP7_75t_L g5493 ( 
.A1(n_5451),
.A2(n_3714),
.B1(n_3738),
.B2(n_3739),
.C(n_3773),
.Y(n_5493)
);

NOR3xp33_ASAP7_75t_L g5494 ( 
.A(n_5468),
.B(n_3724),
.C(n_3739),
.Y(n_5494)
);

NOR2x1p5_ASAP7_75t_L g5495 ( 
.A(n_5455),
.B(n_3724),
.Y(n_5495)
);

NAND2xp5_ASAP7_75t_L g5496 ( 
.A(n_5473),
.B(n_5452),
.Y(n_5496)
);

NOR4xp25_ASAP7_75t_L g5497 ( 
.A(n_5445),
.B(n_3776),
.C(n_3846),
.D(n_3778),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_5447),
.Y(n_5498)
);

INVx1_ASAP7_75t_L g5499 ( 
.A(n_5462),
.Y(n_5499)
);

AOI221xp5_ASAP7_75t_L g5500 ( 
.A1(n_5453),
.A2(n_5464),
.B1(n_5471),
.B2(n_5467),
.C(n_5454),
.Y(n_5500)
);

NAND2xp5_ASAP7_75t_L g5501 ( 
.A(n_5456),
.B(n_3861),
.Y(n_5501)
);

INVx1_ASAP7_75t_L g5502 ( 
.A(n_5449),
.Y(n_5502)
);

NOR4xp25_ASAP7_75t_L g5503 ( 
.A(n_5454),
.B(n_3846),
.C(n_3778),
.D(n_3783),
.Y(n_5503)
);

AND2x2_ASAP7_75t_L g5504 ( 
.A(n_5457),
.B(n_3537),
.Y(n_5504)
);

AOI211xp5_ASAP7_75t_L g5505 ( 
.A1(n_5465),
.A2(n_3776),
.B(n_3835),
.C(n_3773),
.Y(n_5505)
);

AOI211xp5_ASAP7_75t_L g5506 ( 
.A1(n_5479),
.A2(n_3776),
.B(n_3810),
.C(n_3835),
.Y(n_5506)
);

NAND3x1_ASAP7_75t_L g5507 ( 
.A(n_5458),
.B(n_3875),
.C(n_3866),
.Y(n_5507)
);

AOI221xp5_ASAP7_75t_L g5508 ( 
.A1(n_5461),
.A2(n_3739),
.B1(n_3778),
.B2(n_3783),
.C(n_3784),
.Y(n_5508)
);

AOI221x1_ASAP7_75t_L g5509 ( 
.A1(n_5477),
.A2(n_3868),
.B1(n_3922),
.B2(n_3867),
.C(n_3888),
.Y(n_5509)
);

OAI211xp5_ASAP7_75t_L g5510 ( 
.A1(n_5466),
.A2(n_5463),
.B(n_5460),
.C(n_5476),
.Y(n_5510)
);

NOR2x1_ASAP7_75t_L g5511 ( 
.A(n_5478),
.B(n_3863),
.Y(n_5511)
);

NOR2x1_ASAP7_75t_L g5512 ( 
.A(n_5469),
.B(n_3863),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5475),
.Y(n_5513)
);

NOR3xp33_ASAP7_75t_L g5514 ( 
.A(n_5446),
.B(n_3738),
.C(n_3783),
.Y(n_5514)
);

NAND3xp33_ASAP7_75t_L g5515 ( 
.A(n_5443),
.B(n_3816),
.C(n_3789),
.Y(n_5515)
);

INVx1_ASAP7_75t_L g5516 ( 
.A(n_5474),
.Y(n_5516)
);

OAI22xp33_ASAP7_75t_L g5517 ( 
.A1(n_5450),
.A2(n_3803),
.B1(n_3810),
.B2(n_3816),
.Y(n_5517)
);

AOI22xp5_ASAP7_75t_L g5518 ( 
.A1(n_5444),
.A2(n_3784),
.B1(n_3789),
.B2(n_3803),
.Y(n_5518)
);

NAND3xp33_ASAP7_75t_L g5519 ( 
.A(n_5443),
.B(n_3816),
.C(n_3789),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5504),
.Y(n_5520)
);

NOR2xp67_ASAP7_75t_SL g5521 ( 
.A(n_5516),
.B(n_3866),
.Y(n_5521)
);

AOI21xp5_ASAP7_75t_L g5522 ( 
.A1(n_5496),
.A2(n_3803),
.B(n_3810),
.Y(n_5522)
);

AOI221x1_ASAP7_75t_L g5523 ( 
.A1(n_5487),
.A2(n_3888),
.B1(n_3922),
.B2(n_3897),
.C(n_3868),
.Y(n_5523)
);

HB1xp67_ASAP7_75t_L g5524 ( 
.A(n_5491),
.Y(n_5524)
);

AOI22xp5_ASAP7_75t_L g5525 ( 
.A1(n_5513),
.A2(n_3835),
.B1(n_3827),
.B2(n_3738),
.Y(n_5525)
);

AOI221xp5_ASAP7_75t_L g5526 ( 
.A1(n_5497),
.A2(n_3827),
.B1(n_3826),
.B2(n_3824),
.C(n_3784),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_5488),
.Y(n_5527)
);

AOI222xp33_ASAP7_75t_L g5528 ( 
.A1(n_5500),
.A2(n_3824),
.B1(n_3827),
.B2(n_3826),
.C1(n_3922),
.C2(n_3867),
.Y(n_5528)
);

INVx2_ASAP7_75t_L g5529 ( 
.A(n_5495),
.Y(n_5529)
);

OAI21xp33_ASAP7_75t_L g5530 ( 
.A1(n_5518),
.A2(n_5492),
.B(n_5490),
.Y(n_5530)
);

BUFx6f_ASAP7_75t_L g5531 ( 
.A(n_5498),
.Y(n_5531)
);

NAND2xp5_ASAP7_75t_L g5532 ( 
.A(n_5486),
.B(n_3875),
.Y(n_5532)
);

AND2x2_ASAP7_75t_L g5533 ( 
.A(n_5484),
.B(n_5502),
.Y(n_5533)
);

AND2x4_ASAP7_75t_L g5534 ( 
.A(n_5485),
.B(n_3824),
.Y(n_5534)
);

AOI21xp5_ASAP7_75t_L g5535 ( 
.A1(n_5510),
.A2(n_3826),
.B(n_3853),
.Y(n_5535)
);

INVx1_ASAP7_75t_SL g5536 ( 
.A(n_5483),
.Y(n_5536)
);

NAND4xp25_ASAP7_75t_L g5537 ( 
.A(n_5482),
.B(n_3452),
.C(n_3381),
.D(n_3888),
.Y(n_5537)
);

AOI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5494),
.A2(n_3867),
.B1(n_3868),
.B2(n_3897),
.Y(n_5538)
);

NAND2xp5_ASAP7_75t_SL g5539 ( 
.A(n_5515),
.B(n_5519),
.Y(n_5539)
);

NAND3xp33_ASAP7_75t_SL g5540 ( 
.A(n_5489),
.B(n_3897),
.C(n_3912),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5501),
.Y(n_5541)
);

NAND2xp5_ASAP7_75t_L g5542 ( 
.A(n_5511),
.B(n_3886),
.Y(n_5542)
);

AOI322xp5_ASAP7_75t_L g5543 ( 
.A1(n_5499),
.A2(n_3935),
.A3(n_3910),
.B1(n_3907),
.B2(n_3901),
.C1(n_3899),
.C2(n_3892),
.Y(n_5543)
);

OAI211xp5_ASAP7_75t_L g5544 ( 
.A1(n_5512),
.A2(n_3907),
.B(n_3890),
.C(n_3853),
.Y(n_5544)
);

NOR2xp33_ASAP7_75t_L g5545 ( 
.A(n_5517),
.B(n_3890),
.Y(n_5545)
);

AOI21xp5_ASAP7_75t_L g5546 ( 
.A1(n_5503),
.A2(n_3860),
.B(n_3853),
.Y(n_5546)
);

AOI211xp5_ASAP7_75t_L g5547 ( 
.A1(n_5514),
.A2(n_3452),
.B(n_3935),
.C(n_3833),
.Y(n_5547)
);

OAI22xp33_ASAP7_75t_L g5548 ( 
.A1(n_5509),
.A2(n_3935),
.B1(n_3860),
.B2(n_3628),
.Y(n_5548)
);

NAND3xp33_ASAP7_75t_L g5549 ( 
.A(n_5505),
.B(n_5506),
.C(n_5493),
.Y(n_5549)
);

INVx1_ASAP7_75t_L g5550 ( 
.A(n_5542),
.Y(n_5550)
);

NAND2xp5_ASAP7_75t_L g5551 ( 
.A(n_5520),
.B(n_5507),
.Y(n_5551)
);

OAI22xp5_ASAP7_75t_L g5552 ( 
.A1(n_5525),
.A2(n_5505),
.B1(n_5506),
.B2(n_5508),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5521),
.Y(n_5553)
);

INVx1_ASAP7_75t_L g5554 ( 
.A(n_5524),
.Y(n_5554)
);

AND2x4_ASAP7_75t_L g5555 ( 
.A(n_5527),
.B(n_3540),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5532),
.Y(n_5556)
);

XOR2xp5_ASAP7_75t_L g5557 ( 
.A(n_5549),
.B(n_3833),
.Y(n_5557)
);

NAND2xp5_ASAP7_75t_L g5558 ( 
.A(n_5547),
.B(n_3550),
.Y(n_5558)
);

NOR2x1_ASAP7_75t_L g5559 ( 
.A(n_5529),
.B(n_3860),
.Y(n_5559)
);

XOR2xp5_ASAP7_75t_L g5560 ( 
.A(n_5533),
.B(n_3477),
.Y(n_5560)
);

NOR2xp67_ASAP7_75t_L g5561 ( 
.A(n_5540),
.B(n_3628),
.Y(n_5561)
);

AND2x4_ASAP7_75t_L g5562 ( 
.A(n_5536),
.B(n_5531),
.Y(n_5562)
);

NOR2x1p5_ASAP7_75t_L g5563 ( 
.A(n_5531),
.B(n_3628),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_5531),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_5530),
.B(n_3550),
.Y(n_5565)
);

INVx2_ASAP7_75t_SL g5566 ( 
.A(n_5534),
.Y(n_5566)
);

INVx2_ASAP7_75t_L g5567 ( 
.A(n_5534),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_5539),
.Y(n_5568)
);

INVxp33_ASAP7_75t_L g5569 ( 
.A(n_5541),
.Y(n_5569)
);

NOR2xp33_ASAP7_75t_L g5570 ( 
.A(n_5537),
.B(n_3860),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_L g5571 ( 
.A(n_5555),
.B(n_5545),
.Y(n_5571)
);

AND2x4_ASAP7_75t_L g5572 ( 
.A(n_5563),
.B(n_5522),
.Y(n_5572)
);

NOR3xp33_ASAP7_75t_SL g5573 ( 
.A(n_5551),
.B(n_5544),
.C(n_5535),
.Y(n_5573)
);

NAND3x2_ASAP7_75t_L g5574 ( 
.A(n_5562),
.B(n_5523),
.C(n_5543),
.Y(n_5574)
);

NOR3xp33_ASAP7_75t_L g5575 ( 
.A(n_5554),
.B(n_5546),
.C(n_5548),
.Y(n_5575)
);

NAND2x1p5_ASAP7_75t_L g5576 ( 
.A(n_5562),
.B(n_5538),
.Y(n_5576)
);

NOR3xp33_ASAP7_75t_L g5577 ( 
.A(n_5568),
.B(n_5526),
.C(n_5528),
.Y(n_5577)
);

NOR2x2_ASAP7_75t_L g5578 ( 
.A(n_5567),
.B(n_5560),
.Y(n_5578)
);

NOR2xp33_ASAP7_75t_L g5579 ( 
.A(n_5555),
.B(n_3742),
.Y(n_5579)
);

NAND3x1_ASAP7_75t_L g5580 ( 
.A(n_5564),
.B(n_5553),
.C(n_5550),
.Y(n_5580)
);

NAND3xp33_ASAP7_75t_L g5581 ( 
.A(n_5556),
.B(n_3742),
.C(n_3735),
.Y(n_5581)
);

NOR4xp75_ASAP7_75t_L g5582 ( 
.A(n_5552),
.B(n_3469),
.C(n_3458),
.D(n_3456),
.Y(n_5582)
);

XNOR2xp5_ASAP7_75t_L g5583 ( 
.A(n_5557),
.B(n_3424),
.Y(n_5583)
);

OAI22xp5_ASAP7_75t_L g5584 ( 
.A1(n_5565),
.A2(n_3364),
.B1(n_3377),
.B2(n_3626),
.Y(n_5584)
);

OR2x2_ASAP7_75t_L g5585 ( 
.A(n_5558),
.B(n_3550),
.Y(n_5585)
);

NOR3xp33_ASAP7_75t_SL g5586 ( 
.A(n_5570),
.B(n_3657),
.C(n_3627),
.Y(n_5586)
);

INVx2_ASAP7_75t_L g5587 ( 
.A(n_5583),
.Y(n_5587)
);

NOR2xp33_ASAP7_75t_L g5588 ( 
.A(n_5571),
.B(n_5569),
.Y(n_5588)
);

CKINVDCx5p33_ASAP7_75t_R g5589 ( 
.A(n_5573),
.Y(n_5589)
);

CKINVDCx5p33_ASAP7_75t_R g5590 ( 
.A(n_5572),
.Y(n_5590)
);

HB1xp67_ASAP7_75t_L g5591 ( 
.A(n_5572),
.Y(n_5591)
);

NOR2x1p5_ASAP7_75t_L g5592 ( 
.A(n_5585),
.B(n_5566),
.Y(n_5592)
);

INVx2_ASAP7_75t_L g5593 ( 
.A(n_5578),
.Y(n_5593)
);

OAI221xp5_ASAP7_75t_L g5594 ( 
.A1(n_5575),
.A2(n_5559),
.B1(n_5561),
.B2(n_3742),
.C(n_3735),
.Y(n_5594)
);

INVx1_ASAP7_75t_SL g5595 ( 
.A(n_5580),
.Y(n_5595)
);

BUFx2_ASAP7_75t_L g5596 ( 
.A(n_5574),
.Y(n_5596)
);

CKINVDCx20_ASAP7_75t_R g5597 ( 
.A(n_5577),
.Y(n_5597)
);

OAI211xp5_ASAP7_75t_SL g5598 ( 
.A1(n_5595),
.A2(n_5576),
.B(n_5586),
.C(n_5584),
.Y(n_5598)
);

AOI322xp5_ASAP7_75t_L g5599 ( 
.A1(n_5588),
.A2(n_5579),
.A3(n_5582),
.B1(n_5581),
.B2(n_3480),
.C1(n_3448),
.C2(n_3414),
.Y(n_5599)
);

INVx1_ASAP7_75t_L g5600 ( 
.A(n_5591),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5596),
.B(n_3742),
.Y(n_5601)
);

AOI322xp5_ASAP7_75t_L g5602 ( 
.A1(n_5593),
.A2(n_3480),
.A3(n_3448),
.B1(n_3437),
.B2(n_3414),
.C1(n_3424),
.C2(n_3377),
.Y(n_5602)
);

NOR3xp33_ASAP7_75t_L g5603 ( 
.A(n_5589),
.B(n_3364),
.C(n_3540),
.Y(n_5603)
);

OAI22xp5_ASAP7_75t_L g5604 ( 
.A1(n_5597),
.A2(n_3735),
.B1(n_3663),
.B2(n_3626),
.Y(n_5604)
);

AOI322xp5_ASAP7_75t_L g5605 ( 
.A1(n_5587),
.A2(n_3480),
.A3(n_3437),
.B1(n_3491),
.B2(n_3458),
.C1(n_3456),
.C2(n_3468),
.Y(n_5605)
);

OAI211xp5_ASAP7_75t_SL g5606 ( 
.A1(n_5592),
.A2(n_3550),
.B(n_3367),
.C(n_3391),
.Y(n_5606)
);

AO22x2_ASAP7_75t_L g5607 ( 
.A1(n_5600),
.A2(n_5590),
.B1(n_5594),
.B2(n_3468),
.Y(n_5607)
);

AOI22xp5_ASAP7_75t_L g5608 ( 
.A1(n_5598),
.A2(n_3735),
.B1(n_3454),
.B2(n_3597),
.Y(n_5608)
);

HB1xp67_ASAP7_75t_L g5609 ( 
.A(n_5601),
.Y(n_5609)
);

AOI22xp5_ASAP7_75t_L g5610 ( 
.A1(n_5603),
.A2(n_3454),
.B1(n_3597),
.B2(n_3556),
.Y(n_5610)
);

OAI22xp5_ASAP7_75t_L g5611 ( 
.A1(n_5604),
.A2(n_3537),
.B1(n_3663),
.B2(n_3600),
.Y(n_5611)
);

NOR3xp33_ASAP7_75t_L g5612 ( 
.A(n_5609),
.B(n_5607),
.C(n_5608),
.Y(n_5612)
);

NAND4xp25_ASAP7_75t_SL g5613 ( 
.A(n_5610),
.B(n_5599),
.C(n_5602),
.D(n_5605),
.Y(n_5613)
);

NOR3xp33_ASAP7_75t_SL g5614 ( 
.A(n_5611),
.B(n_5606),
.C(n_3652),
.Y(n_5614)
);

AOI21xp5_ASAP7_75t_SL g5615 ( 
.A1(n_5613),
.A2(n_3480),
.B(n_3499),
.Y(n_5615)
);

AO21x1_ASAP7_75t_L g5616 ( 
.A1(n_5615),
.A2(n_5612),
.B(n_5614),
.Y(n_5616)
);

OAI22xp5_ASAP7_75t_L g5617 ( 
.A1(n_5616),
.A2(n_3587),
.B1(n_3556),
.B2(n_3624),
.Y(n_5617)
);

AOI21xp5_ASAP7_75t_L g5618 ( 
.A1(n_5617),
.A2(n_3624),
.B(n_3499),
.Y(n_5618)
);

AOI22xp5_ASAP7_75t_L g5619 ( 
.A1(n_5618),
.A2(n_3485),
.B1(n_3491),
.B2(n_3502),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_SL g5620 ( 
.A(n_5619),
.B(n_3491),
.Y(n_5620)
);

BUFx2_ASAP7_75t_SL g5621 ( 
.A(n_5620),
.Y(n_5621)
);

AOI221xp5_ASAP7_75t_L g5622 ( 
.A1(n_5621),
.A2(n_3485),
.B1(n_3491),
.B2(n_3502),
.C(n_3504),
.Y(n_5622)
);

AOI21xp5_ASAP7_75t_L g5623 ( 
.A1(n_5622),
.A2(n_3366),
.B(n_3367),
.Y(n_5623)
);

AOI211xp5_ASAP7_75t_L g5624 ( 
.A1(n_5623),
.A2(n_3391),
.B(n_3592),
.C(n_3504),
.Y(n_5624)
);


endmodule