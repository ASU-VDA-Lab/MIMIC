module fake_jpeg_3778_n_59 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_56;
wire n_31;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_4),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_22),
.A2(n_34),
.B1(n_18),
.B2(n_20),
.Y(n_39)
);

AO21x2_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_22),
.A2(n_17),
.B1(n_18),
.B2(n_20),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_30),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_26),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_17),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_48),
.A2(n_45),
.B(n_42),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_48),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_48),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_51),
.A2(n_52),
.B1(n_42),
.B2(n_46),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_53),
.B(n_54),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_43),
.B(n_47),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_56),
.A2(n_37),
.B(n_44),
.C(n_32),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g58 ( 
.A(n_57),
.B(n_55),
.C(n_21),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_31),
.Y(n_59)
);


endmodule