module fake_netlist_6_3190_n_1619 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1619);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1619;

wire n_992;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_163;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_148;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_147;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_153;
wire n_842;
wire n_1432;
wire n_156;
wire n_145;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_154;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_150;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_146;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_144;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_152;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_151;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_149;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_6),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_121),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g146 ( 
.A(n_74),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_67),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_12),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_38),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_17),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_66),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_41),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_143),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_60),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_52),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_59),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_62),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_96),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_88),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_84),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_70),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_65),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_53),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_35),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_23),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_47),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_37),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_46),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_31),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_135),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_137),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_109),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_22),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_49),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_15),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_39),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_85),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_61),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_57),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_117),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_4),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_16),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_42),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_32),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_69),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_118),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_139),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_71),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_123),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_9),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_58),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_119),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_29),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_93),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_83),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_46),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_10),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_76),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_44),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_1),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_81),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_129),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_106),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_134),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_77),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_111),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_17),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_108),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_24),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_27),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_142),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_41),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_13),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_18),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_12),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_127),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_72),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_20),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_79),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_49),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_132),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_122),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_26),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_7),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_75),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_45),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_73),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_114),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_13),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_22),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_103),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_32),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_136),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_97),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_48),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_124),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_28),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_39),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_107),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_36),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_33),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_24),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_34),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_28),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_140),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_68),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_101),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_47),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_43),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_92),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_113),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_63),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_112),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_42),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_10),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_37),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_145),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_147),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_149),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_157),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_158),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_189),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_152),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_274),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_274),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_274),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_206),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_206),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_197),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_198),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_221),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_224),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_278),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_160),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_161),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_156),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_224),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_198),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_268),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_268),
.Y(n_315)
);

BUFx2_ASAP7_75t_SL g316 ( 
.A(n_168),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_213),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_213),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_213),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_250),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

INVx2_ASAP7_75t_SL g322 ( 
.A(n_250),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_162),
.Y(n_323)
);

INVxp33_ASAP7_75t_SL g324 ( 
.A(n_144),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_154),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_154),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_237),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_230),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_148),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_179),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_164),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_179),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_184),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_184),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_185),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_230),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_185),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_193),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_193),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_155),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_204),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_212),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_212),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_217),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_166),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_217),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_228),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_169),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_229),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_229),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_235),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_293),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_285),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_285),
.B(n_216),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_285),
.B(n_216),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_294),
.B(n_195),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_283),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_291),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_284),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_296),
.B(n_220),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g367 ( 
.A1(n_328),
.A2(n_230),
.B(n_151),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_289),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_295),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_295),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_297),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_297),
.B(n_220),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_322),
.B(n_168),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_290),
.A2(n_265),
.B1(n_247),
.B2(n_153),
.Y(n_375)
);

AOI22x1_ASAP7_75t_SL g376 ( 
.A1(n_300),
.A2(n_194),
.B1(n_281),
.B2(n_280),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_302),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_336),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_325),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

OA21x2_ASAP7_75t_L g383 ( 
.A1(n_298),
.A2(n_151),
.B(n_150),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_326),
.Y(n_384)
);

AND2x6_ASAP7_75t_L g385 ( 
.A(n_301),
.B(n_220),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_326),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_243),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_299),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_287),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_303),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_150),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_317),
.B(n_318),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_303),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_304),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_288),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_316),
.B(n_170),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_292),
.Y(n_401)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_304),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_306),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_306),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_171),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_333),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_294),
.B(n_210),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_310),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_310),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_334),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_318),
.B(n_175),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_395),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_395),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_360),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_395),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_353),
.B(n_307),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_362),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_367),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_360),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_353),
.B(n_308),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_402),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_394),
.B(n_319),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_356),
.B(n_340),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_366),
.B(n_319),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_367),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_352),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_362),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_357),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_356),
.B(n_340),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_400),
.B(n_324),
.Y(n_440)
);

AND3x2_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_163),
.C(n_159),
.Y(n_441)
);

INVx2_ASAP7_75t_SL g442 ( 
.A(n_402),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

AOI21x1_ASAP7_75t_L g445 ( 
.A1(n_358),
.A2(n_314),
.B(n_311),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_353),
.B(n_323),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

BUFx10_ASAP7_75t_L g450 ( 
.A(n_361),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_400),
.B(n_331),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_R g452 ( 
.A(n_363),
.B(n_391),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_359),
.B(n_345),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_359),
.B(n_348),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_365),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_362),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_368),
.Y(n_461)
);

BUFx8_ASAP7_75t_SL g462 ( 
.A(n_352),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_379),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_402),
.B(n_327),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_409),
.B(n_181),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_379),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g469 ( 
.A(n_412),
.B(n_178),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_362),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_354),
.B(n_309),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_394),
.B(n_320),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_402),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_362),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_381),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_399),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_359),
.B(n_313),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_409),
.B(n_320),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_381),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_402),
.B(n_390),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_390),
.B(n_165),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_370),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_377),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_355),
.B(n_321),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_416),
.B(n_199),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_369),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_371),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_369),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_401),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_377),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_394),
.B(n_355),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_371),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_369),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_378),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_L g499 ( 
.A1(n_372),
.A2(n_245),
.B1(n_251),
.B2(n_256),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_377),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_404),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_416),
.B(n_321),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_404),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_378),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_387),
.B(n_334),
.Y(n_507)
);

OR2x6_ASAP7_75t_L g508 ( 
.A(n_387),
.B(n_245),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_366),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

NAND2xp33_ASAP7_75t_L g511 ( 
.A(n_385),
.B(n_182),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_R g512 ( 
.A(n_376),
.B(n_172),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_373),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_372),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_373),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_380),
.Y(n_517)
);

AOI21x1_ASAP7_75t_L g518 ( 
.A1(n_383),
.A2(n_314),
.B(n_311),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_380),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_366),
.B(n_315),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_382),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_382),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_396),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_366),
.B(n_315),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_384),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_396),
.Y(n_529)
);

AO21x2_ASAP7_75t_L g530 ( 
.A1(n_374),
.A2(n_163),
.B(n_159),
.Y(n_530)
);

INVxp67_ASAP7_75t_SL g531 ( 
.A(n_366),
.Y(n_531)
);

NAND3xp33_ASAP7_75t_L g532 ( 
.A(n_375),
.B(n_174),
.C(n_173),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_372),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g534 ( 
.A(n_385),
.B(n_183),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_386),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_396),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_386),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_374),
.B(n_305),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_396),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_388),
.B(n_210),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_385),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_376),
.B(n_176),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_396),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_396),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_388),
.Y(n_545)
);

BUFx6f_ASAP7_75t_SL g546 ( 
.A(n_385),
.Y(n_546)
);

CKINVDCx20_ASAP7_75t_R g547 ( 
.A(n_383),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_397),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_396),
.Y(n_549)
);

INVx3_ASAP7_75t_L g550 ( 
.A(n_398),
.Y(n_550)
);

AND3x2_ASAP7_75t_L g551 ( 
.A(n_397),
.B(n_180),
.C(n_167),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_398),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_385),
.B(n_190),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_406),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_406),
.B(n_210),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_398),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_408),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_408),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_504),
.B(n_410),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_547),
.A2(n_383),
.B1(n_264),
.B2(n_235),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_471),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_494),
.B(n_385),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_507),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_521),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_494),
.B(n_385),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_482),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_479),
.B(n_385),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_452),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_417),
.A2(n_383),
.B1(n_251),
.B2(n_271),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_521),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_419),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_486),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g574 ( 
.A(n_471),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_440),
.B(n_177),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_503),
.B(n_383),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_451),
.B(n_167),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_507),
.A2(n_256),
.B(n_239),
.Y(n_579)
);

A2O1A1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_487),
.A2(n_239),
.B(n_271),
.C(n_264),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_488),
.B(n_421),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_419),
.Y(n_583)
);

INVxp33_ASAP7_75t_L g584 ( 
.A(n_462),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_437),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_482),
.B(n_191),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_509),
.B(n_180),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_527),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_482),
.B(n_200),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_485),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_531),
.B(n_188),
.Y(n_591)
);

INVx8_ASAP7_75t_L g592 ( 
.A(n_546),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_444),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_486),
.B(n_188),
.Y(n_594)
);

A2O1A1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_417),
.A2(n_261),
.B(n_248),
.C(n_263),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_486),
.B(n_219),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_219),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_427),
.B(n_186),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_418),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_482),
.B(n_202),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_493),
.B(n_222),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_425),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_482),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_533),
.B(n_514),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

NOR2x1p5_ASAP7_75t_L g607 ( 
.A(n_477),
.B(n_187),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_538),
.A2(n_146),
.B1(n_227),
.B2(n_269),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_447),
.B(n_192),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_493),
.B(n_498),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_498),
.B(n_222),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_533),
.B(n_203),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_418),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_504),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_533),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_485),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_448),
.Y(n_617)
);

AO22x2_ASAP7_75t_L g618 ( 
.A1(n_532),
.A2(n_438),
.B1(n_432),
.B2(n_542),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_425),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_420),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_501),
.B(n_240),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_506),
.B(n_248),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_420),
.A2(n_270),
.B(n_263),
.C(n_261),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_433),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_530),
.A2(n_422),
.B1(n_428),
.B2(n_424),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_433),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_483),
.B(n_196),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_533),
.B(n_207),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_533),
.B(n_208),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_433),
.B(n_411),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_514),
.B(n_211),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_431),
.B(n_411),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_477),
.B(n_415),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_506),
.B(n_270),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_431),
.B(n_415),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_513),
.B(n_398),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_513),
.B(n_398),
.Y(n_638)
);

INVx2_ASAP7_75t_SL g639 ( 
.A(n_473),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_481),
.B(n_214),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_530),
.A2(n_195),
.B1(n_205),
.B2(n_342),
.Y(n_641)
);

AOI221xp5_ASAP7_75t_L g642 ( 
.A1(n_469),
.A2(n_259),
.B1(n_253),
.B2(n_244),
.C(n_257),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_450),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_516),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_453),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_473),
.B(n_195),
.Y(n_646)
);

O2A1O1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_422),
.A2(n_347),
.B(n_337),
.C(n_338),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_455),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_508),
.B(n_195),
.Y(n_650)
);

BUFx6f_ASAP7_75t_L g651 ( 
.A(n_541),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_517),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_492),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_517),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_467),
.A2(n_223),
.B1(n_277),
.B2(n_276),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_441),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_454),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_466),
.A2(n_218),
.B1(n_275),
.B2(n_272),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_519),
.B(n_398),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_530),
.A2(n_205),
.B1(n_351),
.B2(n_350),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_554),
.B(n_519),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_492),
.B(n_233),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_508),
.B(n_205),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_524),
.B(n_403),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_528),
.B(n_403),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_508),
.B(n_205),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_535),
.B(n_403),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_541),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_L g669 ( 
.A1(n_430),
.A2(n_414),
.B(n_413),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_535),
.B(n_403),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_430),
.A2(n_434),
.B1(n_558),
.B2(n_557),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_508),
.B(n_335),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_537),
.B(n_403),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_537),
.A2(n_258),
.B1(n_238),
.B2(n_242),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_545),
.B(n_201),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_548),
.B(n_403),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_434),
.B(n_246),
.Y(n_677)
);

INVxp67_ASAP7_75t_L g678 ( 
.A(n_435),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_548),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_557),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_543),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_558),
.A2(n_511),
.B1(n_534),
.B2(n_553),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_455),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_551),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_456),
.B(n_209),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_543),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_456),
.B(n_225),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_457),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_497),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_439),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_497),
.B(n_335),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_450),
.B(n_337),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_429),
.A2(n_414),
.B(n_413),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_450),
.B(n_338),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_457),
.B(n_403),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_461),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_540),
.B(n_339),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_461),
.B(n_413),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_463),
.B(n_249),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_463),
.B(n_407),
.Y(n_700)
);

OAI22xp33_ASAP7_75t_L g701 ( 
.A1(n_555),
.A2(n_282),
.B1(n_226),
.B2(n_231),
.Y(n_701)
);

NOR3xp33_ASAP7_75t_L g702 ( 
.A(n_505),
.B(n_260),
.C(n_232),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_499),
.B(n_339),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_484),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_484),
.A2(n_342),
.B1(n_341),
.B2(n_343),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_490),
.B(n_389),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_495),
.B(n_536),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_443),
.B(n_389),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_495),
.B(n_407),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_442),
.B(n_407),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_500),
.B(n_252),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_446),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_536),
.B(n_236),
.Y(n_713)
);

OAI22xp5_ASAP7_75t_L g714 ( 
.A1(n_443),
.A2(n_255),
.B1(n_254),
.B2(n_279),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_446),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_500),
.B(n_210),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_590),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_576),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_576),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_581),
.B(n_442),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_567),
.B(n_515),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_651),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_651),
.B(n_474),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_562),
.B(n_542),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_585),
.Y(n_725)
);

AND2x4_ASAP7_75t_SL g726 ( 
.A(n_616),
.B(n_341),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_585),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_SL g728 ( 
.A(n_575),
.B(n_512),
.C(n_505),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_651),
.B(n_470),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_573),
.B(n_426),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_651),
.Y(n_731)
);

INVx6_ASAP7_75t_L g732 ( 
.A(n_590),
.Y(n_732)
);

NOR2x2_ASAP7_75t_L g733 ( 
.A(n_618),
.B(n_515),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_567),
.B(n_520),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_593),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_593),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_578),
.B(n_426),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_596),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_575),
.A2(n_343),
.B(n_344),
.C(n_346),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_596),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_574),
.B(n_344),
.Y(n_741)
);

INVx6_ASAP7_75t_L g742 ( 
.A(n_631),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_661),
.B(n_426),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_668),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_661),
.B(n_436),
.Y(n_745)
);

NOR2x2_ASAP7_75t_L g746 ( 
.A(n_618),
.B(n_520),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_569),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_561),
.A2(n_546),
.B1(n_472),
.B2(n_476),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_561),
.A2(n_570),
.B1(n_613),
.B2(n_600),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_617),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_653),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_620),
.B(n_628),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_628),
.B(n_436),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_649),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_565),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_582),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_633),
.B(n_436),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_668),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_346),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_567),
.B(n_522),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_636),
.B(n_644),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_668),
.B(n_546),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_572),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_571),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_691),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_606),
.Y(n_768)
);

AND2x6_ASAP7_75t_SL g769 ( 
.A(n_599),
.B(n_347),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_648),
.B(n_449),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_668),
.B(n_470),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_631),
.B(n_349),
.Y(n_772)
);

INVx5_ASAP7_75t_L g773 ( 
.A(n_592),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_689),
.A2(n_241),
.B1(n_262),
.B2(n_266),
.Y(n_774)
);

NOR3xp33_ASAP7_75t_L g775 ( 
.A(n_645),
.B(n_267),
.C(n_273),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_583),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_643),
.Y(n_777)
);

AND2x6_ASAP7_75t_SL g778 ( 
.A(n_599),
.B(n_349),
.Y(n_778)
);

AND3x2_ASAP7_75t_SL g779 ( 
.A(n_618),
.B(n_0),
.C(n_1),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_564),
.B(n_449),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_692),
.B(n_350),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_643),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_603),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_669),
.A2(n_470),
.B(n_559),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_570),
.A2(n_468),
.B1(n_480),
.B2(n_476),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_567),
.B(n_522),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_694),
.B(n_351),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_588),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_604),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_625),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_652),
.B(n_449),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_654),
.B(n_460),
.Y(n_792)
);

INVx1_ASAP7_75t_SL g793 ( 
.A(n_560),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_627),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_614),
.Y(n_795)
);

AND2x6_ASAP7_75t_SL g796 ( 
.A(n_609),
.B(n_2),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_460),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_619),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_657),
.B(n_460),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_626),
.A2(n_525),
.B1(n_556),
.B2(n_523),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_672),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_646),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_679),
.B(n_536),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_680),
.B(n_550),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_683),
.B(n_550),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_688),
.B(n_550),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_650),
.Y(n_807)
);

AOI22xp5_ASAP7_75t_L g808 ( 
.A1(n_609),
.A2(n_523),
.B1(n_556),
.B2(n_525),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_696),
.B(n_526),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_704),
.B(n_526),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_697),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_663),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_604),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_698),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_671),
.B(n_529),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_610),
.A2(n_470),
.B(n_552),
.Y(n_816)
);

INVxp67_ASAP7_75t_SL g817 ( 
.A(n_604),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_SL g818 ( 
.A(n_607),
.B(n_470),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_R g819 ( 
.A(n_592),
.B(n_656),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_604),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_700),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_678),
.B(n_464),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_563),
.A2(n_539),
.B1(n_529),
.B2(n_549),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_671),
.B(n_539),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_706),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_684),
.Y(n_826)
);

BUFx12f_ASAP7_75t_L g827 ( 
.A(n_666),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_690),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_712),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_675),
.B(n_544),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_566),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_675),
.B(n_549),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_615),
.B(n_543),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_592),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_634),
.B(n_464),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_708),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_685),
.B(n_465),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_647),
.A2(n_580),
.B(n_595),
.C(n_624),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_709),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_626),
.A2(n_472),
.B1(n_480),
.B2(n_468),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_632),
.A2(n_489),
.B1(n_491),
.B2(n_496),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_632),
.A2(n_640),
.B1(n_677),
.B2(n_612),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_685),
.B(n_465),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_715),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_615),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_681),
.Y(n_846)
);

AND3x2_ASAP7_75t_SL g847 ( 
.A(n_641),
.B(n_580),
.C(n_660),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_687),
.B(n_707),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_637),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_638),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_703),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_687),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_608),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_587),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_664),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_707),
.B(n_489),
.Y(n_857)
);

NOR2xp67_ASAP7_75t_L g858 ( 
.A(n_662),
.B(n_518),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_605),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_708),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_640),
.A2(n_496),
.B1(n_491),
.B2(n_559),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_568),
.B(n_552),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_699),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_591),
.B(n_459),
.Y(n_864)
);

NOR3xp33_ASAP7_75t_SL g865 ( 
.A(n_701),
.B(n_2),
.C(n_3),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_699),
.B(n_458),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_665),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_595),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_577),
.B(n_552),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_702),
.B(n_518),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_605),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_586),
.B(n_559),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_713),
.B(n_660),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_682),
.B(n_552),
.Y(n_874)
);

AND2x6_ASAP7_75t_L g875 ( 
.A(n_594),
.B(n_597),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_641),
.A2(n_459),
.B1(n_392),
.B2(n_393),
.Y(n_876)
);

BUFx4f_ASAP7_75t_L g877 ( 
.A(n_584),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_667),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_586),
.B(n_559),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_579),
.A2(n_392),
.B1(n_393),
.B2(n_405),
.Y(n_880)
);

NOR2x2_ASAP7_75t_L g881 ( 
.A(n_642),
.B(n_4),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_716),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_705),
.B(n_392),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_677),
.A2(n_559),
.B1(n_552),
.B2(n_543),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_670),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_L g886 ( 
.A1(n_611),
.A2(n_405),
.B1(n_393),
.B2(n_543),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_673),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_676),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_695),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_621),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_852),
.A2(n_716),
.B(n_624),
.C(n_589),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_727),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_873),
.A2(n_630),
.B1(n_589),
.B2(n_629),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_754),
.B(n_674),
.Y(n_894)
);

AOI21x1_ASAP7_75t_L g895 ( 
.A1(n_869),
.A2(n_635),
.B(n_623),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_848),
.B(n_602),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_749),
.A2(n_598),
.B1(n_612),
.B2(n_629),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_760),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_767),
.B(n_714),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_732),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_729),
.A2(n_693),
.B(n_681),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_890),
.B(n_814),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_756),
.Y(n_903)
);

INVx4_ASAP7_75t_L g904 ( 
.A(n_732),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_771),
.A2(n_686),
.B(n_601),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_821),
.B(n_630),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_869),
.A2(n_862),
.B(n_874),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_825),
.B(n_601),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_756),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_842),
.A2(n_710),
.B(n_711),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_853),
.B(n_658),
.C(n_655),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_851),
.B(n_711),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_732),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_758),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_839),
.B(n_405),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_718),
.Y(n_916)
);

INVx4_ASAP7_75t_L g917 ( 
.A(n_760),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_760),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_749),
.A2(n_445),
.B1(n_475),
.B2(n_423),
.Y(n_919)
);

NAND3xp33_ASAP7_75t_L g920 ( 
.A(n_775),
.B(n_863),
.C(n_724),
.Y(n_920)
);

OAI22xp33_ASAP7_75t_L g921 ( 
.A1(n_802),
.A2(n_445),
.B1(n_510),
.B2(n_475),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_738),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_811),
.B(n_510),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_855),
.B(n_9),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_760),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_758),
.B(n_11),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_801),
.B(n_763),
.Y(n_927)
);

OAI21xp33_ASAP7_75t_L g928 ( 
.A1(n_781),
.A2(n_11),
.B(n_14),
.Y(n_928)
);

HB1xp67_ASAP7_75t_L g929 ( 
.A(n_768),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_855),
.B(n_475),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_768),
.B(n_15),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_831),
.B(n_475),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_845),
.A2(n_510),
.B(n_475),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_787),
.B(n_510),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_R g935 ( 
.A(n_751),
.B(n_64),
.Y(n_935)
);

OAI22xp5_ASAP7_75t_L g936 ( 
.A1(n_720),
.A2(n_475),
.B1(n_423),
.B2(n_510),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_845),
.A2(n_510),
.B(n_423),
.Y(n_937)
);

XOR2xp5_ASAP7_75t_L g938 ( 
.A(n_747),
.B(n_56),
.Y(n_938)
);

O2A1O1Ixp5_ASAP7_75t_SL g939 ( 
.A1(n_874),
.A2(n_19),
.B(n_21),
.C(n_25),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_831),
.B(n_423),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_887),
.B(n_423),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_846),
.A2(n_423),
.B(n_78),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_887),
.B(n_55),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_795),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_849),
.B(n_54),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_788),
.B(n_80),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_719),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_870),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_725),
.Y(n_949)
);

AO32x1_ASAP7_75t_L g950 ( 
.A1(n_800),
.A2(n_840),
.A3(n_884),
.B1(n_882),
.B2(n_735),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_850),
.B(n_87),
.Y(n_951)
);

AOI21x1_ASAP7_75t_L g952 ( 
.A1(n_862),
.A2(n_86),
.B(n_138),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_854),
.B(n_50),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_788),
.B(n_90),
.Y(n_954)
);

BUFx12f_ASAP7_75t_L g955 ( 
.A(n_827),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_736),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_755),
.A2(n_91),
.B(n_126),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_740),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_R g959 ( 
.A(n_818),
.B(n_141),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_722),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_739),
.A2(n_30),
.B(n_33),
.C(n_35),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_857),
.A2(n_94),
.B(n_104),
.Y(n_962)
);

BUFx2_ASAP7_75t_L g963 ( 
.A(n_717),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_795),
.B(n_30),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_757),
.B(n_766),
.Y(n_965)
);

INVxp67_ASAP7_75t_L g966 ( 
.A(n_741),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_807),
.B(n_36),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_812),
.A2(n_95),
.B1(n_100),
.B2(n_99),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_877),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_856),
.B(n_885),
.Y(n_970)
);

AO31x2_ASAP7_75t_L g971 ( 
.A1(n_739),
.A2(n_38),
.A3(n_40),
.B(n_43),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_748),
.A2(n_98),
.B1(n_125),
.B2(n_45),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_784),
.A2(n_40),
.B(n_44),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_724),
.B(n_775),
.C(n_774),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_794),
.B(n_772),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_726),
.B(n_772),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_794),
.B(n_761),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_761),
.B(n_822),
.Y(n_978)
);

INVx3_ASAP7_75t_SL g979 ( 
.A(n_881),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_726),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_773),
.B(n_835),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_737),
.A2(n_745),
.B(n_743),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_888),
.B(n_889),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_769),
.B(n_778),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_864),
.A2(n_830),
.B(n_730),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_834),
.B(n_777),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_742),
.B(n_826),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_L g988 ( 
.A1(n_832),
.A2(n_837),
.B(n_843),
.C(n_734),
.Y(n_988)
);

O2A1O1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_815),
.A2(n_824),
.B(n_786),
.C(n_721),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_816),
.A2(n_759),
.B(n_817),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_773),
.B(n_790),
.Y(n_991)
);

O2A1O1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_865),
.A2(n_799),
.B(n_797),
.C(n_838),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_750),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_817),
.A2(n_858),
.B(n_748),
.Y(n_994)
);

NOR3xp33_ASAP7_75t_SL g995 ( 
.A(n_779),
.B(n_797),
.C(n_746),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_773),
.B(n_820),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_742),
.B(n_782),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_773),
.B(n_820),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_832),
.A2(n_859),
.B(n_871),
.C(n_868),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_833),
.A2(n_859),
.B(n_871),
.Y(n_1000)
);

NAND2xp33_ASAP7_75t_L g1001 ( 
.A(n_764),
.B(n_860),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_722),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_866),
.A2(n_780),
.B(n_752),
.C(n_753),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_780),
.A2(n_728),
.B(n_810),
.C(n_809),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_733),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_834),
.B(n_836),
.Y(n_1006)
);

NOR2x1_ASAP7_75t_R g1007 ( 
.A(n_779),
.B(n_836),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_728),
.A2(n_806),
.B(n_803),
.C(n_804),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_833),
.A2(n_872),
.B(n_879),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_860),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_731),
.A2(n_744),
.B1(n_879),
.B2(n_872),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_721),
.A2(n_762),
.B(n_786),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_867),
.B(n_878),
.Y(n_1013)
);

INVx6_ASAP7_75t_L g1014 ( 
.A(n_860),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_877),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_883),
.B(n_819),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_734),
.A2(n_762),
.B(n_792),
.C(n_791),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_765),
.Y(n_1018)
);

OR2x2_ASAP7_75t_L g1019 ( 
.A(n_783),
.B(n_828),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_765),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_819),
.B(n_828),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_789),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_SL g1023 ( 
.A1(n_796),
.A2(n_847),
.B1(n_860),
.B2(n_723),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_985),
.A2(n_723),
.B(n_770),
.Y(n_1024)
);

CKINVDCx16_ASAP7_75t_R g1025 ( 
.A(n_969),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_966),
.B(n_844),
.Y(n_1026)
);

AO32x2_ASAP7_75t_L g1027 ( 
.A1(n_1023),
.A2(n_847),
.A3(n_876),
.B1(n_875),
.B2(n_808),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_929),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_976),
.B(n_1016),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_SL g1030 ( 
.A1(n_928),
.A2(n_876),
.B1(n_880),
.B2(n_805),
.C(n_785),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_992),
.A2(n_823),
.B(n_841),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_920),
.B(n_844),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_909),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_894),
.A2(n_861),
.B(n_776),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_902),
.B(n_867),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_902),
.B(n_878),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_970),
.B(n_776),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_986),
.B(n_813),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_1000),
.A2(n_829),
.B(n_798),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_898),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_988),
.A2(n_875),
.B(n_886),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_944),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_916),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_993),
.Y(n_1044)
);

AO31x2_ASAP7_75t_L g1045 ( 
.A1(n_999),
.A2(n_875),
.A3(n_785),
.B(n_880),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_965),
.Y(n_1046)
);

CKINVDCx11_ASAP7_75t_R g1047 ( 
.A(n_955),
.Y(n_1047)
);

NOR3xp33_ASAP7_75t_SL g1048 ( 
.A(n_984),
.B(n_813),
.C(n_875),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1018),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_914),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_895),
.A2(n_764),
.B(n_907),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_978),
.B(n_1005),
.Y(n_1052)
);

AO32x2_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_764),
.A3(n_1011),
.B1(n_972),
.B2(n_919),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_904),
.B(n_913),
.Y(n_1054)
);

AO32x2_ASAP7_75t_L g1055 ( 
.A1(n_950),
.A2(n_939),
.A3(n_995),
.B1(n_917),
.B2(n_1007),
.Y(n_1055)
);

OAI21x1_ASAP7_75t_L g1056 ( 
.A1(n_1012),
.A2(n_990),
.B(n_1009),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_898),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1019),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1020),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_892),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_898),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_899),
.B(n_979),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_891),
.A2(n_911),
.B(n_908),
.C(n_906),
.Y(n_1063)
);

AOI221x1_ASAP7_75t_L g1064 ( 
.A1(n_973),
.A2(n_974),
.B1(n_994),
.B2(n_982),
.C(n_910),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_986),
.B(n_1006),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_1017),
.A2(n_901),
.B(n_905),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1021),
.B(n_964),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_1003),
.A2(n_943),
.A3(n_951),
.B(n_945),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_903),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_906),
.A2(n_908),
.B(n_1004),
.C(n_1008),
.Y(n_1070)
);

NAND4xp25_ASAP7_75t_SL g1071 ( 
.A(n_948),
.B(n_961),
.C(n_980),
.D(n_924),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_926),
.B(n_931),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_983),
.B(n_896),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1013),
.B(n_977),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_947),
.Y(n_1075)
);

OR2x2_ASAP7_75t_L g1076 ( 
.A(n_927),
.B(n_912),
.Y(n_1076)
);

AOI21x1_ASAP7_75t_L g1077 ( 
.A1(n_934),
.A2(n_943),
.B(n_953),
.Y(n_1077)
);

AOI21x1_ASAP7_75t_L g1078 ( 
.A1(n_945),
.A2(n_953),
.B(n_951),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_954),
.B(n_975),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_952),
.A2(n_933),
.B(n_937),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1001),
.A2(n_989),
.B(n_893),
.Y(n_1081)
);

NAND3x1_ASAP7_75t_L g1082 ( 
.A(n_967),
.B(n_987),
.C(n_997),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_949),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_956),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_950),
.A2(n_981),
.B(n_915),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_950),
.A2(n_915),
.B(n_941),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_1006),
.B(n_904),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_900),
.B(n_963),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_958),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_922),
.Y(n_1090)
);

AO21x2_ASAP7_75t_L g1091 ( 
.A1(n_921),
.A2(n_940),
.B(n_932),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_930),
.B(n_1022),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_930),
.B(n_960),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_960),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_957),
.A2(n_962),
.B(n_968),
.C(n_942),
.Y(n_1095)
);

AOI211x1_ASAP7_75t_L g1096 ( 
.A1(n_946),
.A2(n_923),
.B(n_991),
.C(n_996),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_938),
.B(n_935),
.Y(n_1097)
);

AOI21x1_ASAP7_75t_L g1098 ( 
.A1(n_936),
.A2(n_998),
.B(n_971),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_1014),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_1002),
.A2(n_918),
.B(n_959),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_1015),
.Y(n_1101)
);

NAND2xp33_ASAP7_75t_L g1102 ( 
.A(n_1010),
.B(n_925),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_971),
.A2(n_992),
.B(n_988),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_971),
.A2(n_985),
.B(n_771),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_902),
.B(n_581),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_913),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_992),
.A2(n_988),
.B(n_999),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_902),
.A2(n_852),
.B1(n_749),
.B2(n_848),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_992),
.A2(n_575),
.B(n_581),
.C(n_852),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_916),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_992),
.A2(n_575),
.B(n_581),
.C(n_852),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_920),
.B(n_852),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_902),
.B(n_581),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_992),
.A2(n_575),
.B(n_581),
.C(n_852),
.Y(n_1114)
);

AO32x2_ASAP7_75t_L g1115 ( 
.A1(n_1023),
.A2(n_897),
.A3(n_1011),
.B1(n_972),
.B2(n_840),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_929),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_985),
.A2(n_771),
.B(n_729),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_999),
.A2(n_910),
.B(n_982),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_916),
.Y(n_1119)
);

OR2x6_ASAP7_75t_L g1120 ( 
.A(n_954),
.B(n_732),
.Y(n_1120)
);

OAI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_902),
.A2(n_356),
.B1(n_853),
.B2(n_767),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_976),
.B(n_793),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_986),
.B(n_1006),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_920),
.B(n_852),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_974),
.A2(n_575),
.B1(n_853),
.B2(n_852),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_902),
.B(n_581),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_916),
.Y(n_1127)
);

INVxp67_ASAP7_75t_SL g1128 ( 
.A(n_929),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_902),
.A2(n_852),
.B1(n_749),
.B2(n_848),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_916),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_902),
.B(n_581),
.Y(n_1131)
);

NAND3x1_ASAP7_75t_L g1132 ( 
.A(n_974),
.B(n_984),
.C(n_724),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_916),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_916),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_902),
.B(n_581),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_902),
.B(n_581),
.Y(n_1136)
);

AO31x2_ASAP7_75t_L g1137 ( 
.A1(n_999),
.A2(n_897),
.A3(n_982),
.B(n_1003),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_929),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_976),
.B(n_793),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_985),
.A2(n_771),
.B(n_729),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_914),
.Y(n_1141)
);

CKINVDCx14_ASAP7_75t_R g1142 ( 
.A(n_969),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_914),
.B(n_853),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_916),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_914),
.B(n_853),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_999),
.A2(n_897),
.A3(n_982),
.B(n_1003),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1043),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1114),
.C(n_1136),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_1088),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1044),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1125),
.A2(n_1062),
.B1(n_1124),
.B2(n_1112),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1105),
.A2(n_1113),
.B(n_1126),
.C(n_1135),
.Y(n_1152)
);

NAND2x1p5_ASAP7_75t_L g1153 ( 
.A(n_1087),
.B(n_1100),
.Y(n_1153)
);

OR2x6_ASAP7_75t_L g1154 ( 
.A(n_1120),
.B(n_1096),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_1121),
.A2(n_1072),
.B1(n_1125),
.B2(n_1071),
.C(n_1063),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1110),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1131),
.B(n_1073),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1067),
.B(n_1029),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1039),
.A2(n_1051),
.B(n_1024),
.Y(n_1159)
);

AND2x4_ASAP7_75t_L g1160 ( 
.A(n_1120),
.B(n_1065),
.Y(n_1160)
);

AO31x2_ASAP7_75t_L g1161 ( 
.A1(n_1104),
.A2(n_1064),
.A3(n_1086),
.B(n_1085),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1081),
.A2(n_1041),
.B(n_1107),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1041),
.A2(n_1077),
.B(n_1098),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_R g1164 ( 
.A(n_1048),
.B(n_1120),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1078),
.A2(n_1034),
.B(n_1107),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1031),
.A2(n_1103),
.B(n_1093),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1095),
.A2(n_1118),
.B(n_1070),
.Y(n_1167)
);

AOI21xp33_ASAP7_75t_L g1168 ( 
.A1(n_1032),
.A2(n_1129),
.B(n_1108),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_1103),
.A2(n_1046),
.B1(n_1116),
.B2(n_1141),
.C(n_1050),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1122),
.B(n_1139),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1047),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1087),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1035),
.A2(n_1036),
.B1(n_1076),
.B2(n_1058),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1030),
.A2(n_1037),
.B(n_1115),
.C(n_1074),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1060),
.A2(n_1092),
.B(n_1094),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1119),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1033),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1127),
.A2(n_1144),
.B(n_1134),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1030),
.A2(n_1115),
.B(n_1079),
.C(n_1130),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1049),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1133),
.A2(n_1059),
.B(n_1089),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1101),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_L g1183 ( 
.A1(n_1052),
.A2(n_1145),
.B1(n_1143),
.B2(n_1083),
.Y(n_1183)
);

OA21x2_ASAP7_75t_L g1184 ( 
.A1(n_1075),
.A2(n_1146),
.B(n_1137),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1084),
.A2(n_1090),
.B(n_1082),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1065),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1132),
.A2(n_1026),
.B(n_1042),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1141),
.A2(n_1128),
.B1(n_1096),
.B2(n_1028),
.Y(n_1188)
);

INVx1_ASAP7_75t_SL g1189 ( 
.A(n_1138),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1054),
.A2(n_1045),
.B(n_1146),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_1123),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1045),
.A2(n_1137),
.B(n_1068),
.Y(n_1192)
);

NOR2xp67_ASAP7_75t_L g1193 ( 
.A(n_1106),
.B(n_1099),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1123),
.B(n_1038),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1038),
.B(n_1097),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1068),
.A2(n_1091),
.B(n_1053),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1068),
.A2(n_1091),
.B(n_1053),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1040),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1053),
.A2(n_1115),
.B(n_1027),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1027),
.A2(n_1055),
.B(n_1102),
.Y(n_1200)
);

NOR4xp25_ASAP7_75t_L g1201 ( 
.A(n_1027),
.B(n_1055),
.C(n_1142),
.D(n_1025),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1055),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1057),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_1061),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1061),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1043),
.Y(n_1206)
);

AND2x4_ASAP7_75t_L g1207 ( 
.A(n_1120),
.B(n_1065),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1120),
.B(n_1065),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1087),
.B(n_773),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1047),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1125),
.A2(n_575),
.B1(n_853),
.B2(n_974),
.Y(n_1213)
);

CKINVDCx6p67_ASAP7_75t_R g1214 ( 
.A(n_1047),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1043),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1125),
.A2(n_1113),
.B1(n_1126),
.B2(n_1105),
.Y(n_1216)
);

HB1xp67_ASAP7_75t_L g1217 ( 
.A(n_1107),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1069),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1080),
.A2(n_1066),
.B(n_1056),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1120),
.B(n_1096),
.Y(n_1220)
);

BUFx3_ASAP7_75t_L g1221 ( 
.A(n_1065),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1076),
.B(n_1058),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_L g1223 ( 
.A(n_1125),
.B(n_575),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1114),
.C(n_575),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1080),
.A2(n_1056),
.B(n_1066),
.Y(n_1225)
);

BUFx2_ASAP7_75t_SL g1226 ( 
.A(n_1101),
.Y(n_1226)
);

AND2x4_ASAP7_75t_L g1227 ( 
.A(n_1120),
.B(n_1065),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1069),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1109),
.B(n_1111),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1088),
.Y(n_1230)
);

INVx6_ASAP7_75t_L g1231 ( 
.A(n_1087),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1050),
.B(n_751),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1233)
);

AO31x2_ASAP7_75t_L g1234 ( 
.A1(n_1104),
.A2(n_1064),
.A3(n_1086),
.B(n_1085),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1125),
.A2(n_1113),
.B1(n_1126),
.B2(n_1105),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1114),
.C(n_575),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1117),
.A2(n_1140),
.B(n_1095),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1120),
.B(n_1065),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1069),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1087),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1125),
.B(n_575),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1117),
.A2(n_1140),
.B(n_1095),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1109),
.A2(n_575),
.B(n_1111),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1125),
.A2(n_575),
.B1(n_974),
.B2(n_928),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_1047),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_SL g1246 ( 
.A(n_1109),
.B(n_1111),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1217),
.B(n_1184),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1178),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1223),
.A2(n_1241),
.B(n_1224),
.C(n_1236),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1222),
.B(n_1158),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1154),
.B(n_1220),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1216),
.B(n_1235),
.Y(n_1252)
);

AOI21x1_ASAP7_75t_SL g1253 ( 
.A1(n_1209),
.A2(n_1233),
.B(n_1210),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1170),
.B(n_1149),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1230),
.B(n_1151),
.Y(n_1255)
);

AOI221x1_ASAP7_75t_SL g1256 ( 
.A1(n_1241),
.A2(n_1168),
.B1(n_1188),
.B2(n_1232),
.C(n_1157),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1152),
.B(n_1173),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1213),
.A2(n_1244),
.B1(n_1155),
.B2(n_1183),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1154),
.B(n_1220),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1237),
.A2(n_1242),
.B(n_1224),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1244),
.B(n_1189),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1217),
.B(n_1184),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1187),
.A2(n_1148),
.B1(n_1169),
.B2(n_1220),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1154),
.B(n_1160),
.Y(n_1265)
);

OA21x2_ASAP7_75t_L g1266 ( 
.A1(n_1163),
.A2(n_1165),
.B(n_1196),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1184),
.B(n_1199),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1201),
.B(n_1166),
.Y(n_1268)
);

AOI21x1_ASAP7_75t_SL g1269 ( 
.A1(n_1195),
.A2(n_1160),
.B(n_1207),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1226),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1162),
.B(n_1200),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1174),
.A2(n_1179),
.B(n_1238),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1202),
.B(n_1179),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1178),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1193),
.A2(n_1191),
.B1(n_1186),
.B2(n_1231),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1212),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1186),
.A2(n_1191),
.B1(n_1231),
.B2(n_1221),
.Y(n_1277)
);

AOI211xp5_ASAP7_75t_SL g1278 ( 
.A1(n_1172),
.A2(n_1240),
.B(n_1150),
.C(n_1215),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_SL g1279 ( 
.A1(n_1207),
.A2(n_1238),
.B(n_1208),
.Y(n_1279)
);

AND2x4_ASAP7_75t_L g1280 ( 
.A(n_1208),
.B(n_1227),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1197),
.A2(n_1185),
.B(n_1175),
.C(n_1190),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1147),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1177),
.B(n_1180),
.Y(n_1283)
);

INVx3_ASAP7_75t_SL g1284 ( 
.A(n_1182),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1192),
.A2(n_1159),
.B(n_1219),
.Y(n_1285)
);

INVx2_ASAP7_75t_SL g1286 ( 
.A(n_1156),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1212),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_SL g1288 ( 
.A1(n_1164),
.A2(n_1245),
.B(n_1214),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1177),
.B(n_1180),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1218),
.B(n_1239),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1176),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_L g1292 ( 
.A1(n_1206),
.A2(n_1182),
.B1(n_1153),
.B2(n_1211),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1228),
.B(n_1181),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1153),
.A2(n_1211),
.B1(n_1205),
.B2(n_1203),
.Y(n_1294)
);

O2A1O1Ixp5_ASAP7_75t_L g1295 ( 
.A1(n_1198),
.A2(n_1204),
.B(n_1161),
.C(n_1234),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1171),
.A2(n_1245),
.B1(n_1161),
.B2(n_1234),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1161),
.B(n_1234),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1225),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1188),
.Y(n_1299)
);

AND2x4_ASAP7_75t_L g1300 ( 
.A(n_1154),
.B(n_1220),
.Y(n_1300)
);

HB1xp67_ASAP7_75t_L g1301 ( 
.A(n_1188),
.Y(n_1301)
);

BUFx2_ASAP7_75t_SL g1302 ( 
.A(n_1232),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1154),
.B(n_1220),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1188),
.Y(n_1304)
);

O2A1O1Ixp5_ASAP7_75t_L g1305 ( 
.A1(n_1243),
.A2(n_1229),
.B(n_1246),
.C(n_1241),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1213),
.A2(n_1223),
.B1(n_1241),
.B2(n_1244),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1223),
.A2(n_1241),
.B(n_1224),
.C(n_1111),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1170),
.Y(n_1308)
);

CKINVDCx16_ASAP7_75t_R g1309 ( 
.A(n_1226),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_1188),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1216),
.B(n_1235),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1223),
.A2(n_1241),
.B(n_1167),
.C(n_1236),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1167),
.A2(n_1103),
.B(n_1163),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1217),
.B(n_1184),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1248),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1251),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1274),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1247),
.B(n_1263),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1252),
.B(n_1311),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1314),
.B(n_1271),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1267),
.B(n_1314),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1267),
.B(n_1297),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1293),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1297),
.B(n_1273),
.Y(n_1324)
);

OAI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1306),
.A2(n_1312),
.B1(n_1258),
.B2(n_1249),
.C(n_1305),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1273),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1281),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1281),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1279),
.B(n_1260),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1268),
.B(n_1313),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1295),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1268),
.B(n_1313),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1312),
.B(n_1257),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1266),
.B(n_1259),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1286),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1285),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1286),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1266),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1282),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1296),
.B(n_1298),
.Y(n_1340)
);

HB1xp67_ASAP7_75t_L g1341 ( 
.A(n_1291),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1283),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1289),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1307),
.A2(n_1269),
.B(n_1272),
.Y(n_1344)
);

INVx5_ASAP7_75t_L g1345 ( 
.A(n_1259),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1299),
.B(n_1310),
.Y(n_1346)
);

HB1xp67_ASAP7_75t_L g1347 ( 
.A(n_1301),
.Y(n_1347)
);

OR2x6_ASAP7_75t_L g1348 ( 
.A(n_1279),
.B(n_1303),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1304),
.B(n_1300),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1315),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1315),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1335),
.Y(n_1352)
);

OAI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1325),
.A2(n_1264),
.B1(n_1278),
.B2(n_1262),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1322),
.B(n_1272),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1323),
.B(n_1256),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1335),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1315),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1317),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1325),
.B(n_1255),
.Y(n_1360)
);

INVx4_ASAP7_75t_L g1361 ( 
.A(n_1348),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1317),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1317),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1321),
.B(n_1265),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1345),
.B(n_1280),
.Y(n_1365)
);

INVx4_ASAP7_75t_R g1366 ( 
.A(n_1316),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1345),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1321),
.B(n_1290),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1323),
.B(n_1250),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1337),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_1319),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1324),
.B(n_1261),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1320),
.B(n_1254),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1323),
.B(n_1308),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1320),
.B(n_1292),
.Y(n_1375)
);

OAI33xp33_ASAP7_75t_L g1376 ( 
.A1(n_1319),
.A2(n_1294),
.A3(n_1275),
.B1(n_1287),
.B2(n_1277),
.B3(n_1253),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1324),
.B(n_1330),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1326),
.B(n_1270),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1353),
.A2(n_1333),
.B1(n_1329),
.B2(n_1344),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1350),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1353),
.A2(n_1333),
.B(n_1332),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1350),
.Y(n_1382)
);

AOI221xp5_ASAP7_75t_L g1383 ( 
.A1(n_1360),
.A2(n_1332),
.B1(n_1330),
.B2(n_1347),
.C(n_1328),
.Y(n_1383)
);

NAND4xp25_ASAP7_75t_SL g1384 ( 
.A(n_1354),
.B(n_1276),
.C(n_1330),
.D(n_1332),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1365),
.B(n_1367),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1377),
.B(n_1324),
.Y(n_1386)
);

INVx2_ASAP7_75t_SL g1387 ( 
.A(n_1366),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1377),
.B(n_1358),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1360),
.A2(n_1329),
.B1(n_1346),
.B2(n_1348),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1355),
.B(n_1347),
.C(n_1328),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1351),
.A2(n_1331),
.B(n_1336),
.Y(n_1391)
);

OAI221xp5_ASAP7_75t_L g1392 ( 
.A1(n_1355),
.A2(n_1329),
.B1(n_1302),
.B2(n_1346),
.C(n_1284),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1369),
.B(n_1346),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1352),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1378),
.B(n_1328),
.C(n_1327),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1371),
.B(n_1309),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1357),
.Y(n_1397)
);

OR2x2_ASAP7_75t_L g1398 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1398)
);

OR2x2_ASAP7_75t_L g1399 ( 
.A(n_1373),
.B(n_1318),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1357),
.A2(n_1331),
.B(n_1336),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1359),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1375),
.A2(n_1329),
.B1(n_1327),
.B2(n_1340),
.C(n_1349),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1377),
.B(n_1334),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1359),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1375),
.B(n_1318),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1352),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1367),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1376),
.A2(n_1329),
.B1(n_1344),
.B2(n_1348),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1376),
.A2(n_1329),
.B1(n_1344),
.B2(n_1354),
.Y(n_1409)
);

AOI221xp5_ASAP7_75t_L g1410 ( 
.A1(n_1374),
.A2(n_1327),
.B1(n_1331),
.B2(n_1342),
.C(n_1343),
.Y(n_1410)
);

INVxp67_ASAP7_75t_L g1411 ( 
.A(n_1369),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1362),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1374),
.A2(n_1343),
.B1(n_1342),
.B2(n_1341),
.C(n_1339),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1362),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1363),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1411),
.B(n_1368),
.Y(n_1416)
);

INVx3_ASAP7_75t_L g1417 ( 
.A(n_1385),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1394),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1380),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1410),
.B(n_1368),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1380),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1405),
.B(n_1356),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_SL g1423 ( 
.A(n_1390),
.B(n_1345),
.Y(n_1423)
);

NOR2xp33_ASAP7_75t_SL g1424 ( 
.A(n_1381),
.B(n_1371),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1382),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1383),
.A2(n_1336),
.B(n_1338),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1391),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1382),
.Y(n_1428)
);

INVx4_ASAP7_75t_SL g1429 ( 
.A(n_1387),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1403),
.B(n_1354),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1406),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1397),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1385),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1397),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1401),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1385),
.Y(n_1436)
);

INVx3_ASAP7_75t_L g1437 ( 
.A(n_1407),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_R g1438 ( 
.A(n_1396),
.B(n_1276),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1407),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1400),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1413),
.B(n_1370),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1392),
.B(n_1378),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1400),
.Y(n_1443)
);

BUFx8_ASAP7_75t_L g1444 ( 
.A(n_1387),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1405),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1419),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_L g1447 ( 
.A(n_1423),
.B(n_1395),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1419),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1421),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1442),
.B(n_1420),
.Y(n_1450)
);

AOI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1424),
.A2(n_1384),
.B(n_1389),
.C(n_1402),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1421),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1430),
.B(n_1386),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1429),
.B(n_1361),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1425),
.Y(n_1455)
);

INVx2_ASAP7_75t_SL g1456 ( 
.A(n_1444),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1427),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1425),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1442),
.B(n_1372),
.Y(n_1459)
);

INVx1_ASAP7_75t_SL g1460 ( 
.A(n_1438),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1430),
.B(n_1386),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1445),
.B(n_1398),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1430),
.B(n_1388),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1428),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1428),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1432),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

OAI33xp33_ASAP7_75t_L g1468 ( 
.A1(n_1441),
.A2(n_1370),
.A3(n_1414),
.B1(n_1412),
.B2(n_1415),
.B3(n_1404),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1445),
.B(n_1422),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1420),
.B(n_1372),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1424),
.B(n_1379),
.Y(n_1473)
);

INVx2_ASAP7_75t_SL g1474 ( 
.A(n_1444),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1429),
.B(n_1403),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1429),
.B(n_1398),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1422),
.B(n_1399),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1434),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1429),
.B(n_1399),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1418),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1429),
.B(n_1358),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1433),
.B(n_1358),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1433),
.B(n_1364),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1435),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1422),
.B(n_1393),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1447),
.B(n_1423),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1469),
.B(n_1481),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1475),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1446),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1457),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1475),
.B(n_1476),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1446),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1483),
.B(n_1436),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1450),
.B(n_1441),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1448),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1457),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1477),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1483),
.B(n_1436),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1448),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1449),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1472),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1469),
.B(n_1431),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

NOR2x1_ASAP7_75t_L g1506 ( 
.A(n_1460),
.B(n_1439),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1462),
.B(n_1478),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1476),
.B(n_1433),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1463),
.B(n_1417),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.B(n_1417),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1484),
.B(n_1417),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1452),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1459),
.B(n_1431),
.Y(n_1513)
);

AO22x1_ASAP7_75t_L g1514 ( 
.A1(n_1456),
.A2(n_1287),
.B1(n_1284),
.B2(n_1444),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1452),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1471),
.B(n_1416),
.Y(n_1516)
);

NOR2x1_ASAP7_75t_L g1517 ( 
.A(n_1473),
.B(n_1439),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1484),
.B(n_1417),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1462),
.B(n_1418),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1456),
.B(n_1417),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1485),
.B(n_1453),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1485),
.B(n_1437),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1506),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1489),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1496),
.B(n_1453),
.Y(n_1525)
);

INVx1_ASAP7_75t_SL g1526 ( 
.A(n_1504),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1517),
.A2(n_1468),
.B1(n_1361),
.B2(n_1409),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1489),
.B(n_1461),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1504),
.B(n_1461),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1513),
.B(n_1519),
.Y(n_1530)
);

AND3x1_ASAP7_75t_L g1531 ( 
.A(n_1490),
.B(n_1451),
.C(n_1474),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1514),
.B(n_1474),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1493),
.B(n_1477),
.Y(n_1533)
);

INVx4_ASAP7_75t_L g1534 ( 
.A(n_1520),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1493),
.B(n_1480),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1480),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_SL g1537 ( 
.A1(n_1488),
.A2(n_1438),
.B1(n_1426),
.B2(n_1454),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1488),
.A2(n_1408),
.B1(n_1478),
.B2(n_1487),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1491),
.Y(n_1539)
);

OAI21xp33_ASAP7_75t_L g1540 ( 
.A1(n_1488),
.A2(n_1487),
.B(n_1464),
.Y(n_1540)
);

INVx1_ASAP7_75t_SL g1541 ( 
.A(n_1519),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1507),
.B(n_1455),
.Y(n_1542)
);

CKINVDCx16_ASAP7_75t_R g1543 ( 
.A(n_1488),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1514),
.B(n_1454),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1508),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1521),
.B(n_1416),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1490),
.Y(n_1547)
);

INVx1_ASAP7_75t_SL g1548 ( 
.A(n_1523),
.Y(n_1548)
);

AOI32xp33_ASAP7_75t_L g1549 ( 
.A1(n_1531),
.A2(n_1508),
.A3(n_1500),
.B1(n_1495),
.B2(n_1499),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1543),
.A2(n_1527),
.B1(n_1537),
.B2(n_1544),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1541),
.B(n_1526),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1534),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1553)
);

AOI21xp5_ASAP7_75t_L g1554 ( 
.A1(n_1540),
.A2(n_1499),
.B(n_1520),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1534),
.Y(n_1555)
);

AOI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1532),
.A2(n_1533),
.B1(n_1535),
.B2(n_1536),
.Y(n_1556)
);

AOI21xp5_ASAP7_75t_L g1557 ( 
.A1(n_1538),
.A2(n_1520),
.B(n_1516),
.Y(n_1557)
);

OAI31xp33_ASAP7_75t_L g1558 ( 
.A1(n_1524),
.A2(n_1497),
.A3(n_1491),
.B(n_1515),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1547),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1495),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_SL g1561 ( 
.A(n_1534),
.B(n_1500),
.Y(n_1561)
);

OR2x2_ASAP7_75t_L g1562 ( 
.A(n_1528),
.B(n_1494),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1547),
.Y(n_1563)
);

OAI32xp33_ASAP7_75t_L g1564 ( 
.A1(n_1545),
.A2(n_1518),
.A3(n_1511),
.B1(n_1522),
.B2(n_1512),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1539),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1539),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_SL g1567 ( 
.A(n_1548),
.B(n_1544),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1548),
.B(n_1545),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1559),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1563),
.B(n_1533),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1551),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1560),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1561),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1552),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1565),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1555),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1556),
.B(n_1535),
.Y(n_1577)
);

AOI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1573),
.A2(n_1553),
.B(n_1549),
.Y(n_1578)
);

NOR2xp67_ASAP7_75t_L g1579 ( 
.A(n_1573),
.B(n_1554),
.Y(n_1579)
);

AOI221x1_ASAP7_75t_L g1580 ( 
.A1(n_1569),
.A2(n_1566),
.B1(n_1550),
.B2(n_1557),
.C(n_1536),
.Y(n_1580)
);

AOI21xp33_ASAP7_75t_L g1581 ( 
.A1(n_1567),
.A2(n_1564),
.B(n_1558),
.Y(n_1581)
);

OAI21xp33_ASAP7_75t_L g1582 ( 
.A1(n_1577),
.A2(n_1529),
.B(n_1525),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1577),
.B(n_1544),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1568),
.Y(n_1584)
);

AOI222xp33_ASAP7_75t_L g1585 ( 
.A1(n_1571),
.A2(n_1558),
.B1(n_1494),
.B2(n_1505),
.C1(n_1501),
.C2(n_1502),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1572),
.A2(n_1544),
.B(n_1562),
.Y(n_1586)
);

OAI32xp33_ASAP7_75t_L g1587 ( 
.A1(n_1572),
.A2(n_1542),
.A3(n_1502),
.B1(n_1501),
.B2(n_1505),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1570),
.Y(n_1588)
);

AOI21xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1581),
.A2(n_1574),
.B(n_1575),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1584),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1583),
.Y(n_1591)
);

OAI221xp5_ASAP7_75t_L g1592 ( 
.A1(n_1578),
.A2(n_1579),
.B1(n_1582),
.B2(n_1586),
.C(n_1576),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1587),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1591),
.B(n_1588),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1591),
.B(n_1585),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1593),
.B(n_1580),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1589),
.B(n_1585),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1590),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1594),
.Y(n_1600)
);

AO22x2_ASAP7_75t_L g1601 ( 
.A1(n_1597),
.A2(n_1512),
.B1(n_1515),
.B2(n_1498),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1595),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1596),
.B(n_1546),
.Y(n_1603)
);

INVx3_ASAP7_75t_SL g1604 ( 
.A(n_1598),
.Y(n_1604)
);

NOR3xp33_ASAP7_75t_L g1605 ( 
.A(n_1602),
.B(n_1599),
.C(n_1498),
.Y(n_1605)
);

AOI322xp5_ASAP7_75t_L g1606 ( 
.A1(n_1603),
.A2(n_1518),
.A3(n_1511),
.B1(n_1492),
.B2(n_1503),
.C1(n_1509),
.C2(n_1510),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1600),
.A2(n_1503),
.B1(n_1492),
.B2(n_1509),
.Y(n_1607)
);

OR3x1_ASAP7_75t_L g1608 ( 
.A(n_1605),
.B(n_1604),
.C(n_1601),
.Y(n_1608)
);

NOR3xp33_ASAP7_75t_L g1609 ( 
.A(n_1608),
.B(n_1601),
.C(n_1607),
.Y(n_1609)
);

OR4x1_ASAP7_75t_L g1610 ( 
.A(n_1609),
.B(n_1606),
.C(n_1455),
.D(n_1458),
.Y(n_1610)
);

AOI22x1_ASAP7_75t_L g1611 ( 
.A1(n_1610),
.A2(n_1472),
.B1(n_1510),
.B2(n_1522),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1611),
.A2(n_1454),
.B1(n_1482),
.B2(n_1479),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1612),
.A2(n_1486),
.B1(n_1482),
.B2(n_1479),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1613),
.A2(n_1454),
.B1(n_1470),
.B2(n_1467),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1614),
.B(n_1458),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1614),
.A2(n_1486),
.B(n_1470),
.Y(n_1616)
);

AOI22x1_ASAP7_75t_L g1617 ( 
.A1(n_1616),
.A2(n_1288),
.B1(n_1467),
.B2(n_1466),
.Y(n_1617)
);

OAI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1617),
.A2(n_1615),
.B1(n_1466),
.B2(n_1465),
.Y(n_1618)
);

AOI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1618),
.A2(n_1465),
.B(n_1443),
.C(n_1440),
.Y(n_1619)
);


endmodule