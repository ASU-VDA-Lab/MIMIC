module fake_jpeg_9679_n_73 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_55;
wire n_27;
wire n_64;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_24;
wire n_36;
wire n_62;
wire n_56;
wire n_31;
wire n_25;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_3),
.B(n_19),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_7),
.A2(n_5),
.B(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_0),
.B(n_11),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_0),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_1),
.C(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_44),
.B(n_49),
.Y(n_54)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_47),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_30),
.Y(n_51)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_39),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_59),
.B(n_43),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_34),
.Y(n_62)
);

A2O1A1O1Ixp25_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_57),
.B(n_54),
.C(n_51),
.D(n_26),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_51),
.A3(n_23),
.B1(n_37),
.B2(n_49),
.C(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_23),
.C(n_22),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_31),
.B1(n_33),
.B2(n_25),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_48),
.B1(n_32),
.B2(n_43),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_SL g69 ( 
.A1(n_67),
.A2(n_28),
.B(n_40),
.C(n_46),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_30),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_70),
.B(n_24),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_50),
.Y(n_73)
);


endmodule