module fake_jpeg_8873_n_234 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_234);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_234;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_23),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_55),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_29),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_60),
.B(n_62),
.C(n_63),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_49),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_22),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_26),
.B1(n_23),
.B2(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_63),
.B1(n_42),
.B2(n_18),
.Y(n_66)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_41),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_32),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_16),
.B1(n_31),
.B2(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_22),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_18),
.Y(n_65)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_78),
.B(n_47),
.C(n_65),
.Y(n_99)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_67),
.A2(n_73),
.B1(n_82),
.B2(n_68),
.Y(n_94)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_75),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_69),
.B(n_77),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_62),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_38),
.B1(n_41),
.B2(n_57),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_17),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_41),
.B1(n_44),
.B2(n_17),
.Y(n_78)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_60),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_87),
.Y(n_105)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_95),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_48),
.C(n_53),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_104),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_53),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_56),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_99),
.A2(n_58),
.B1(n_46),
.B2(n_61),
.Y(n_113)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_100),
.Y(n_133)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_44),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_55),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_58),
.B1(n_61),
.B2(n_50),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_97),
.B1(n_110),
.B2(n_103),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_0),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_108),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_59),
.B(n_25),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_80),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_40),
.B1(n_43),
.B2(n_16),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_123),
.A2(n_126),
.B1(n_130),
.B2(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_20),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_105),
.A2(n_40),
.B1(n_31),
.B2(n_33),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_92),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_92),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_33),
.B1(n_28),
.B2(n_20),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_34),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_90),
.C(n_93),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_110),
.B1(n_88),
.B2(n_100),
.Y(n_140)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_132),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_135),
.B(n_136),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_116),
.A2(n_102),
.B1(n_101),
.B2(n_97),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_140),
.B1(n_117),
.B2(n_125),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_141),
.B(n_145),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_150),
.B(n_154),
.C(n_138),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_34),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_111),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_117),
.B(n_13),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_150),
.A2(n_152),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_91),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_106),
.B(n_108),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_114),
.B(n_130),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_165),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_151),
.A2(n_116),
.B(n_121),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_174),
.B(n_32),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_131),
.Y(n_162)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_162),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_112),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_143),
.C(n_171),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_173),
.B1(n_134),
.B2(n_30),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_34),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_170),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_155),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_176),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_184),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_160),
.B(n_159),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_139),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_180),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_153),
.C(n_144),
.Y(n_180)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_167),
.C(n_170),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_168),
.B1(n_172),
.B2(n_156),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_30),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_187),
.B(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_19),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_190),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_172),
.B(n_15),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_183),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_201),
.B(n_182),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_157),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_197),
.B(n_202),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_200),
.B(n_176),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_156),
.B(n_174),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_157),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_201),
.B(n_175),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_173),
.B1(n_177),
.B2(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_195),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_206),
.B(n_195),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_158),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_158),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_203),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_194),
.B(n_198),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_167),
.C(n_19),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_210),
.B(n_15),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_215),
.C(n_210),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_9),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_211),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_9),
.Y(n_220)
);

NAND3xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_199),
.C(n_10),
.Y(n_218)
);

AOI31xp67_ASAP7_75t_SL g223 ( 
.A1(n_218),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_216),
.C(n_212),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_222),
.A2(n_223),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_224),
.B(n_3),
.C(n_4),
.Y(n_228)
);

AOI311xp33_ASAP7_75t_L g229 ( 
.A1(n_227),
.A2(n_3),
.A3(n_4),
.B(n_5),
.C(n_6),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_3),
.Y(n_230)
);

AOI322xp5_ASAP7_75t_L g231 ( 
.A1(n_229),
.A2(n_4),
.A3(n_5),
.B1(n_224),
.B2(n_225),
.C1(n_226),
.C2(n_223),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

BUFx24_ASAP7_75t_SL g233 ( 
.A(n_232),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_233),
.B(n_231),
.Y(n_234)
);


endmodule