module real_aes_6688_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_741;
wire n_283;
wire n_252;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g480 ( .A1(n_0), .A2(n_184), .B(n_481), .C(n_484), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_1), .B(n_475), .Y(n_486) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVx1_ASAP7_75t_L g233 ( .A(n_3), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_4), .B(n_172), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_5), .A2(n_459), .B(n_529), .Y(n_528) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_6), .A2(n_9), .B1(n_442), .B2(n_758), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_6), .Y(n_758) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_7), .A2(n_189), .B(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_40), .B1(n_145), .B2(n_157), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_9), .A2(n_129), .B1(n_130), .B2(n_442), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_9), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_10), .B(n_189), .Y(n_222) );
AND2x6_ASAP7_75t_L g160 ( .A(n_11), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_12), .A2(n_160), .B(n_462), .C(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_13), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_14), .B(n_41), .Y(n_115) );
INVx1_ASAP7_75t_L g141 ( .A(n_15), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_16), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g227 ( .A(n_17), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g102 ( .A1(n_18), .A2(n_103), .B1(n_116), .B2(n_763), .Y(n_102) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_19), .B(n_172), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_20), .B(n_187), .Y(n_205) );
AO32x2_ASAP7_75t_L g181 ( .A1(n_21), .A2(n_182), .A3(n_186), .B1(n_188), .B2(n_189), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_22), .A2(n_100), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_22), .Y(n_124) );
AND2x2_ASAP7_75t_L g523 ( .A(n_23), .B(n_137), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_24), .B(n_145), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_25), .B(n_187), .Y(n_235) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_26), .A2(n_56), .B1(n_145), .B2(n_157), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g198 ( .A1(n_27), .A2(n_82), .B1(n_145), .B2(n_149), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_28), .B(n_145), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_29), .A2(n_188), .B(n_462), .C(n_464), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_30), .A2(n_188), .B(n_462), .C(n_541), .Y(n_540) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_31), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_32), .B(n_137), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_33), .A2(n_459), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_34), .B(n_137), .Y(n_179) );
INVx2_ASAP7_75t_L g147 ( .A(n_35), .Y(n_147) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_36), .A2(n_493), .B(n_494), .C(n_498), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_37), .B(n_145), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_38), .B(n_137), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_39), .B(n_152), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_42), .B(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_43), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_44), .B(n_172), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_45), .B(n_459), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_46), .A2(n_493), .B(n_498), .C(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_47), .B(n_145), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g118 ( .A(n_48), .B(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g482 ( .A(n_49), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_50), .A2(n_91), .B1(n_157), .B2(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g521 ( .A(n_51), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_52), .B(n_145), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_53), .B(n_145), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_54), .B(n_459), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_55), .B(n_220), .Y(n_219) );
AOI22xp33_ASAP7_75t_SL g209 ( .A1(n_57), .A2(n_61), .B1(n_145), .B2(n_149), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_58), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_59), .B(n_145), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_60), .B(n_145), .Y(n_246) );
INVx1_ASAP7_75t_L g161 ( .A(n_62), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_63), .B(n_459), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_64), .B(n_475), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_65), .A2(n_220), .B(n_230), .C(n_532), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_66), .B(n_145), .Y(n_234) );
INVx1_ASAP7_75t_L g140 ( .A(n_67), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_68), .Y(n_752) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_69), .B(n_172), .Y(n_496) );
AO32x2_ASAP7_75t_L g194 ( .A1(n_70), .A2(n_188), .A3(n_189), .B1(n_195), .B2(n_199), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_71), .B(n_173), .Y(n_552) );
INVx1_ASAP7_75t_L g245 ( .A(n_72), .Y(n_245) );
INVx1_ASAP7_75t_L g170 ( .A(n_73), .Y(n_170) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_74), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_75), .B(n_466), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_76), .A2(n_462), .B(n_498), .C(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g754 ( .A(n_77), .B(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_77), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_78), .B(n_149), .Y(n_171) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_79), .Y(n_530) );
INVx1_ASAP7_75t_L g109 ( .A(n_80), .Y(n_109) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_81), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_83), .B(n_157), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_84), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_85), .B(n_149), .Y(n_176) );
INVx2_ASAP7_75t_L g138 ( .A(n_86), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_87), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_88), .B(n_159), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_89), .B(n_149), .Y(n_216) );
OR2x2_ASAP7_75t_L g111 ( .A(n_90), .B(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g445 ( .A(n_90), .B(n_113), .Y(n_445) );
INVx2_ASAP7_75t_L g740 ( .A(n_90), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_92), .A2(n_101), .B1(n_149), .B2(n_150), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_93), .B(n_459), .Y(n_491) );
INVx1_ASAP7_75t_L g495 ( .A(n_94), .Y(n_495) );
INVxp67_ASAP7_75t_L g533 ( .A(n_95), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_96), .B(n_149), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_97), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g508 ( .A(n_98), .Y(n_508) );
INVx1_ASAP7_75t_L g548 ( .A(n_99), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_100), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx6p67_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_L g764 ( .A(n_106), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_110), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_SL g119 ( .A(n_111), .Y(n_119) );
INVx1_ASAP7_75t_SL g762 ( .A(n_111), .Y(n_762) );
NOR2x2_ASAP7_75t_L g748 ( .A(n_112), .B(n_740), .Y(n_748) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g739 ( .A(n_113), .B(n_740), .Y(n_739) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_120), .Y(n_117) );
OAI32xp33_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_745), .A3(n_749), .B1(n_750), .B2(n_753), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_125), .B1(n_741), .B2(n_742), .Y(n_121) );
INVx1_ASAP7_75t_L g741 ( .A(n_122), .Y(n_741) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22x1_ASAP7_75t_SL g126 ( .A1(n_127), .A2(n_443), .B1(n_446), .B2(n_737), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_128), .A2(n_447), .B1(n_737), .B2(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_SL g755 ( .A1(n_129), .A2(n_130), .B1(n_756), .B2(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_364), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_283), .C(n_298), .D(n_324), .E(n_346), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_263), .Y(n_132) );
OAI221xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_200), .B1(n_236), .B2(n_252), .C(n_253), .Y(n_133) );
NOR2xp33_ASAP7_75t_SL g134 ( .A(n_135), .B(n_190), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_135), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g440 ( .A(n_135), .Y(n_440) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_163), .Y(n_135) );
INVx1_ASAP7_75t_L g280 ( .A(n_136), .Y(n_280) );
AND2x2_ASAP7_75t_L g282 ( .A(n_136), .B(n_181), .Y(n_282) );
AND2x2_ASAP7_75t_L g292 ( .A(n_136), .B(n_180), .Y(n_292) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_136), .Y(n_310) );
INVx1_ASAP7_75t_L g320 ( .A(n_136), .Y(n_320) );
OR2x2_ASAP7_75t_L g358 ( .A(n_136), .B(n_257), .Y(n_358) );
INVx2_ASAP7_75t_L g408 ( .A(n_136), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_136), .B(n_256), .Y(n_425) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_142), .B(n_162), .Y(n_136) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_137), .A2(n_167), .B(n_179), .Y(n_166) );
INVx2_ASAP7_75t_L g199 ( .A(n_137), .Y(n_199) );
INVx1_ASAP7_75t_L g472 ( .A(n_137), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_137), .A2(n_491), .B(n_492), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_137), .A2(n_518), .B(n_519), .Y(n_517) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_L g187 ( .A(n_138), .B(n_139), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_154), .B(n_160), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_148), .B(n_151), .Y(n_143) );
INVx3_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_145), .Y(n_510) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
BUFx3_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
AND2x6_ASAP7_75t_L g462 ( .A(n_146), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx1_ASAP7_75t_L g221 ( .A(n_147), .Y(n_221) );
INVx2_ASAP7_75t_L g228 ( .A(n_149), .Y(n_228) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
INVx3_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_153), .Y(n_178) );
AND2x2_ASAP7_75t_L g460 ( .A(n_153), .B(n_221), .Y(n_460) );
INVx1_ASAP7_75t_L g463 ( .A(n_153), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_158), .Y(n_154) );
O2A1O1Ixp5_ASAP7_75t_L g244 ( .A1(n_158), .A2(n_232), .B(n_245), .C(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g182 ( .A1(n_159), .A2(n_183), .B1(n_184), .B2(n_185), .Y(n_182) );
OAI22xp5_ASAP7_75t_SL g195 ( .A1(n_159), .A2(n_173), .B1(n_196), .B2(n_198), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_159), .A2(n_184), .B1(n_208), .B2(n_209), .Y(n_207) );
INVx4_ASAP7_75t_L g483 ( .A(n_159), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g167 ( .A1(n_160), .A2(n_168), .B(n_174), .Y(n_167) );
BUFx3_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_214), .B(n_217), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_160), .A2(n_226), .B(n_231), .Y(n_225) );
AND2x4_ASAP7_75t_L g459 ( .A(n_160), .B(n_460), .Y(n_459) );
INVx4_ASAP7_75t_SL g485 ( .A(n_160), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_160), .B(n_460), .Y(n_549) );
NOR2xp67_ASAP7_75t_L g163 ( .A(n_164), .B(n_180), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_165), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_165), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_SL g340 ( .A(n_165), .B(n_280), .Y(n_340) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
INVx2_ASAP7_75t_L g257 ( .A(n_166), .Y(n_257) );
OR2x2_ASAP7_75t_L g319 ( .A(n_166), .B(n_320), .Y(n_319) );
O2A1O1Ixp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_172), .Y(n_168) );
INVx2_ASAP7_75t_L g184 ( .A(n_172), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_172), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_172), .A2(n_242), .B(n_243), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_172), .B(n_533), .Y(n_532) );
INVx5_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .B(n_177), .Y(n_174) );
INVx1_ASAP7_75t_L g230 ( .A(n_177), .Y(n_230) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g466 ( .A(n_178), .Y(n_466) );
AND2x2_ASAP7_75t_L g258 ( .A(n_180), .B(n_194), .Y(n_258) );
AND2x2_ASAP7_75t_L g275 ( .A(n_180), .B(n_255), .Y(n_275) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AND2x2_ASAP7_75t_L g193 ( .A(n_181), .B(n_194), .Y(n_193) );
BUFx2_ASAP7_75t_L g278 ( .A(n_181), .Y(n_278) );
AND2x2_ASAP7_75t_L g407 ( .A(n_181), .B(n_408), .Y(n_407) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_184), .A2(n_218), .B(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g231 ( .A1(n_184), .A2(n_232), .B(n_233), .C(n_234), .Y(n_231) );
INVx2_ASAP7_75t_L g224 ( .A(n_186), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_186), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_187), .Y(n_189) );
NAND3xp33_ASAP7_75t_L g206 ( .A(n_188), .B(n_207), .C(n_210), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g240 ( .A1(n_188), .A2(n_241), .B(n_244), .Y(n_240) );
INVx4_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_213), .B(n_222), .Y(n_212) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_189), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_189), .A2(n_539), .B(n_540), .Y(n_538) );
INVx1_ASAP7_75t_L g252 ( .A(n_190), .Y(n_252) );
AND2x2_ASAP7_75t_L g190 ( .A(n_191), .B(n_193), .Y(n_190) );
AND2x2_ASAP7_75t_L g370 ( .A(n_191), .B(n_258), .Y(n_370) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g371 ( .A(n_192), .B(n_282), .Y(n_371) );
O2A1O1Ixp33_ASAP7_75t_L g338 ( .A1(n_193), .A2(n_339), .B(n_341), .C(n_343), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_193), .B(n_339), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_193), .A2(n_269), .B1(n_412), .B2(n_413), .C(n_415), .Y(n_411) );
INVx1_ASAP7_75t_L g255 ( .A(n_194), .Y(n_255) );
INVx1_ASAP7_75t_L g291 ( .A(n_194), .Y(n_291) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_194), .Y(n_300) );
INVx2_ASAP7_75t_L g484 ( .A(n_197), .Y(n_484) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_197), .Y(n_497) );
INVx1_ASAP7_75t_L g469 ( .A(n_199), .Y(n_469) );
INVx1_ASAP7_75t_SL g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
AND2x2_ASAP7_75t_L g317 ( .A(n_202), .B(n_262), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_202), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_203), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g409 ( .A(n_203), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g441 ( .A(n_203), .Y(n_441) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g271 ( .A(n_204), .Y(n_271) );
AND2x2_ASAP7_75t_L g297 ( .A(n_204), .B(n_251), .Y(n_297) );
NOR2x1_ASAP7_75t_L g306 ( .A(n_204), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g313 ( .A(n_204), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
INVx1_ASAP7_75t_L g249 ( .A(n_205), .Y(n_249) );
AO21x1_ASAP7_75t_L g248 ( .A1(n_207), .A2(n_210), .B(n_249), .Y(n_248) );
INVx3_ASAP7_75t_L g475 ( .A(n_210), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_210), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_210), .A2(n_505), .B(n_512), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_210), .B(n_513), .Y(n_512) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_210), .A2(n_547), .B(n_554), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_211), .B(n_353), .Y(n_388) );
INVx1_ASAP7_75t_SL g392 ( .A(n_211), .Y(n_392) );
AND2x2_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
INVx3_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
AND2x2_ASAP7_75t_L g262 ( .A(n_212), .B(n_239), .Y(n_262) );
AND2x2_ASAP7_75t_L g284 ( .A(n_212), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g329 ( .A(n_212), .B(n_323), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_212), .B(n_261), .Y(n_410) );
INVx2_ASAP7_75t_L g232 ( .A(n_220), .Y(n_232) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g250 ( .A(n_223), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g261 ( .A(n_223), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_223), .B(n_239), .Y(n_286) );
AND2x2_ASAP7_75t_L g322 ( .A(n_223), .B(n_323), .Y(n_322) );
OA21x2_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_235), .Y(n_223) );
OA21x2_ASAP7_75t_L g239 ( .A1(n_224), .A2(n_240), .B(n_247), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .C(n_230), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_228), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_228), .A2(n_552), .B(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_230), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_232), .A2(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_250), .Y(n_237) );
INVx1_ASAP7_75t_L g302 ( .A(n_238), .Y(n_302) );
AND2x2_ASAP7_75t_L g344 ( .A(n_238), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_238), .B(n_265), .Y(n_350) );
AOI21xp5_ASAP7_75t_SL g424 ( .A1(n_238), .A2(n_256), .B(n_279), .Y(n_424) );
AND2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_248), .Y(n_238) );
OR2x2_ASAP7_75t_L g267 ( .A(n_239), .B(n_248), .Y(n_267) );
AND2x2_ASAP7_75t_L g314 ( .A(n_239), .B(n_251), .Y(n_314) );
INVx2_ASAP7_75t_L g323 ( .A(n_239), .Y(n_323) );
INVx1_ASAP7_75t_L g429 ( .A(n_239), .Y(n_429) );
AND2x2_ASAP7_75t_L g353 ( .A(n_248), .B(n_323), .Y(n_353) );
INVx1_ASAP7_75t_L g378 ( .A(n_248), .Y(n_378) );
AND2x2_ASAP7_75t_L g287 ( .A(n_250), .B(n_271), .Y(n_287) );
AND2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_SL g417 ( .A(n_250), .Y(n_417) );
INVx2_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
AND2x2_ASAP7_75t_L g345 ( .A(n_251), .B(n_261), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_251), .B(n_429), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_258), .B(n_259), .Y(n_253) );
AND2x2_ASAP7_75t_L g360 ( .A(n_254), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g414 ( .A(n_254), .Y(n_414) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
BUFx2_ASAP7_75t_L g433 ( .A(n_255), .Y(n_433) );
BUFx2_ASAP7_75t_L g304 ( .A(n_256), .Y(n_304) );
AND2x2_ASAP7_75t_L g406 ( .A(n_256), .B(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g389 ( .A(n_257), .Y(n_389) );
AND2x4_ASAP7_75t_L g316 ( .A(n_258), .B(n_279), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_258), .B(n_340), .Y(n_352) );
AOI32xp33_ASAP7_75t_L g276 ( .A1(n_259), .A2(n_277), .A3(n_279), .B1(n_281), .B2(n_282), .Y(n_276) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx3_ASAP7_75t_L g265 ( .A(n_260), .Y(n_265) );
OR2x2_ASAP7_75t_L g401 ( .A(n_260), .B(n_357), .Y(n_401) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g270 ( .A(n_261), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g377 ( .A(n_261), .B(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g269 ( .A(n_262), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g281 ( .A(n_262), .B(n_271), .Y(n_281) );
INVx1_ASAP7_75t_L g402 ( .A(n_262), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_262), .B(n_377), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_268), .B(n_272), .C(n_276), .Y(n_263) );
OAI322xp33_ASAP7_75t_L g372 ( .A1(n_264), .A2(n_309), .A3(n_373), .B1(n_375), .B2(n_379), .C1(n_380), .C2(n_384), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVxp67_ASAP7_75t_L g337 ( .A(n_265), .Y(n_337) );
INVx1_ASAP7_75t_SL g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g391 ( .A(n_267), .B(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_267), .B(n_307), .Y(n_438) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g330 ( .A(n_270), .Y(n_330) );
OR2x2_ASAP7_75t_L g416 ( .A(n_271), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_274), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g325 ( .A(n_275), .B(n_304), .Y(n_325) );
AND2x2_ASAP7_75t_L g396 ( .A(n_275), .B(n_309), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_275), .B(n_383), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g283 ( .A1(n_277), .A2(n_284), .B1(n_287), .B2(n_288), .C(n_293), .Y(n_283) );
OR2x2_ASAP7_75t_L g294 ( .A(n_277), .B(n_290), .Y(n_294) );
AND2x2_ASAP7_75t_L g382 ( .A(n_277), .B(n_383), .Y(n_382) );
AOI32xp33_ASAP7_75t_L g421 ( .A1(n_277), .A2(n_307), .A3(n_422), .B1(n_423), .B2(n_426), .Y(n_421) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_278), .B(n_314), .C(n_337), .Y(n_355) );
AND2x2_ASAP7_75t_L g381 ( .A(n_278), .B(n_374), .Y(n_381) );
INVxp67_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
BUFx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_282), .B(n_334), .Y(n_390) );
INVx2_ASAP7_75t_L g400 ( .A(n_282), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_282), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g369 ( .A(n_285), .Y(n_369) );
OR2x2_ASAP7_75t_L g295 ( .A(n_286), .B(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_288), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_291), .Y(n_374) );
AND2x2_ASAP7_75t_L g333 ( .A(n_292), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g379 ( .A(n_292), .Y(n_379) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_292), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI21xp33_ASAP7_75t_SL g318 ( .A1(n_294), .A2(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g412 ( .A(n_297), .B(n_322), .Y(n_412) );
AOI211xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_301), .B(n_311), .C(n_318), .Y(n_298) );
AND2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_310), .Y(n_342) );
INVx2_ASAP7_75t_L g357 ( .A(n_300), .Y(n_357) );
OR2x2_ASAP7_75t_L g395 ( .A(n_300), .B(n_358), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_300), .B(n_438), .Y(n_437) );
AOI211xp5_ASAP7_75t_SL g301 ( .A1(n_302), .A2(n_303), .B(n_305), .C(n_308), .Y(n_301) );
INVxp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_304), .B(n_342), .Y(n_341) );
OAI211xp5_ASAP7_75t_L g423 ( .A1(n_305), .A2(n_400), .B(n_424), .C(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_306), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g363 ( .A(n_307), .B(n_353), .Y(n_363) );
INVx1_ASAP7_75t_L g368 ( .A(n_307), .Y(n_368) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g311 ( .A(n_312), .B(n_315), .Y(n_311) );
INVxp33_ASAP7_75t_L g419 ( .A(n_313), .Y(n_419) );
AND2x2_ASAP7_75t_L g398 ( .A(n_314), .B(n_377), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_319), .A2(n_381), .B(n_382), .Y(n_380) );
OAI322xp33_ASAP7_75t_L g399 ( .A1(n_321), .A2(n_400), .A3(n_401), .B1(n_402), .B2(n_403), .C1(n_405), .C2(n_409), .Y(n_399) );
AOI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_326), .B1(n_331), .B2(n_335), .C(n_338), .Y(n_324) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_328), .B(n_330), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g376 ( .A(n_329), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g420 ( .A(n_333), .Y(n_420) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_336), .B(n_356), .Y(n_422) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g385 ( .A(n_345), .B(n_353), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_349), .B1(n_351), .B2(n_353), .C(n_354), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_349), .A2(n_366), .B1(n_370), .B2(n_371), .C(n_372), .Y(n_365) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_353), .B(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_356), .B1(n_359), .B2(n_362), .Y(n_354) );
OR2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx2_ASAP7_75t_SL g383 ( .A(n_358), .Y(n_383) );
INVxp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND5xp2_ASAP7_75t_L g364 ( .A(n_365), .B(n_386), .C(n_411), .D(n_421), .E(n_431), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
NOR4xp25_ASAP7_75t_L g439 ( .A(n_368), .B(n_374), .C(n_440), .D(n_441), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_371), .A2(n_432), .B1(n_434), .B2(n_436), .C(n_439), .Y(n_431) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
OAI322xp33_ASAP7_75t_L g387 ( .A1(n_381), .A2(n_388), .A3(n_389), .B1(n_390), .B2(n_391), .C1(n_393), .C2(n_397), .Y(n_387) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_399), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_394), .B(n_396), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g432 ( .A(n_407), .B(n_433), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVxp67_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g744 ( .A(n_444), .Y(n_744) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_448), .B(n_692), .Y(n_447) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_449), .B(n_627), .Y(n_448) );
NAND4xp25_ASAP7_75t_SL g449 ( .A(n_450), .B(n_572), .C(n_596), .D(n_619), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_514), .B1(n_544), .B2(n_556), .C(n_559), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_453), .B(n_487), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_453), .A2(n_473), .B1(n_515), .B2(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_453), .B(n_488), .Y(n_630) );
AND2x2_ASAP7_75t_L g649 ( .A(n_453), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_453), .B(n_633), .Y(n_719) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_473), .Y(n_453) );
AND2x2_ASAP7_75t_L g587 ( .A(n_454), .B(n_488), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_454), .B(n_602), .Y(n_601) );
OR2x2_ASAP7_75t_L g610 ( .A(n_454), .B(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g615 ( .A(n_454), .B(n_474), .Y(n_615) );
INVx2_ASAP7_75t_L g647 ( .A(n_454), .Y(n_647) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_454), .Y(n_691) );
AND2x2_ASAP7_75t_L g708 ( .A(n_454), .B(n_585), .Y(n_708) );
INVx5_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g626 ( .A(n_455), .B(n_585), .Y(n_626) );
AND2x4_ASAP7_75t_L g640 ( .A(n_455), .B(n_473), .Y(n_640) );
HB1xp67_ASAP7_75t_L g644 ( .A(n_455), .Y(n_644) );
AND2x2_ASAP7_75t_L g664 ( .A(n_455), .B(n_579), .Y(n_664) );
AND2x2_ASAP7_75t_L g714 ( .A(n_455), .B(n_489), .Y(n_714) );
AND2x2_ASAP7_75t_L g724 ( .A(n_455), .B(n_474), .Y(n_724) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_470), .Y(n_455) );
AOI21xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_461), .B(n_469), .Y(n_456) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx5_ASAP7_75t_L g479 ( .A(n_462), .Y(n_479) );
INVx2_ASAP7_75t_L g468 ( .A(n_466), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_468), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_L g520 ( .A1(n_468), .A2(n_497), .B(n_521), .C(n_522), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x2_ASAP7_75t_L g580 ( .A(n_473), .B(n_488), .Y(n_580) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_473), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_473), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g670 ( .A(n_473), .Y(n_670) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g558 ( .A(n_474), .B(n_503), .Y(n_558) );
AND2x2_ASAP7_75t_L g585 ( .A(n_474), .B(n_504), .Y(n_585) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_486), .Y(n_474) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_479), .B(n_480), .C(n_485), .Y(n_477) );
INVx2_ASAP7_75t_L g493 ( .A(n_479), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_479), .A2(n_485), .B(n_530), .C(n_531), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g498 ( .A(n_485), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_487), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_501), .Y(n_487) );
OR2x2_ASAP7_75t_L g611 ( .A(n_488), .B(n_502), .Y(n_611) );
AND2x2_ASAP7_75t_L g648 ( .A(n_488), .B(n_558), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_488), .B(n_579), .Y(n_659) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_488), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_488), .B(n_615), .Y(n_732) );
INVx5_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
AND2x2_ASAP7_75t_L g566 ( .A(n_489), .B(n_502), .Y(n_566) );
AND2x2_ASAP7_75t_L g682 ( .A(n_489), .B(n_577), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_489), .B(n_615), .Y(n_704) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_502), .Y(n_650) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_503), .Y(n_602) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx2_ASAP7_75t_L g579 ( .A(n_504), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_511), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_515), .B(n_592), .Y(n_711) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_516), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g563 ( .A(n_516), .B(n_564), .Y(n_563) );
INVx5_ASAP7_75t_SL g571 ( .A(n_516), .Y(n_571) );
OR2x2_ASAP7_75t_L g594 ( .A(n_516), .B(n_564), .Y(n_594) );
OR2x2_ASAP7_75t_L g604 ( .A(n_516), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g667 ( .A(n_516), .B(n_526), .Y(n_667) );
AND2x2_ASAP7_75t_SL g705 ( .A(n_516), .B(n_525), .Y(n_705) );
NOR4xp25_ASAP7_75t_L g726 ( .A(n_516), .B(n_647), .C(n_727), .D(n_728), .Y(n_726) );
AND2x2_ASAP7_75t_L g736 ( .A(n_516), .B(n_568), .Y(n_736) );
OR2x6_ASAP7_75t_L g516 ( .A(n_517), .B(n_523), .Y(n_516) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_557), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_525), .B(n_563), .Y(n_730) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_535), .Y(n_525) );
OR2x2_ASAP7_75t_L g570 ( .A(n_526), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_526), .B(n_546), .Y(n_589) );
INVxp67_ASAP7_75t_L g592 ( .A(n_526), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_526), .B(n_564), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_526), .B(n_536), .Y(n_658) );
AND2x2_ASAP7_75t_L g673 ( .A(n_526), .B(n_568), .Y(n_673) );
OR2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_536), .Y(n_702) );
OA21x2_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_534), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_535), .B(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_535), .B(n_571), .Y(n_710) );
OR2x2_ASAP7_75t_L g731 ( .A(n_535), .B(n_608), .Y(n_731) );
INVx1_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g545 ( .A(n_536), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g568 ( .A(n_536), .B(n_564), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_536), .B(n_546), .Y(n_583) );
AND2x2_ASAP7_75t_L g653 ( .A(n_536), .B(n_577), .Y(n_653) );
AND2x2_ASAP7_75t_L g687 ( .A(n_536), .B(n_571), .Y(n_687) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_537), .B(n_571), .Y(n_590) );
AND2x2_ASAP7_75t_L g618 ( .A(n_537), .B(n_546), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_544), .B(n_626), .Y(n_625) );
AOI221xp5_ASAP7_75t_L g685 ( .A1(n_545), .A2(n_633), .B1(n_669), .B2(n_686), .C(n_688), .Y(n_685) );
INVx5_ASAP7_75t_SL g564 ( .A(n_546), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B(n_550), .Y(n_547) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g584 ( .A1(n_557), .A2(n_585), .A3(n_586), .B1(n_588), .B2(n_591), .B3(n_595), .Y(n_584) );
OR2x2_ASAP7_75t_L g600 ( .A(n_557), .B(n_601), .Y(n_600) );
AOI322xp5_ASAP7_75t_L g709 ( .A1(n_557), .A2(n_626), .A3(n_633), .B1(n_710), .B2(n_711), .C1(n_712), .C2(n_715), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_557), .B(n_585), .Y(n_727) );
A2O1A1Ixp33_ASAP7_75t_SL g733 ( .A1(n_557), .A2(n_585), .B(n_734), .C(n_736), .Y(n_733) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_558), .A2(n_573), .B1(n_578), .B2(n_581), .C(n_584), .Y(n_572) );
INVx1_ASAP7_75t_L g665 ( .A(n_558), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_558), .B(n_714), .Y(n_713) );
OAI22xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_562), .B1(n_565), .B2(n_567), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g642 ( .A(n_563), .B(n_577), .Y(n_642) );
AND2x2_ASAP7_75t_L g700 ( .A(n_563), .B(n_701), .Y(n_700) );
OR2x2_ASAP7_75t_L g608 ( .A(n_564), .B(n_571), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_564), .B(n_577), .Y(n_636) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_566), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_566), .B(n_644), .Y(n_698) );
OAI321xp33_ASAP7_75t_L g717 ( .A1(n_566), .A2(n_639), .A3(n_718), .B1(n_719), .B2(n_720), .C(n_721), .Y(n_717) );
INVx1_ASAP7_75t_L g684 ( .A(n_567), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_568), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g623 ( .A(n_568), .B(n_571), .Y(n_623) );
AOI321xp33_ASAP7_75t_L g681 ( .A1(n_568), .A2(n_585), .A3(n_682), .B1(n_683), .B2(n_684), .C(n_685), .Y(n_681) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g598 ( .A(n_570), .B(n_583), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_571), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_571), .B(n_653), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_571), .B(n_657), .Y(n_694) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x4_ASAP7_75t_L g617 ( .A(n_575), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g582 ( .A(n_576), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g690 ( .A(n_577), .Y(n_690) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_580), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g613 ( .A(n_585), .Y(n_613) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_587), .B(n_622), .Y(n_671) );
OR2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
OR2x2_ASAP7_75t_L g635 ( .A(n_590), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g680 ( .A(n_590), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_591), .A2(n_638), .B1(n_641), .B2(n_643), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
OR2x2_ASAP7_75t_L g735 ( .A(n_594), .B(n_658), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B1(n_603), .B2(n_609), .C(n_612), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g633 ( .A(n_602), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_SL g679 ( .A(n_605), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_607), .B(n_657), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g674 ( .A1(n_607), .A2(n_675), .B(n_677), .Y(n_674) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g720 ( .A(n_608), .B(n_702), .Y(n_720) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_SL g622 ( .A(n_611), .Y(n_622) );
AOI21xp33_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_616), .Y(n_612) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g666 ( .A(n_618), .B(n_667), .Y(n_666) );
INVxp67_ASAP7_75t_L g728 ( .A(n_618), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_624), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_622), .B(n_640), .Y(n_676) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g697 ( .A(n_626), .Y(n_697) );
NAND5xp2_ASAP7_75t_L g627 ( .A(n_628), .B(n_645), .C(n_654), .D(n_674), .E(n_681), .Y(n_627) );
O2A1O1Ixp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_634), .C(n_637), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g669 ( .A(n_633), .Y(n_669) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_641), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g683 ( .A(n_643), .Y(n_683) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_649), .B(n_651), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_646), .A2(n_700), .B1(n_703), .B2(n_705), .C(n_706), .Y(n_699) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AOI321xp33_ASAP7_75t_L g654 ( .A1(n_647), .A2(n_655), .A3(n_659), .B1(n_660), .B2(n_666), .C(n_668), .Y(n_654) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g725 ( .A(n_659), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g660 ( .A(n_661), .B(n_665), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g677 ( .A(n_662), .B(n_678), .Y(n_677) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NOR2xp67_ASAP7_75t_SL g689 ( .A(n_663), .B(n_670), .Y(n_689) );
AOI321xp33_ASAP7_75t_SL g721 ( .A1(n_666), .A2(n_722), .A3(n_723), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_721) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B(n_671), .C(n_672), .Y(n_668) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_679), .B(n_687), .Y(n_716) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_691), .Y(n_688) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_717), .C(n_729), .Y(n_692) );
OAI211xp5_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_695), .B(n_699), .C(n_709), .Y(n_693) );
INVxp67_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OAI221xp5_ASAP7_75t_L g729 ( .A1(n_698), .A2(n_730), .B1(n_731), .B2(n_732), .C(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g718 ( .A(n_700), .Y(n_718) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_SL g722 ( .A(n_720), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
CKINVDCx14_ASAP7_75t_R g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
INVx3_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_759), .C(n_762), .Y(n_753) );
INVx1_ASAP7_75t_L g761 ( .A(n_755), .Y(n_761) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
endmodule