module fake_jpeg_28610_n_528 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_528);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_528;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx11_ASAP7_75t_SL g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_18),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_54),
.B(n_58),
.Y(n_136)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_56),
.Y(n_119)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_18),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_59),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_60),
.B(n_62),
.Y(n_112)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_24),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_24),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_68),
.B(n_71),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_73),
.B(n_79),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_37),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_0),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_37),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_96),
.Y(n_129)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_86),
.Y(n_148)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g125 ( 
.A(n_90),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_23),
.B(n_16),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_94),
.Y(n_153)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_23),
.B(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_95),
.Y(n_150)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_46),
.Y(n_97)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_97),
.Y(n_147)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_98),
.Y(n_145)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_24),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_103),
.B(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_34),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_39),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_77),
.A2(n_30),
.B1(n_31),
.B2(n_29),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_163),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_80),
.A2(n_29),
.B(n_16),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_109),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_117),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_78),
.A2(n_15),
.B(n_3),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_131),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_59),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_55),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_134),
.B(n_73),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_57),
.A2(n_39),
.B1(n_34),
.B2(n_40),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g174 ( 
.A(n_135),
.B(n_44),
.Y(n_174)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_137),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_139),
.B(n_67),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_90),
.A2(n_30),
.B1(n_31),
.B2(n_40),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_100),
.B1(n_101),
.B2(n_56),
.Y(n_176)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_83),
.B(n_38),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_45),
.Y(n_167)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_91),
.A2(n_31),
.B1(n_30),
.B2(n_28),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_99),
.B1(n_53),
.B2(n_86),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_61),
.A2(n_31),
.B1(n_45),
.B2(n_35),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g164 ( 
.A(n_129),
.B(n_65),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_154),
.C(n_157),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_89),
.B1(n_93),
.B2(n_95),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_111),
.Y(n_166)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_166),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_167),
.B(n_173),
.Y(n_236)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_169),
.Y(n_264)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_124),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_171),
.B(n_182),
.Y(n_253)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_160),
.Y(n_172)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_172),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_110),
.A2(n_96),
.B(n_35),
.C(n_33),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_174),
.B(n_178),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_176),
.A2(n_162),
.B1(n_63),
.B2(n_74),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_103),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_50),
.B(n_32),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_183),
.Y(n_232)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

NAND2xp33_ASAP7_75t_SL g182 ( 
.A(n_144),
.B(n_88),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_188),
.Y(n_238)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_108),
.B(n_66),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_185),
.B(n_213),
.Y(n_250)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_209),
.B1(n_69),
.B2(n_72),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_106),
.Y(n_191)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_191),
.Y(n_251)
);

BUFx4f_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

BUFx2_ASAP7_75t_SL g255 ( 
.A(n_192),
.Y(n_255)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_195),
.B(n_207),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g196 ( 
.A(n_147),
.Y(n_196)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_105),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_198),
.Y(n_242)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_150),
.Y(n_201)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_204),
.Y(n_229)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_141),
.B(n_71),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_136),
.B(n_68),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_210),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_135),
.A2(n_85),
.B1(n_81),
.B2(n_82),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_112),
.B(n_64),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_211),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_125),
.A2(n_36),
.B1(n_28),
.B2(n_20),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_159),
.B(n_32),
.Y(n_213)
);

NAND2xp33_ASAP7_75t_SL g214 ( 
.A(n_159),
.B(n_32),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_214),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_147),
.B(n_28),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_216),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_116),
.B(n_28),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_132),
.B(n_28),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_218),
.Y(n_243)
);

INVx6_ASAP7_75t_SL g219 ( 
.A(n_123),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_219),
.Y(n_260)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_220),
.Y(n_246)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_142),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_221),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_231),
.B(n_192),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_193),
.A2(n_154),
.B1(n_148),
.B2(n_123),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_233),
.A2(n_256),
.B(n_49),
.Y(n_299)
);

AO22x2_ASAP7_75t_L g234 ( 
.A1(n_185),
.A2(n_174),
.B1(n_187),
.B2(n_214),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g279 ( 
.A1(n_234),
.A2(n_171),
.B1(n_201),
.B2(n_44),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_146),
.B1(n_127),
.B2(n_133),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_193),
.A2(n_148),
.B1(n_49),
.B2(n_50),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_205),
.A2(n_151),
.B1(n_158),
.B2(n_119),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_263),
.B1(n_152),
.B2(n_126),
.Y(n_282)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_173),
.A2(n_185),
.B1(n_205),
.B2(n_164),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_258),
.A2(n_180),
.B1(n_181),
.B2(n_199),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_161),
.B1(n_126),
.B2(n_146),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_261),
.A2(n_169),
.B1(n_191),
.B2(n_204),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_164),
.B(n_158),
.C(n_151),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_269),
.C(n_206),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_175),
.B(n_84),
.C(n_76),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_185),
.B(n_182),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_270),
.A2(n_286),
.B1(n_292),
.B2(n_296),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx3_ASAP7_75t_SL g345 ( 
.A(n_271),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_238),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_272),
.Y(n_334)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_254),
.Y(n_273)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_288),
.Y(n_323)
);

O2A1O1Ixp33_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_192),
.B(n_190),
.C(n_217),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_275),
.Y(n_335)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_277),
.Y(n_321)
);

AND2x6_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_202),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_278),
.B(n_280),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_279),
.A2(n_284),
.B(n_297),
.Y(n_328)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_177),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_281),
.B(n_283),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_282),
.A2(n_266),
.B1(n_227),
.B2(n_256),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_232),
.B(n_186),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_295),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_236),
.B(n_243),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_291),
.Y(n_333)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_249),
.Y(n_290)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_259),
.A2(n_133),
.B1(n_127),
.B2(n_152),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_240),
.Y(n_293)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_293),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_294),
.B(n_303),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_203),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_244),
.A2(n_121),
.B1(n_155),
.B2(n_161),
.Y(n_296)
);

OR2x4_ASAP7_75t_L g297 ( 
.A(n_234),
.B(n_253),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_222),
.A2(n_121),
.B1(n_155),
.B2(n_194),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_302),
.B1(n_311),
.B2(n_296),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_299),
.A2(n_312),
.B1(n_172),
.B2(n_200),
.Y(n_350)
);

INVx6_ASAP7_75t_SL g300 ( 
.A(n_268),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_301),
.Y(n_343)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_254),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_222),
.A2(n_166),
.B1(n_170),
.B2(n_189),
.Y(n_302)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_268),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_267),
.B(n_200),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_304),
.B(n_306),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_260),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_307),
.Y(n_346)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

OR2x4_ASAP7_75t_L g308 ( 
.A(n_234),
.B(n_50),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_308),
.A2(n_49),
.B(n_228),
.Y(n_351)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_309),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_243),
.B(n_186),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_310),
.B(n_242),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_262),
.A2(n_231),
.B1(n_234),
.B2(n_239),
.Y(n_311)
);

INVx5_ASAP7_75t_SL g312 ( 
.A(n_260),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_247),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_314),
.B(n_326),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_297),
.A2(n_239),
.B1(n_253),
.B2(n_233),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_315),
.A2(n_317),
.B1(n_319),
.B2(n_324),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_304),
.B1(n_279),
.B2(n_295),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_279),
.A2(n_253),
.B1(n_302),
.B2(n_298),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_320),
.B(n_271),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_322),
.A2(n_286),
.B1(n_292),
.B2(n_277),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_285),
.A2(n_269),
.B1(n_257),
.B2(n_263),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_265),
.C(n_246),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_338),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_223),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_327),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_278),
.A2(n_227),
.B1(n_266),
.B2(n_229),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_329),
.A2(n_332),
.B1(n_342),
.B2(n_300),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_275),
.A2(n_252),
.B1(n_226),
.B2(n_237),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_299),
.A2(n_264),
.B(n_237),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_337),
.B(n_340),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_273),
.B(n_242),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_235),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_312),
.A2(n_252),
.B1(n_264),
.B2(n_168),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_332),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_351),
.Y(n_376)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_343),
.Y(n_352)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_353),
.B(n_372),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_346),
.B(n_309),
.Y(n_355)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_355),
.Y(n_404)
);

OAI21xp33_ASAP7_75t_L g357 ( 
.A1(n_327),
.A2(n_305),
.B(n_280),
.Y(n_357)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_371),
.B(n_315),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_334),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_367),
.Y(n_386)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_343),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_359),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_340),
.B(n_306),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_365),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_336),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_363),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_339),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_369),
.B1(n_329),
.B2(n_321),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_345),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_341),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_368),
.A2(n_378),
.B1(n_316),
.B2(n_317),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_335),
.A2(n_290),
.B1(n_276),
.B2(n_287),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_375),
.Y(n_402)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_330),
.B(n_303),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_307),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_373),
.A2(n_382),
.B1(n_337),
.B2(n_344),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_331),
.B(n_280),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_225),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_377),
.B(n_384),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_335),
.A2(n_225),
.B1(n_248),
.B2(n_246),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_320),
.A2(n_235),
.B(n_248),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_379),
.A2(n_378),
.B(n_382),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_349),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_380),
.B(n_381),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_318),
.B(n_349),
.Y(n_381)
);

OAI22x1_ASAP7_75t_L g382 ( 
.A1(n_328),
.A2(n_291),
.B1(n_202),
.B2(n_149),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_318),
.B(n_177),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_383),
.B(n_385),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_319),
.B(n_230),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_341),
.B(n_230),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_366),
.A2(n_322),
.B1(n_316),
.B2(n_328),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_387),
.A2(n_393),
.B1(n_398),
.B2(n_408),
.Y(n_433)
);

AOI21xp33_ASAP7_75t_L g441 ( 
.A1(n_389),
.A2(n_44),
.B(n_5),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_385),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_391),
.B(n_412),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_356),
.B(n_326),
.Y(n_392)
);

NAND3xp33_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_365),
.C(n_3),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_394),
.A2(n_376),
.B1(n_365),
.B2(n_370),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_395),
.A2(n_401),
.B1(n_405),
.B2(n_411),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_325),
.C(n_314),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_406),
.C(n_374),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_366),
.A2(n_324),
.B1(n_323),
.B2(n_348),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_373),
.A2(n_323),
.B1(n_338),
.B2(n_344),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_373),
.A2(n_348),
.B1(n_345),
.B2(n_313),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_351),
.C(n_313),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_355),
.B(n_321),
.Y(n_407)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_407),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_384),
.A2(n_345),
.B1(n_224),
.B2(n_221),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_360),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_149),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_364),
.A2(n_224),
.B1(n_220),
.B2(n_211),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_352),
.A2(n_359),
.B1(n_379),
.B2(n_353),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_369),
.A2(n_145),
.B1(n_41),
.B2(n_4),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_413),
.A2(n_362),
.B1(n_36),
.B2(n_20),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_36),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_415),
.A2(n_44),
.B(n_5),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_439),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_399),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_418),
.B(n_434),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_361),
.C(n_372),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_419),
.B(n_440),
.C(n_403),
.Y(n_453)
);

OAI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_404),
.A2(n_368),
.B1(n_371),
.B2(n_367),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_420),
.A2(n_422),
.B1(n_427),
.B2(n_431),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_437),
.B(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_426),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_428),
.B(n_429),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_410),
.B(n_36),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_401),
.B(n_36),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_436),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_396),
.A2(n_20),
.B1(n_3),
.B2(n_5),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_399),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_386),
.B(n_2),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_390),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_48),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_438),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_398),
.B(n_409),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_48),
.C(n_44),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_396),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_442),
.A2(n_393),
.B1(n_408),
.B2(n_413),
.Y(n_463)
);

FAx1_ASAP7_75t_L g444 ( 
.A(n_423),
.B(n_412),
.CI(n_415),
.CON(n_444),
.SN(n_444)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_444),
.B(n_454),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_419),
.B(n_417),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_455),
.C(n_457),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_432),
.B(n_386),
.Y(n_449)
);

CKINVDCx14_ASAP7_75t_R g479 ( 
.A(n_449),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_423),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_450),
.Y(n_469)
);

XNOR2x1_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_456),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_387),
.C(n_388),
.Y(n_455)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_395),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_388),
.C(n_404),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_391),
.C(n_416),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_421),
.C(n_424),
.Y(n_466)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_426),
.Y(n_461)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_461),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_433),
.A2(n_394),
.B1(n_411),
.B2(n_416),
.Y(n_462)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_462),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_463),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_475),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_444),
.A2(n_437),
.B(n_438),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_458),
.B(n_10),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_SL g468 ( 
.A(n_445),
.B(n_414),
.C(n_407),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_468),
.B(n_473),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_460),
.A2(n_433),
.B1(n_405),
.B2(n_403),
.Y(n_471)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_456),
.B(n_429),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_472),
.B(n_476),
.Y(n_481)
);

AOI322xp5_ASAP7_75t_SL g473 ( 
.A1(n_451),
.A2(n_442),
.A3(n_392),
.B1(n_431),
.B2(n_430),
.C1(n_402),
.C2(n_427),
.Y(n_473)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_447),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_440),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_463),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_480),
.A2(n_452),
.B1(n_459),
.B2(n_455),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_446),
.C(n_443),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_484),
.C(n_489),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_479),
.B(n_466),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_486),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_443),
.C(n_453),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_465),
.B(n_457),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_470),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_448),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_490),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_478),
.B(n_444),
.Y(n_490)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_491),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_458),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_472),
.Y(n_503)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_469),
.B(n_9),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g504 ( 
.A(n_495),
.Y(n_504)
);

OAI21x1_ASAP7_75t_L g496 ( 
.A1(n_488),
.A2(n_478),
.B(n_485),
.Y(n_496)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_496),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_502),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_490),
.A2(n_467),
.B(n_469),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_500),
.A2(n_481),
.B(n_11),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_474),
.C(n_471),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_505),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_474),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_475),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_506),
.B(n_507),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_493),
.B1(n_494),
.B2(n_468),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_511),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_470),
.B1(n_480),
.B2(n_492),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_512),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_499),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_515),
.A2(n_503),
.B1(n_497),
.B2(n_481),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_498),
.C(n_502),
.Y(n_518)
);

AO21x1_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_508),
.B(n_505),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_SL g519 ( 
.A1(n_517),
.A2(n_499),
.B(n_514),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_519),
.B(n_520),
.Y(n_523)
);

AOI321xp33_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_515),
.A3(n_513),
.B1(n_516),
.B2(n_13),
.C(n_10),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_10),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_524),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_523),
.C(n_12),
.Y(n_526)
);

O2A1O1Ixp33_ASAP7_75t_SL g527 ( 
.A1(n_526),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_527),
.A2(n_48),
.B1(n_504),
.B2(n_525),
.Y(n_528)
);


endmodule