module real_jpeg_2683_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_1),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_2),
.A2(n_34),
.B1(n_36),
.B2(n_39),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_4),
.A2(n_68),
.B1(n_69),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_76),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_76),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_5),
.A2(n_68),
.B1(n_69),
.B2(n_82),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_5),
.A2(n_34),
.B1(n_36),
.B2(n_82),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_6),
.A2(n_83),
.B1(n_86),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_6),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_97),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_6),
.A2(n_28),
.B1(n_29),
.B2(n_97),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_97),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_8),
.A2(n_83),
.B1(n_86),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_8),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_8),
.A2(n_68),
.B1(n_69),
.B2(n_112),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_112),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_112),
.Y(n_222)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_11),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_11),
.A2(n_60),
.B1(n_68),
.B2(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_86),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_15),
.B(n_113),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_15),
.A2(n_67),
.B(n_68),
.C(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_15),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_15),
.B(n_73),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_15),
.A2(n_68),
.B1(n_69),
.B2(n_162),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_31),
.C(n_34),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_162),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_15),
.B(n_46),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_15),
.B(n_61),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_139),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_138),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_21),
.B(n_114),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_99),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_24),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_25),
.A2(n_33),
.B1(n_155),
.B2(n_189),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_25),
.A2(n_157),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_26),
.A2(n_38),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_26),
.A2(n_59),
.B1(n_61),
.B2(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_26),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_26),
.B(n_158),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_28),
.A2(n_29),
.B1(n_67),
.B2(n_74),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_28),
.A2(n_74),
.B(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_29),
.B(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_33),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_33),
.A2(n_178),
.B(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_34),
.B(n_218),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B(n_47),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_43),
.A2(n_46),
.B1(n_56),
.B2(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_43),
.A2(n_162),
.B(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_44),
.A2(n_45),
.B1(n_48),
.B2(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_44),
.A2(n_45),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_44),
.A2(n_45),
.B1(n_136),
.B2(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_44),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_44),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_44),
.A2(n_45),
.B1(n_193),
.B2(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_45),
.A2(n_152),
.B(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_45),
.B(n_166),
.Y(n_195)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_46),
.A2(n_165),
.B(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_62),
.B1(n_63),
.B2(n_98),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_53),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_61),
.B(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_79),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_65),
.A2(n_127),
.B(n_129),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_65),
.A2(n_129),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_66),
.B(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_66),
.A2(n_73),
.B1(n_128),
.B2(n_146),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B(n_72),
.C(n_73),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_69),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_68),
.A2(n_83),
.A3(n_90),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_69),
.B(n_92),
.Y(n_133)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_73),
.B(n_109),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_77),
.B(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_77),
.A2(n_108),
.B(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_87),
.B(n_94),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_88),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_86),
.B1(n_90),
.B2(n_92),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_83),
.A2(n_87),
.B(n_162),
.C(n_171),
.Y(n_170)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_93),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_90),
.Y(n_92)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_95),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.C(n_110),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_101),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_102),
.B(n_104),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_103),
.Y(n_177)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_110),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_111),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_119),
.C(n_121),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_115),
.B(n_119),
.Y(n_242)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_121),
.B(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.C(n_130),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_122),
.B(n_126),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_130),
.B(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI31xp33_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_239),
.A3(n_249),
.B(n_254),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_183),
.B(n_238),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_167),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_142),
.B(n_167),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_153),
.C(n_159),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_143),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_148),
.C(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_153),
.B(n_159),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_163),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_179),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_168),
.B(n_180),
.C(n_182),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_169),
.B(n_174),
.C(n_175),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_233),
.B(n_237),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_202),
.B(n_232),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_196),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_196),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_190),
.C(n_191),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_192),
.B1(n_211),
.B2(n_213),
.Y(n_210)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_214),
.B(n_231),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_210),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_211),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_225),
.B(n_230),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_220),
.B(n_224),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_221),
.B(n_223),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_222),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_228),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI21xp33_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_241),
.B(n_243),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_246),
.A2(n_247),
.B1(n_248),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_253),
.Y(n_255)
);


endmodule