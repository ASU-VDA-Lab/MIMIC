module fake_aes_3691_n_476 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_476);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_476;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_67;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
HB1xp67_ASAP7_75t_L g65 ( .A(n_50), .Y(n_65) );
INVx1_ASAP7_75t_L g66 ( .A(n_43), .Y(n_66) );
INVxp67_ASAP7_75t_SL g67 ( .A(n_19), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_9), .Y(n_68) );
INVxp33_ASAP7_75t_SL g69 ( .A(n_29), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_62), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_27), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_13), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_5), .Y(n_73) );
CKINVDCx20_ASAP7_75t_R g74 ( .A(n_7), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_24), .Y(n_75) );
INVxp33_ASAP7_75t_L g76 ( .A(n_45), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_25), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_64), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_6), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_51), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_0), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_55), .B(n_9), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_13), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_14), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_35), .Y(n_85) );
BUFx10_ASAP7_75t_L g86 ( .A(n_38), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_33), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_53), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_20), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_63), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_18), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_26), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_57), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
BUFx3_ASAP7_75t_L g96 ( .A(n_23), .Y(n_96) );
BUFx3_ASAP7_75t_L g97 ( .A(n_41), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_3), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_65), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_85), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_85), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_83), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_99), .B(n_0), .Y(n_104) );
NAND2xp33_ASAP7_75t_R g105 ( .A(n_69), .B(n_39), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_83), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_99), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_88), .Y(n_108) );
BUFx2_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_94), .B(n_1), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_94), .B(n_1), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_89), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_68), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_66), .Y(n_115) );
OR2x6_ASAP7_75t_L g116 ( .A(n_72), .B(n_2), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_72), .B(n_3), .Y(n_117) );
INVx2_ASAP7_75t_L g118 ( .A(n_89), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_66), .Y(n_119) );
NAND2xp33_ASAP7_75t_SL g120 ( .A(n_76), .B(n_4), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_73), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_101), .Y(n_124) );
BUFx3_ASAP7_75t_L g125 ( .A(n_118), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_108), .Y(n_126) );
INVx4_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_115), .B(n_71), .Y(n_128) );
AND2x6_ASAP7_75t_L g129 ( .A(n_104), .B(n_96), .Y(n_129) );
NAND2xp5_ASAP7_75t_SL g130 ( .A(n_100), .B(n_86), .Y(n_130) );
INVxp33_ASAP7_75t_L g131 ( .A(n_109), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_104), .B(n_96), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_113), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_102), .Y(n_134) );
AO22x2_ASAP7_75t_L g135 ( .A1(n_104), .A2(n_98), .B1(n_71), .B2(n_75), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_109), .B(n_86), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_117), .A2(n_73), .B1(n_79), .B2(n_81), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_113), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_107), .B(n_86), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_116), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_115), .B(n_70), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
XOR2xp5_ASAP7_75t_L g145 ( .A(n_108), .B(n_74), .Y(n_145) );
INVxp67_ASAP7_75t_SL g146 ( .A(n_119), .Y(n_146) );
NAND2xp33_ASAP7_75t_SL g147 ( .A(n_105), .B(n_79), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_135), .A2(n_116), .B1(n_117), .B2(n_120), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_125), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_135), .A2(n_117), .B1(n_120), .B2(n_119), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_123), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_124), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_146), .B(n_110), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_141), .B(n_114), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_124), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_127), .B(n_121), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_125), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_135), .A2(n_122), .B1(n_118), .B2(n_111), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_141), .B(n_112), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_127), .Y(n_164) );
INVx5_ASAP7_75t_L g165 ( .A(n_129), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_143), .A2(n_122), .B(n_90), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g167 ( .A(n_131), .B(n_78), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_133), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_136), .B(n_86), .Y(n_169) );
CKINVDCx8_ASAP7_75t_R g170 ( .A(n_126), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_133), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_134), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_133), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_136), .B(n_103), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_145), .Y(n_176) );
INVx1_ASAP7_75t_SL g177 ( .A(n_145), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_127), .Y(n_178) );
AND2x6_ASAP7_75t_L g179 ( .A(n_142), .B(n_75), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_142), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
BUFx12f_ASAP7_75t_L g182 ( .A(n_179), .Y(n_182) );
CKINVDCx11_ASAP7_75t_R g183 ( .A(n_170), .Y(n_183) );
AOI21xp33_ASAP7_75t_L g184 ( .A1(n_167), .A2(n_144), .B(n_142), .Y(n_184) );
BUFx2_ASAP7_75t_L g185 ( .A(n_157), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_169), .B(n_138), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_151), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_157), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_157), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
AOI21x1_ASAP7_75t_L g191 ( .A1(n_166), .A2(n_135), .B(n_128), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx5_ASAP7_75t_SL g193 ( .A(n_157), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g194 ( .A1(n_170), .A2(n_144), .B1(n_142), .B2(n_128), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
INVx2_ASAP7_75t_SL g199 ( .A(n_165), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_169), .B(n_144), .Y(n_200) );
INVx4_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_156), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_165), .B(n_144), .Y(n_204) );
OR2x6_ASAP7_75t_L g205 ( .A(n_171), .B(n_135), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_148), .A2(n_130), .B1(n_139), .B2(n_92), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_150), .A2(n_129), .B1(n_132), .B2(n_147), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_162), .A2(n_140), .B(n_139), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_163), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_176), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_183), .Y(n_213) );
BUFx4f_ASAP7_75t_SL g214 ( .A(n_211), .Y(n_214) );
OR2x2_ASAP7_75t_L g215 ( .A(n_186), .B(n_177), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_192), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_181), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_SL g218 ( .A1(n_192), .A2(n_163), .B(n_173), .C(n_159), .Y(n_218) );
INVx2_ASAP7_75t_SL g219 ( .A(n_182), .Y(n_219) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_205), .A2(n_161), .B1(n_173), .B2(n_155), .Y(n_220) );
AO31x2_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_140), .A3(n_77), .B(n_80), .Y(n_221) );
INVx2_ASAP7_75t_SL g222 ( .A(n_182), .Y(n_222) );
AOI22xp33_ASAP7_75t_SL g223 ( .A1(n_205), .A2(n_179), .B1(n_171), .B2(n_132), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_210), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_185), .A2(n_129), .B1(n_132), .B2(n_179), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_210), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_210), .Y(n_228) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_205), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_200), .B(n_185), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_205), .Y(n_231) );
NOR2xp33_ASAP7_75t_SL g232 ( .A(n_205), .B(n_179), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_188), .A2(n_175), .B1(n_154), .B2(n_178), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_189), .B(n_164), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_187), .Y(n_235) );
OAI21xp5_ASAP7_75t_L g236 ( .A1(n_209), .A2(n_158), .B(n_149), .Y(n_236) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_140), .B(n_77), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g238 ( .A(n_193), .Y(n_238) );
BUFx4f_ASAP7_75t_L g239 ( .A(n_231), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_216), .B(n_187), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_216), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_215), .A2(n_207), .B1(n_132), .B2(n_129), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
OAI221xp5_ASAP7_75t_L g244 ( .A1(n_215), .A2(n_208), .B1(n_184), .B2(n_189), .C(n_206), .Y(n_244) );
OR2x6_ASAP7_75t_L g245 ( .A(n_231), .B(n_195), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_228), .Y(n_246) );
OAI221xp5_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_206), .B1(n_190), .B2(n_197), .C(n_106), .Y(n_247) );
OAI221xp5_ASAP7_75t_SL g248 ( .A1(n_235), .A2(n_194), .B1(n_95), .B2(n_81), .C(n_91), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_217), .B(n_190), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_230), .A2(n_132), .B1(n_129), .B2(n_179), .Y(n_250) );
CKINVDCx9p33_ASAP7_75t_R g251 ( .A(n_214), .Y(n_251) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_236), .A2(n_226), .B(n_224), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_226), .B(n_195), .Y(n_254) );
AOI22xp33_ASAP7_75t_SL g255 ( .A1(n_232), .A2(n_193), .B1(n_179), .B2(n_197), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_227), .Y(n_256) );
OAI221xp5_ASAP7_75t_L g257 ( .A1(n_223), .A2(n_202), .B1(n_191), .B2(n_95), .C(n_84), .Y(n_257) );
OAI221xp5_ASAP7_75t_SL g258 ( .A1(n_225), .A2(n_91), .B1(n_84), .B2(n_87), .C(n_80), .Y(n_258) );
OAI22xp33_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_202), .B1(n_164), .B2(n_180), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_241), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_248), .B(n_213), .C(n_82), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_253), .A2(n_218), .B(n_237), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_239), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_240), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_257), .A2(n_233), .B1(n_238), .B2(n_132), .Y(n_265) );
AND2x4_ASAP7_75t_L g266 ( .A(n_245), .B(n_221), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_244), .A2(n_238), .B1(n_129), .B2(n_132), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_241), .B(n_237), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_245), .B(n_221), .Y(n_269) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_239), .A2(n_193), .B1(n_237), .B2(n_222), .Y(n_270) );
OAI31xp33_ASAP7_75t_L g271 ( .A1(n_258), .A2(n_219), .A3(n_222), .B(n_90), .Y(n_271) );
NAND3xp33_ASAP7_75t_L g272 ( .A(n_247), .B(n_237), .C(n_113), .Y(n_272) );
AOI33xp33_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_87), .A3(n_93), .B1(n_98), .B2(n_219), .B3(n_8), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_253), .B(n_221), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_252), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_243), .B(n_221), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_252), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_243), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_253), .B(n_221), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_246), .B(n_193), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_260), .Y(n_281) );
OAI31xp33_ASAP7_75t_L g282 ( .A1(n_271), .A2(n_259), .A3(n_249), .B(n_246), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_264), .B(n_240), .Y(n_284) );
OAI31xp33_ASAP7_75t_L g285 ( .A1(n_271), .A2(n_249), .A3(n_242), .B(n_254), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_264), .B(n_254), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_260), .B(n_278), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g288 ( .A(n_263), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_278), .B(n_213), .Y(n_289) );
INVx4_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_276), .B(n_245), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_263), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g294 ( .A1(n_261), .A2(n_239), .B1(n_255), .B2(n_245), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_274), .B(n_245), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVxp33_ASAP7_75t_L g297 ( .A(n_280), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_275), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_265), .A2(n_239), .B1(n_249), .B2(n_193), .Y(n_299) );
NOR3xp33_ASAP7_75t_L g300 ( .A(n_273), .B(n_93), .C(n_67), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_275), .Y(n_301) );
AOI21xp33_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_256), .B(n_249), .Y(n_302) );
AOI331xp33_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_251), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_10), .C1(n_11), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_266), .B(n_96), .Y(n_304) );
OAI221xp5_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_250), .B1(n_97), .B2(n_113), .C(n_252), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_277), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_280), .B(n_4), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_272), .A2(n_97), .B1(n_252), .B2(n_180), .C(n_178), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_274), .B(n_97), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_274), .B(n_10), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_283), .B(n_279), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_296), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_288), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_281), .Y(n_314) );
INVx2_ASAP7_75t_SL g315 ( .A(n_288), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_283), .B(n_279), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_284), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_283), .B(n_279), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_284), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_281), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_292), .B(n_277), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_304), .B(n_266), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_291), .B(n_277), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_286), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_292), .B(n_266), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_295), .B(n_269), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_301), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_310), .B(n_269), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_291), .B(n_269), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_295), .B(n_269), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_309), .B(n_269), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_296), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_304), .B(n_268), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_309), .B(n_268), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_300), .A2(n_280), .B1(n_272), .B2(n_262), .C(n_137), .Y(n_336) );
AND2x4_ASAP7_75t_L g337 ( .A(n_304), .B(n_262), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_301), .B(n_11), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_304), .B(n_12), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_310), .B(n_12), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_306), .B(n_15), .Y(n_341) );
NAND3xp33_ASAP7_75t_L g342 ( .A(n_289), .B(n_133), .C(n_137), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_298), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_298), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_297), .B(n_15), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_302), .B(n_16), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_290), .B(n_293), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_293), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_307), .B(n_16), .Y(n_351) );
AOI22x1_ASAP7_75t_L g352 ( .A1(n_313), .A2(n_303), .B1(n_282), .B2(n_285), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_315), .Y(n_353) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_320), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_317), .B(n_299), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g358 ( .A1(n_319), .A2(n_294), .B(n_305), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_328), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_324), .B(n_282), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_328), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_344), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_325), .B(n_285), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_312), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_351), .A2(n_308), .B1(n_129), .B2(n_132), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_335), .B(n_338), .Y(n_367) );
OAI21xp33_ASAP7_75t_L g368 ( .A1(n_340), .A2(n_133), .B(n_137), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_321), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g370 ( .A(n_346), .B(n_17), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_329), .B(n_21), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_311), .B(n_22), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_338), .B(n_129), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_333), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_330), .Y(n_376) );
OAI332xp33_ASAP7_75t_L g377 ( .A1(n_340), .A2(n_159), .A3(n_158), .B1(n_149), .B2(n_199), .B3(n_160), .C1(n_172), .C2(n_179), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_339), .A2(n_348), .B(n_347), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_341), .B(n_28), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_341), .B(n_30), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_323), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_343), .Y(n_382) );
OAI322xp33_ASAP7_75t_L g383 ( .A1(n_339), .A2(n_326), .A3(n_331), .B1(n_327), .B2(n_332), .C1(n_315), .C2(n_348), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_332), .A2(n_201), .B1(n_203), .B2(n_199), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_316), .B(n_31), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_349), .B(n_32), .Y(n_386) );
NOR3xp33_ASAP7_75t_L g387 ( .A(n_342), .B(n_234), .C(n_203), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_318), .B(n_350), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_318), .B(n_36), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_322), .B(n_37), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_371), .B(n_334), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_376), .B(n_334), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_353), .B(n_322), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_381), .B(n_331), .Y(n_394) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_360), .B(n_336), .C(n_327), .D(n_326), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_366), .B(n_334), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_388), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_387), .B(n_337), .Y(n_398) );
AOI321xp33_ASAP7_75t_L g399 ( .A1(n_363), .A2(n_337), .A3(n_345), .B1(n_234), .B2(n_204), .C(n_160), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_356), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_369), .B(n_337), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_357), .B(n_40), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_352), .A2(n_42), .B(n_44), .Y(n_404) );
OAI21xp5_ASAP7_75t_L g405 ( .A1(n_368), .A2(n_204), .B(n_203), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_367), .B(n_46), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_354), .Y(n_407) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_358), .A2(n_204), .B1(n_201), .B2(n_158), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_390), .B(n_212), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_354), .B(n_47), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_355), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_383), .B(n_48), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_364), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_378), .B(n_49), .Y(n_416) );
AND3x1_ASAP7_75t_L g417 ( .A(n_370), .B(n_52), .C(n_54), .Y(n_417) );
NAND3x1_ASAP7_75t_L g418 ( .A(n_373), .B(n_56), .C(n_58), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_364), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_375), .Y(n_420) );
XOR2x2_ASAP7_75t_L g421 ( .A(n_390), .B(n_59), .Y(n_421) );
OAI32xp33_ASAP7_75t_L g422 ( .A1(n_386), .A2(n_201), .A3(n_159), .B1(n_60), .B2(n_61), .Y(n_422) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_365), .A2(n_198), .B(n_196), .Y(n_423) );
OAI31xp33_ASAP7_75t_L g424 ( .A1(n_384), .A2(n_172), .A3(n_196), .B(n_198), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_382), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_382), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_SL g427 ( .A1(n_379), .A2(n_196), .B(n_212), .C(n_168), .Y(n_427) );
NOR2xp33_ASAP7_75t_SL g428 ( .A(n_385), .B(n_212), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_372), .A2(n_196), .B1(n_168), .B2(n_174), .Y(n_429) );
XNOR2x1_ASAP7_75t_L g430 ( .A(n_389), .B(n_380), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_374), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g432 ( .A1(n_377), .A2(n_168), .B(n_174), .C(n_352), .Y(n_432) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_352), .A2(n_174), .B(n_378), .C(n_313), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_360), .A2(n_358), .B1(n_351), .B2(n_363), .Y(n_434) );
AOI211xp5_ASAP7_75t_SL g435 ( .A1(n_383), .A2(n_358), .B(n_368), .C(n_378), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_356), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_371), .B(n_376), .Y(n_437) );
XOR2x2_ASAP7_75t_L g438 ( .A(n_353), .B(n_313), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_356), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_356), .Y(n_440) );
XNOR2xp5_ASAP7_75t_L g441 ( .A(n_353), .B(n_213), .Y(n_441) );
XOR2xp5_ASAP7_75t_L g442 ( .A(n_441), .B(n_438), .Y(n_442) );
OAI21xp5_ASAP7_75t_SL g443 ( .A1(n_435), .A2(n_433), .B(n_432), .Y(n_443) );
BUFx2_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
AOI221xp5_ASAP7_75t_L g445 ( .A1(n_397), .A2(n_434), .B1(n_413), .B2(n_395), .C(n_436), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_420), .Y(n_446) );
NOR4xp25_ASAP7_75t_L g447 ( .A(n_404), .B(n_418), .C(n_399), .D(n_398), .Y(n_447) );
AOI22x1_ASAP7_75t_L g448 ( .A1(n_421), .A2(n_405), .B1(n_393), .B2(n_403), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_440), .A2(n_439), .B1(n_402), .B2(n_400), .C(n_437), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_411), .Y(n_450) );
XOR2xp5_ASAP7_75t_L g451 ( .A(n_430), .B(n_421), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_419), .A2(n_415), .B1(n_412), .B2(n_414), .C(n_401), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_398), .A2(n_408), .B1(n_391), .B2(n_396), .Y(n_453) );
XNOR2xp5_ASAP7_75t_L g454 ( .A(n_417), .B(n_394), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_391), .B(n_392), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_448), .A2(n_409), .B1(n_423), .B2(n_431), .Y(n_456) );
OAI211xp5_ASAP7_75t_SL g457 ( .A1(n_443), .A2(n_423), .B(n_406), .C(n_424), .Y(n_457) );
INVxp33_ASAP7_75t_SL g458 ( .A(n_442), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_451), .B(n_416), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_444), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_443), .B(n_416), .C(n_428), .D(n_424), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_447), .A2(n_422), .B(n_429), .C(n_427), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g463 ( .A(n_461), .B(n_450), .Y(n_463) );
INVxp33_ASAP7_75t_SL g464 ( .A(n_459), .Y(n_464) );
NOR4xp25_ASAP7_75t_L g465 ( .A(n_457), .B(n_445), .C(n_449), .D(n_452), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_462), .B(n_453), .C(n_454), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_460), .A2(n_446), .B1(n_455), .B2(n_426), .C1(n_425), .C2(n_410), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_463), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_466), .Y(n_469) );
OA22x2_ASAP7_75t_L g470 ( .A1(n_465), .A2(n_456), .B1(n_464), .B2(n_458), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_469), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_468), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_472), .Y(n_473) );
OR2x6_ASAP7_75t_L g474 ( .A(n_473), .B(n_470), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_474), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_475), .A2(n_471), .B(n_467), .Y(n_476) );
endmodule