module fake_jpeg_3773_n_328 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_19;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_30),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_16),
.B1(n_14),
.B2(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_18),
.B(n_6),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_13),
.CON(n_41),
.SN(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_13),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_31),
.A2(n_14),
.B1(n_26),
.B2(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_46),
.B1(n_31),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_48),
.B(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_33),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_52),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_44),
.B1(n_54),
.B2(n_47),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_68),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_30),
.C(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_73),
.B1(n_54),
.B2(n_44),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_72),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_45),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_38),
.C(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_75),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_38),
.C(n_12),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_40),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_82),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_83),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_0),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_40),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_86),
.Y(n_106)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_91),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_61),
.B1(n_90),
.B2(n_76),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_54),
.B1(n_44),
.B2(n_39),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_78),
.B1(n_52),
.B2(n_64),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_59),
.B(n_0),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_98),
.B(n_99),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_40),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_65),
.Y(n_122)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_57),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_94),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_87),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_89),
.B1(n_66),
.B2(n_92),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_110),
.B1(n_97),
.B2(n_101),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_SL g109 ( 
.A(n_87),
.Y(n_109)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_109),
.Y(n_145)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_114),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_80),
.A2(n_70),
.B1(n_57),
.B2(n_73),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_119),
.B1(n_124),
.B2(n_88),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_86),
.B(n_43),
.Y(n_147)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_83),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_73),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_100),
.CI(n_96),
.CON(n_130),
.SN(n_130)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_70),
.B1(n_32),
.B2(n_51),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_83),
.B(n_29),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_121),
.A2(n_83),
.B(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_122),
.B(n_94),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_78),
.B1(n_32),
.B2(n_53),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_98),
.B(n_99),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_129),
.B(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_79),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_127),
.B(n_128),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_123),
.B(n_112),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_136),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_135),
.B(n_102),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_95),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_139),
.B1(n_141),
.B2(n_107),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_138),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_108),
.B1(n_117),
.B2(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_140),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_110),
.B1(n_104),
.B2(n_97),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_143),
.A2(n_147),
.B1(n_150),
.B2(n_64),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_106),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_144),
.B(n_64),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_105),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_127),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_100),
.B(n_84),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_148),
.A2(n_149),
.B(n_104),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_118),
.A2(n_100),
.B(n_84),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_SL g150 ( 
.A1(n_118),
.A2(n_29),
.B(n_49),
.C(n_2),
.Y(n_150)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_148),
.CI(n_132),
.CON(n_183),
.SN(n_183)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_122),
.B(n_115),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_158),
.B(n_14),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_149),
.A2(n_115),
.B(n_102),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_164),
.B(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_161),
.Y(n_179)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_167),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_124),
.Y(n_164)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_34),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_168),
.B(n_148),
.C(n_125),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_137),
.A2(n_103),
.B1(n_78),
.B2(n_111),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_169),
.A2(n_172),
.B1(n_178),
.B2(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_171),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_111),
.B1(n_32),
.B2(n_77),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_132),
.B1(n_144),
.B2(n_138),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_26),
.Y(n_174)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_136),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_77),
.B1(n_29),
.B2(n_114),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_169),
.A2(n_147),
.B1(n_143),
.B2(n_128),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_196),
.B1(n_199),
.B2(n_204),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_182),
.A2(n_201),
.B1(n_205),
.B2(n_164),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_200),
.C(n_152),
.Y(n_212)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_151),
.A2(n_125),
.B(n_150),
.C(n_145),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_193),
.B(n_197),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_192),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

OAI31xp33_ASAP7_75t_L g193 ( 
.A1(n_151),
.A2(n_146),
.A3(n_130),
.B(n_150),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_163),
.B1(n_157),
.B2(n_170),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_150),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_172),
.A2(n_150),
.B1(n_130),
.B2(n_77),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_55),
.C(n_34),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_154),
.A2(n_8),
.B(n_12),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_202),
.B(n_161),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_159),
.A2(n_142),
.B1(n_145),
.B2(n_29),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_156),
.A2(n_145),
.B1(n_20),
.B2(n_34),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_207),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_152),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_208),
.B(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_153),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_211),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_213),
.C(n_214),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_179),
.B(n_174),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_200),
.B(n_158),
.C(n_153),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_215),
.C(n_224),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_175),
.C(n_160),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_218),
.B(n_223),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_220),
.A2(n_222),
.B1(n_227),
.B2(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_186),
.B1(n_195),
.B2(n_183),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_167),
.B1(n_171),
.B2(n_157),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_162),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_165),
.C(n_68),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_34),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_68),
.C(n_55),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_205),
.C(n_203),
.Y(n_236)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_226),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_232),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_231),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_180),
.C(n_187),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_199),
.B1(n_194),
.B2(n_190),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_234),
.A2(n_217),
.B1(n_209),
.B2(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_190),
.C(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_227),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_242),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_201),
.C(n_186),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_186),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_248),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_162),
.C(n_68),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_246),
.B(n_247),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_68),
.C(n_55),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_225),
.B(n_55),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_145),
.C(n_74),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_250),
.A2(n_255),
.B1(n_266),
.B2(n_246),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_236),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_253),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_249),
.A2(n_210),
.B1(n_74),
.B2(n_71),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_244),
.B(n_210),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_7),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

AO221x1_ASAP7_75t_L g276 ( 
.A1(n_263),
.A2(n_9),
.B1(n_12),
.B2(n_3),
.C(n_4),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_10),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_265),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_74),
.B1(n_71),
.B2(n_24),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_235),
.B(n_9),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_267),
.B(n_10),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_235),
.C(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_275),
.C(n_283),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g269 ( 
.A(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_7),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_240),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_278),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_282),
.B(n_280),
.Y(n_290)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_273),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_8),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_248),
.C(n_71),
.Y(n_275)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_276),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_260),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_260),
.A2(n_8),
.B1(n_12),
.B2(n_3),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_254),
.A2(n_19),
.B1(n_17),
.B2(n_1),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_266),
.B1(n_265),
.B2(n_261),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_1),
.C(n_2),
.Y(n_283)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_270),
.A2(n_275),
.B1(n_279),
.B2(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_6),
.C(n_10),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_292),
.A2(n_293),
.B(n_7),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_281),
.B(n_256),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g300 ( 
.A(n_294),
.B(n_269),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_283),
.C(n_278),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_271),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_302),
.C(n_304),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_268),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_300),
.B(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_285),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_259),
.C(n_282),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_8),
.C(n_10),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_4),
.B(n_5),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_301),
.A2(n_284),
.B1(n_289),
.B2(n_287),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_315),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_314),
.B(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_313),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_296),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_305),
.B(n_5),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_315),
.C(n_5),
.Y(n_321)
);

NAND2xp33_ASAP7_75t_L g319 ( 
.A(n_312),
.B(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_319),
.B(n_308),
.Y(n_320)
);

AO21x1_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_321),
.B(n_316),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_322),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_323),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_317),
.C(n_5),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_1),
.C(n_2),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_9),
.Y(n_327)
);

AO21x1_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_11),
.B(n_300),
.Y(n_328)
);


endmodule