module fake_jpeg_22694_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_47),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_42),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_49),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_7),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_39),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_54),
.B1(n_62),
.B2(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_37),
.B1(n_24),
.B2(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_60),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_35),
.B1(n_36),
.B2(n_32),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_48),
.A2(n_37),
.B1(n_24),
.B2(n_34),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_39),
.A2(n_37),
.B1(n_38),
.B2(n_34),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_44),
.A2(n_38),
.B1(n_20),
.B2(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_45),
.A2(n_20),
.B1(n_29),
.B2(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_61),
.A2(n_67),
.B1(n_70),
.B2(n_75),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_27),
.B1(n_33),
.B2(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_71),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_66),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_27),
.B1(n_22),
.B2(n_29),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_28),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_28),
.B1(n_18),
.B2(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_0),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_18),
.B1(n_35),
.B2(n_36),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_35),
.C(n_36),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_87),
.Y(n_99)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_35),
.B1(n_26),
.B2(n_23),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_26),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_76),
.B(n_89),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_51),
.A2(n_26),
.B1(n_23),
.B2(n_5),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_82),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_39),
.A2(n_23),
.B1(n_4),
.B2(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_90),
.B1(n_7),
.B2(n_8),
.Y(n_102)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_1),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_39),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_6),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_10),
.Y(n_112)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_95),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_66),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_17),
.B(n_8),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_91),
.B(n_86),
.C(n_81),
.Y(n_126)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_108),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_102),
.A2(n_111),
.B1(n_54),
.B2(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_8),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_89),
.B(n_58),
.Y(n_137)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_109),
.A2(n_59),
.B1(n_74),
.B2(n_73),
.Y(n_141)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_112),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_58),
.B(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_93),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_90),
.A2(n_78),
.B1(n_71),
.B2(n_54),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_54),
.B1(n_69),
.B2(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_126),
.B(n_129),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_76),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_128),
.B(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_69),
.B1(n_82),
.B2(n_80),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_119),
.B1(n_113),
.B2(n_94),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_115),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_139),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_107),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_148),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_147),
.Y(n_157)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_59),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_57),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_96),
.A2(n_57),
.B1(n_88),
.B2(n_73),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_64),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_118),
.B(n_72),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_102),
.A2(n_63),
.B1(n_77),
.B2(n_14),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_156),
.A2(n_117),
.B1(n_120),
.B2(n_129),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_160),
.A2(n_164),
.B1(n_169),
.B2(n_184),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_174),
.B1(n_145),
.B2(n_143),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_162),
.B(n_175),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_101),
.B1(n_114),
.B2(n_121),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_132),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_170),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_138),
.A2(n_122),
.B1(n_101),
.B2(n_114),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_107),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_173),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_146),
.A2(n_140),
.B1(n_144),
.B2(n_131),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_125),
.Y(n_175)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_181),
.Y(n_196)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_153),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_113),
.B(n_100),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_185),
.B1(n_137),
.B2(n_150),
.Y(n_193)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_144),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_130),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_125),
.B1(n_124),
.B2(n_121),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_124),
.B(n_77),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_128),
.Y(n_190)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_146),
.B1(n_147),
.B2(n_128),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_171),
.A2(n_134),
.B1(n_150),
.B2(n_135),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_186),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_104),
.B1(n_130),
.B2(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_108),
.Y(n_203)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_167),
.B(n_136),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_206),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_104),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

OAI21x1_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_104),
.B(n_158),
.Y(n_218)
);

FAx1_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_179),
.CI(n_173),
.CON(n_216),
.SN(n_216)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_216),
.A2(n_225),
.B1(n_176),
.B2(n_207),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g217 ( 
.A1(n_205),
.A2(n_166),
.B(n_183),
.Y(n_217)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_218),
.A2(n_180),
.B1(n_178),
.B2(n_196),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_162),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_227),
.C(n_229),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_206),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_208),
.A2(n_185),
.B1(n_179),
.B2(n_177),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_179),
.C(n_166),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_169),
.C(n_160),
.Y(n_229)
);

AOI322xp5_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_198),
.A3(n_187),
.B1(n_188),
.B2(n_203),
.C1(n_202),
.C2(n_197),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_212),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_187),
.B1(n_209),
.B2(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_189),
.C(n_199),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_235),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_228),
.A2(n_163),
.B1(n_204),
.B2(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_237),
.Y(n_253)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_240),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_226),
.A2(n_163),
.B1(n_177),
.B2(n_195),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_239),
.Y(n_246)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_196),
.C(n_200),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_217),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_149),
.C(n_126),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_126),
.C(n_13),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_225),
.Y(n_256)
);

FAx1_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_224),
.CI(n_216),
.CON(n_247),
.SN(n_247)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_247),
.B(n_212),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_219),
.Y(n_261)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_224),
.B(n_222),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_222),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_231),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_232),
.Y(n_260)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_215),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_262),
.A2(n_263),
.B(n_265),
.Y(n_267)
);

BUFx24_ASAP7_75t_SL g263 ( 
.A(n_256),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_246),
.B1(n_245),
.B2(n_250),
.Y(n_270)
);

AOI21xp33_ASAP7_75t_L g265 ( 
.A1(n_252),
.A2(n_213),
.B(n_219),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_231),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_249),
.C(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_233),
.C(n_249),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_273),
.C(n_241),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_213),
.B1(n_248),
.B2(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_268),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_269),
.A2(n_255),
.B(n_220),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_215),
.B(n_220),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_251),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_278),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_272),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_280),
.C(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_273),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_283),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_284),
.A2(n_285),
.B(n_243),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_267),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_287),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_286),
.Y(n_289)
);


endmodule