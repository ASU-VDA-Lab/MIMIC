module fake_aes_9629_n_28 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_3), .B(n_12), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_1), .B(n_5), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_20) );
CKINVDCx20_ASAP7_75t_R g21 ( .A(n_19), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
NOR2x1_ASAP7_75t_L g23 ( .A(n_22), .B(n_17), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .C(n_20), .Y(n_24) );
INVx1_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
OAI22x1_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_17), .B1(n_16), .B2(n_3), .Y(n_26) );
AOI31xp33_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_18), .A3(n_2), .B(n_4), .Y(n_27) );
AOI322xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_0), .A3(n_4), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_13), .Y(n_28) );
endmodule