module fake_jpeg_6937_n_46 (n_3, n_2, n_1, n_0, n_4, n_5, n_46);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_46;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_2),
.Y(n_7)
);

BUFx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_16),
.B(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NAND2x1_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_10),
.B(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_2),
.C(n_5),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_22),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_19),
.C(n_15),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_19),
.C(n_25),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_30),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_36),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_28),
.C(n_20),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_17),
.B1(n_28),
.B2(n_26),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_34),
.B(n_6),
.C(n_12),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_40),
.B(n_42),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_33),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_35),
.B(n_12),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_44),
.A2(n_13),
.B(n_5),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_45),
.A2(n_13),
.B(n_43),
.Y(n_46)
);


endmodule