module fake_netlist_6_2209_n_1779 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1779);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1779;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_125),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_31),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_18),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_70),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_105),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_36),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_41),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_101),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_54),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_26),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_77),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_36),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_8),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_26),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_27),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_28),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_49),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_89),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_18),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_7),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_59),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_67),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_4),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_62),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_40),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_14),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_56),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_122),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_65),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_74),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_9),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_87),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_142),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_76),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_115),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_47),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_37),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_30),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_146),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_78),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_15),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_32),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_5),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_7),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_68),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_81),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_154),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_13),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_104),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_3),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_128),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_111),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_57),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_12),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_134),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_103),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_45),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_91),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_50),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_151),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_56),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_43),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_31),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_84),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_20),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_37),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_34),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_32),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_54),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_16),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_17),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_94),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_92),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_132),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_108),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_88),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_25),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_49),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_96),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_61),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_141),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_20),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_130),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_121),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_27),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_35),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_79),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_110),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_97),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_72),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_51),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_38),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_19),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_119),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_11),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_35),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_23),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_127),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_45),
.Y(n_291)
);

BUFx8_ASAP7_75t_SL g292 ( 
.A(n_90),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_24),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_52),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_16),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_66),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_73),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_51),
.Y(n_299)
);

BUFx2_ASAP7_75t_SL g300 ( 
.A(n_10),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_38),
.Y(n_301)
);

BUFx4f_ASAP7_75t_SL g302 ( 
.A(n_47),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_100),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_10),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_17),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_242),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_219),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_242),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_292),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_155),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_219),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_242),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_242),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_294),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_204),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_295),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_161),
.B(n_0),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_274),
.B(n_0),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_295),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_304),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_257),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_271),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_165),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_304),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_274),
.B(n_2),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_167),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_168),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_187),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_2),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_282),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_187),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_282),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_159),
.B(n_3),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_170),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_174),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_271),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_271),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_176),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_177),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_180),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_291),
.Y(n_364)
);

BUFx10_ASAP7_75t_L g365 ( 
.A(n_258),
.Y(n_365)
);

INVxp33_ASAP7_75t_L g366 ( 
.A(n_156),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_291),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_156),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_169),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_169),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_184),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_173),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_158),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_187),
.B(n_4),
.Y(n_375)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_173),
.B(n_5),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_211),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_188),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_196),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_199),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_178),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_200),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_309),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_309),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_158),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_374),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_374),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

OA21x2_ASAP7_75t_L g390 ( 
.A1(n_311),
.A2(n_317),
.B(n_316),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_337),
.B(n_158),
.Y(n_393)
);

OA21x2_ASAP7_75t_L g394 ( 
.A1(n_317),
.A2(n_186),
.B(n_182),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_321),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_337),
.B(n_351),
.Y(n_398)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_194),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_322),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_L g403 ( 
.A(n_341),
.B(n_258),
.Y(n_403)
);

OAI21x1_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_259),
.B(n_194),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_322),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_333),
.B(n_216),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_324),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_347),
.Y(n_409)
);

CKINVDCx6p67_ASAP7_75t_R g410 ( 
.A(n_342),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_308),
.Y(n_411)
);

BUFx8_ASAP7_75t_L g412 ( 
.A(n_315),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

NOR2x1_ASAP7_75t_L g414 ( 
.A(n_325),
.B(n_194),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_326),
.B(n_259),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_326),
.B(n_259),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_310),
.A2(n_172),
.B1(n_191),
.B2(n_217),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_327),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_365),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_327),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_290),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_328),
.B(n_290),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_328),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_356),
.B(n_290),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_331),
.B(n_159),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_331),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_334),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_334),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_335),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_335),
.B(n_164),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_365),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_354),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_339),
.B(n_164),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_339),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_332),
.B(n_171),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_356),
.B(n_189),
.Y(n_440)
);

AND2x4_ASAP7_75t_L g441 ( 
.A(n_346),
.B(n_189),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_340),
.B(n_192),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_343),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_343),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_349),
.B(n_192),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_349),
.Y(n_447)
);

OA21x2_ASAP7_75t_L g448 ( 
.A1(n_350),
.A2(n_186),
.B(n_182),
.Y(n_448)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_350),
.A2(n_203),
.B(n_197),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_352),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_406),
.A2(n_314),
.B1(n_353),
.B2(n_346),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_411),
.B(n_378),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_439),
.B1(n_441),
.B2(n_403),
.Y(n_455)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_390),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_411),
.B(n_378),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_424),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_424),
.B(n_345),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_388),
.Y(n_461)
);

OAI22xp33_ASAP7_75t_L g462 ( 
.A1(n_439),
.A2(n_376),
.B1(n_366),
.B2(n_234),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_430),
.B(n_313),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_398),
.B(n_318),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_440),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_390),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g471 ( 
.A(n_409),
.B(n_430),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_436),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_427),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_388),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_448),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_387),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_448),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_357),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_430),
.B(n_320),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_398),
.B(n_193),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_441),
.A2(n_376),
.B1(n_203),
.B2(n_212),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_448),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_387),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_440),
.B(n_358),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_387),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_427),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_384),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_384),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_422),
.B(n_193),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_450),
.B(n_323),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_449),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_404),
.B(n_207),
.Y(n_501)
);

AND2x6_ASAP7_75t_L g502 ( 
.A(n_427),
.B(n_258),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_385),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_420),
.B(n_338),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_409),
.A2(n_379),
.B1(n_355),
.B2(n_360),
.Y(n_505)
);

INVx5_ASAP7_75t_L g506 ( 
.A(n_427),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_449),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_399),
.B(n_344),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

INVx4_ASAP7_75t_L g510 ( 
.A(n_427),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_387),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_449),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_420),
.B(n_361),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_392),
.Y(n_514)
);

BUFx8_ASAP7_75t_SL g515 ( 
.A(n_436),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_SL g516 ( 
.A(n_399),
.B(n_312),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_420),
.B(n_362),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_449),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_385),
.Y(n_520)
);

OR2x6_ASAP7_75t_L g521 ( 
.A(n_422),
.B(n_441),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_389),
.Y(n_522)
);

HAxp5_ASAP7_75t_SL g523 ( 
.A(n_418),
.B(n_197),
.CON(n_523),
.SN(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_420),
.B(n_372),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_449),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

OAI22xp33_ASAP7_75t_L g527 ( 
.A1(n_418),
.A2(n_252),
.B1(n_220),
.B2(n_221),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_399),
.B(n_380),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_449),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_410),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_449),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_441),
.A2(n_260),
.B1(n_251),
.B2(n_249),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_440),
.B(n_358),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_394),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_392),
.Y(n_537)
);

OAI22xp33_ASAP7_75t_L g538 ( 
.A1(n_418),
.A2(n_179),
.B1(n_239),
.B2(n_213),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

AND2x2_ASAP7_75t_SL g540 ( 
.A(n_403),
.B(n_258),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_420),
.B(n_381),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_427),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_394),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_396),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_450),
.B(n_383),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_441),
.A2(n_260),
.B1(n_212),
.B2(n_237),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_396),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_394),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_420),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_396),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_394),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_399),
.B(n_201),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_441),
.A2(n_275),
.B1(n_254),
.B2(n_285),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_440),
.B(n_359),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_397),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_410),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_435),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_422),
.B(n_207),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_394),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_399),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_394),
.Y(n_564)
);

OR2x6_ASAP7_75t_L g565 ( 
.A(n_422),
.B(n_300),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_397),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_397),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_416),
.B(n_359),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_399),
.B(n_202),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_410),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_441),
.A2(n_248),
.B1(n_230),
.B2(n_268),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_422),
.A2(n_393),
.B1(n_426),
.B2(n_404),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_399),
.B(n_412),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_422),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_435),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_392),
.Y(n_577)
);

NAND3xp33_ASAP7_75t_L g578 ( 
.A(n_393),
.B(n_364),
.C(n_363),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g579 ( 
.A(n_410),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_393),
.B(n_363),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_435),
.B(n_261),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_422),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_435),
.B(n_393),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_L g584 ( 
.A(n_426),
.B(n_258),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_392),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_416),
.B(n_364),
.Y(n_586)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_426),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_392),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_426),
.A2(n_301),
.B1(n_285),
.B2(n_288),
.Y(n_589)
);

INVx8_ASAP7_75t_L g590 ( 
.A(n_435),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_428),
.B(n_367),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_402),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_416),
.B(n_367),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_416),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_414),
.B(n_258),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_395),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_402),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_445),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_416),
.B(n_270),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_416),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_412),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_459),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_467),
.B(n_416),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_515),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_471),
.B(n_368),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_458),
.B(n_412),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_467),
.B(n_438),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_547),
.Y(n_609)
);

INVx2_ASAP7_75t_SL g610 ( 
.A(n_459),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_455),
.B(n_438),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_537),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_438),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_591),
.B(n_438),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_466),
.B(n_412),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_521),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_499),
.B(n_412),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_547),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_548),
.B(n_412),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_590),
.A2(n_386),
.B(n_401),
.Y(n_620)
);

NAND2x1_ASAP7_75t_L g621 ( 
.A(n_552),
.B(n_438),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_438),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_481),
.B(n_402),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_481),
.B(n_405),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_575),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_537),
.Y(n_627)
);

INVx1_ASAP7_75t_SL g628 ( 
.A(n_454),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_476),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_483),
.A2(n_329),
.B1(n_336),
.B2(n_412),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_568),
.B(n_405),
.Y(n_631)
);

NOR3xp33_ASAP7_75t_L g632 ( 
.A(n_505),
.B(n_297),
.C(n_166),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_586),
.B(n_405),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_495),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_593),
.B(n_408),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_581),
.B(n_408),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_483),
.A2(n_208),
.B1(n_206),
.B2(n_205),
.Y(n_637)
);

NOR3xp33_ASAP7_75t_L g638 ( 
.A(n_527),
.B(n_175),
.C(n_157),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_465),
.B(n_302),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_454),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_563),
.B(n_404),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_580),
.B(n_408),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_L g643 ( 
.A(n_494),
.B(n_428),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_575),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_473),
.Y(n_645)
);

O2A1O1Ixp33_ASAP7_75t_L g646 ( 
.A1(n_478),
.A2(n_401),
.B(n_428),
.C(n_446),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

AOI22xp5_ASAP7_75t_L g648 ( 
.A1(n_483),
.A2(n_243),
.B1(n_214),
.B2(n_215),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_540),
.B(n_419),
.Y(n_649)
);

AOI22xp5_ASAP7_75t_L g650 ( 
.A1(n_483),
.A2(n_280),
.B1(n_225),
.B2(n_226),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_582),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_457),
.B(n_369),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_478),
.A2(n_404),
.B1(n_288),
.B2(n_307),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_540),
.B(n_419),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_540),
.B(n_421),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_547),
.B(n_209),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_521),
.Y(n_657)
);

O2A1O1Ixp33_ASAP7_75t_L g658 ( 
.A1(n_480),
.A2(n_401),
.B(n_434),
.C(n_446),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_489),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_583),
.B(n_421),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_489),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_457),
.B(n_237),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_535),
.B(n_421),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_473),
.B(n_228),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_535),
.B(n_425),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_547),
.B(n_229),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_473),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_557),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_557),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_482),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_537),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_547),
.B(n_231),
.Y(n_673)
);

NOR3xp33_ASAP7_75t_L g674 ( 
.A(n_538),
.B(n_183),
.C(n_181),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_456),
.B(n_425),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_473),
.B(n_232),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_480),
.A2(n_301),
.B(n_303),
.C(n_249),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_456),
.B(n_425),
.Y(n_679)
);

INVxp33_ASAP7_75t_L g680 ( 
.A(n_571),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_462),
.B(n_190),
.Y(n_681)
);

BUFx6f_ASAP7_75t_SL g682 ( 
.A(n_497),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_456),
.B(n_195),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_495),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_453),
.B(n_185),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_477),
.B(n_429),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_185),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_496),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_531),
.B(n_185),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_473),
.B(n_236),
.Y(n_690)
);

OR2x2_ASAP7_75t_SL g691 ( 
.A(n_523),
.B(n_245),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_497),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_477),
.B(n_429),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_559),
.B(n_185),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_477),
.B(n_504),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_L g696 ( 
.A(n_578),
.B(n_599),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_592),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_496),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_513),
.B(n_429),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_517),
.B(n_431),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_564),
.B(n_240),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_524),
.B(n_431),
.Y(n_703)
);

HB1xp67_ASAP7_75t_L g704 ( 
.A(n_565),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_597),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_564),
.B(n_247),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_541),
.B(n_431),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_460),
.B(n_433),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_579),
.B(n_369),
.Y(n_710)
);

INVx3_ASAP7_75t_L g711 ( 
.A(n_521),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_503),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_460),
.B(n_433),
.Y(n_713)
);

NOR3xp33_ASAP7_75t_L g714 ( 
.A(n_472),
.B(n_246),
.C(n_244),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_521),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_503),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_486),
.B(n_370),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_564),
.B(n_256),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_564),
.B(n_266),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_564),
.B(n_267),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_463),
.B(n_433),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_552),
.B(n_269),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_519),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_484),
.A2(n_434),
.B(n_446),
.C(n_442),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_528),
.Y(n_725)
);

O2A1O1Ixp5_ASAP7_75t_L g726 ( 
.A1(n_484),
.A2(n_386),
.B(n_434),
.C(n_437),
.Y(n_726)
);

BUFx3_ASAP7_75t_L g727 ( 
.A(n_497),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_552),
.B(n_273),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_552),
.B(n_277),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_523),
.B(n_578),
.C(n_589),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_574),
.B(n_279),
.Y(n_731)
);

BUFx6f_ASAP7_75t_SL g732 ( 
.A(n_497),
.Y(n_732)
);

INVxp67_ASAP7_75t_SL g733 ( 
.A(n_493),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_596),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_519),
.Y(n_735)
);

A2O1A1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_487),
.A2(n_307),
.B(n_245),
.C(n_275),
.Y(n_736)
);

AOI22xp5_ASAP7_75t_L g737 ( 
.A1(n_565),
.A2(n_284),
.B1(n_286),
.B2(n_293),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_463),
.B(n_464),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_574),
.B(n_493),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_464),
.B(n_210),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_572),
.A2(n_210),
.B1(n_278),
.B2(n_238),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_470),
.B(n_218),
.Y(n_742)
);

NAND3xp33_ASAP7_75t_SL g743 ( 
.A(n_516),
.B(n_198),
.C(n_222),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_561),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_470),
.B(n_218),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_475),
.B(n_227),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_475),
.B(n_223),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_487),
.B(n_233),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_561),
.B(n_370),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_574),
.B(n_223),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_491),
.B(n_492),
.Y(n_751)
);

NAND3xp33_ASAP7_75t_L g752 ( 
.A(n_533),
.B(n_281),
.C(n_235),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_574),
.B(n_224),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_493),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_563),
.B(n_296),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_491),
.B(n_224),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_520),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_508),
.B(n_264),
.C(n_241),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_596),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_493),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_492),
.B(n_238),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_493),
.B(n_305),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_596),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_520),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_529),
.B(n_437),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_498),
.A2(n_437),
.B(n_442),
.C(n_386),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_534),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_498),
.B(n_250),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_479),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_500),
.B(n_272),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_534),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_615),
.A2(n_565),
.B1(n_561),
.B2(n_569),
.Y(n_772)
);

INVx2_ASAP7_75t_SL g773 ( 
.A(n_710),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_671),
.B(n_507),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_680),
.B(n_507),
.Y(n_775)
);

A2O1A1Ixp33_ASAP7_75t_L g776 ( 
.A1(n_617),
.A2(n_532),
.B(n_512),
.C(n_530),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_643),
.B(n_512),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_611),
.A2(n_525),
.B(n_518),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_738),
.B(n_518),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_620),
.A2(n_590),
.B(n_539),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_739),
.A2(n_590),
.B(n_539),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_603),
.B(n_525),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_628),
.B(n_570),
.Y(n_783)
);

O2A1O1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_741),
.A2(n_562),
.B(n_544),
.C(n_536),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_739),
.A2(n_590),
.B(n_539),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_645),
.A2(n_590),
.B(n_539),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_743),
.B(n_573),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_615),
.A2(n_565),
.B1(n_561),
.B2(n_555),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_695),
.A2(n_532),
.B(n_530),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_609),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_738),
.B(n_536),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_751),
.B(n_544),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_602),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_751),
.B(n_551),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_617),
.A2(n_601),
.B1(n_600),
.B2(n_594),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_626),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_699),
.B(n_551),
.Y(n_797)
);

O2A1O1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_677),
.A2(n_554),
.B(n_562),
.C(n_584),
.Y(n_798)
);

OAI21xp33_ASAP7_75t_L g799 ( 
.A1(n_681),
.A2(n_556),
.B(n_549),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_645),
.A2(n_510),
.B(n_546),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_675),
.A2(n_554),
.B(n_501),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_668),
.A2(n_510),
.B(n_546),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_602),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_701),
.B(n_594),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_730),
.A2(n_501),
.B1(n_601),
.B2(n_251),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_668),
.A2(n_510),
.B(n_546),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_679),
.A2(n_501),
.B(n_600),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_767),
.A2(n_510),
.B(n_546),
.Y(n_808)
);

OAI22xp5_ASAP7_75t_L g809 ( 
.A1(n_619),
.A2(n_600),
.B1(n_594),
.B2(n_560),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_644),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_703),
.B(n_594),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_619),
.A2(n_298),
.B(n_278),
.C(n_560),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_708),
.B(n_600),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_613),
.B(n_560),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_609),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_610),
.B(n_296),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_767),
.A2(n_542),
.B(n_534),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_616),
.B(n_371),
.Y(n_818)
);

AO21x1_ASAP7_75t_L g819 ( 
.A1(n_656),
.A2(n_298),
.B(n_526),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_629),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_771),
.A2(n_534),
.B(n_542),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_647),
.Y(n_822)
);

NOR2x1_ASAP7_75t_R g823 ( 
.A(n_605),
.B(n_253),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_683),
.B(n_522),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_651),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_689),
.B(n_694),
.Y(n_826)
);

O2A1O1Ixp5_ASAP7_75t_L g827 ( 
.A1(n_631),
.A2(n_522),
.B(n_545),
.C(n_526),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_616),
.B(n_371),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_683),
.B(n_543),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_685),
.A2(n_303),
.B1(n_254),
.B2(n_595),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_771),
.A2(n_542),
.B(n_534),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_765),
.A2(n_595),
.B1(n_488),
.B2(n_490),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_606),
.Y(n_833)
);

BUFx2_ASAP7_75t_SL g834 ( 
.A(n_682),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_609),
.B(n_542),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_609),
.Y(n_836)
);

BUFx2_ASAP7_75t_L g837 ( 
.A(n_640),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_746),
.B(n_543),
.Y(n_838)
);

AOI22xp5_ASAP7_75t_L g839 ( 
.A1(n_696),
.A2(n_595),
.B1(n_490),
.B2(n_479),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_639),
.B(n_296),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_659),
.A2(n_669),
.B1(n_670),
.B2(n_662),
.Y(n_841)
);

OAI21x1_ASAP7_75t_L g842 ( 
.A1(n_621),
.A2(n_567),
.B(n_545),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_652),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_618),
.B(n_542),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_618),
.A2(n_528),
.B(n_506),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_746),
.B(n_550),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_678),
.B(n_550),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_697),
.Y(n_848)
);

CKINVDCx10_ASAP7_75t_R g849 ( 
.A(n_663),
.Y(n_849)
);

NOR2xp67_ASAP7_75t_L g850 ( 
.A(n_737),
.B(n_479),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_618),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_618),
.A2(n_528),
.B(n_506),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_733),
.A2(n_506),
.B(n_576),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_700),
.B(n_706),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_636),
.B(n_553),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_L g856 ( 
.A1(n_649),
.A2(n_576),
.B1(n_553),
.B2(n_558),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_SL g857 ( 
.A1(n_691),
.A2(n_265),
.B1(n_262),
.B2(n_276),
.Y(n_857)
);

NOR2x2_ASAP7_75t_L g858 ( 
.A(n_663),
.B(n_681),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_604),
.A2(n_506),
.B(n_576),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_686),
.A2(n_558),
.B(n_566),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_642),
.B(n_566),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_607),
.B(n_296),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_748),
.B(n_479),
.Y(n_863)
);

BUFx12f_ASAP7_75t_L g864 ( 
.A(n_663),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_748),
.B(n_485),
.Y(n_865)
);

NAND2xp33_ASAP7_75t_SL g866 ( 
.A(n_755),
.B(n_255),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_768),
.B(n_485),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_693),
.A2(n_585),
.B(n_588),
.Y(n_868)
);

NOR3xp33_ASAP7_75t_L g869 ( 
.A(n_632),
.B(n_442),
.C(n_283),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_724),
.A2(n_377),
.B(n_382),
.C(n_373),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_687),
.Y(n_871)
);

AO21x1_ASAP7_75t_L g872 ( 
.A1(n_656),
.A2(n_423),
.B(n_417),
.Y(n_872)
);

AOI222xp33_ASAP7_75t_L g873 ( 
.A1(n_752),
.A2(n_299),
.B1(n_382),
.B2(n_377),
.C1(n_373),
.C2(n_417),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_727),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_754),
.A2(n_506),
.B(n_576),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_717),
.B(n_485),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_629),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_768),
.B(n_485),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_624),
.B(n_488),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_725),
.B(n_506),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_625),
.B(n_488),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_754),
.A2(n_576),
.B(n_509),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_622),
.B(n_657),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_614),
.B(n_488),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_622),
.B(n_490),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_754),
.A2(n_576),
.B(n_509),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_623),
.B(n_490),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_722),
.A2(n_729),
.B(n_728),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_664),
.B(n_596),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_657),
.B(n_509),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_634),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_749),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_666),
.B(n_461),
.Y(n_893)
);

NOR2x1_ASAP7_75t_L g894 ( 
.A(n_607),
.B(n_414),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_634),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_608),
.A2(n_414),
.B(n_511),
.C(n_415),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_749),
.B(n_461),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_754),
.A2(n_511),
.B(n_598),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_714),
.B(n_423),
.C(n_417),
.Y(n_899)
);

INVx11_ASAP7_75t_L g900 ( 
.A(n_682),
.Y(n_900)
);

NOR2x1p5_ASAP7_75t_L g901 ( 
.A(n_715),
.B(n_415),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_715),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_661),
.B(n_468),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_684),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_711),
.B(n_511),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_726),
.A2(n_588),
.B(n_585),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_677),
.A2(n_415),
.B(n_423),
.C(n_577),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_684),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_633),
.B(n_468),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_760),
.A2(n_598),
.B(n_469),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_727),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_688),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_760),
.A2(n_598),
.B(n_469),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_725),
.B(n_598),
.Y(n_914)
);

OAI321xp33_ASAP7_75t_L g915 ( 
.A1(n_736),
.A2(n_452),
.A3(n_451),
.B1(n_577),
.B2(n_514),
.C(n_407),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_635),
.B(n_474),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_769),
.B(n_654),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_760),
.A2(n_598),
.B(n_474),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_688),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_769),
.B(n_577),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_736),
.A2(n_514),
.B(n_395),
.C(n_451),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_711),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_760),
.A2(n_514),
.B(n_391),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_744),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_709),
.A2(n_391),
.B(n_400),
.Y(n_925)
);

AO21x1_ASAP7_75t_L g926 ( 
.A1(n_667),
.A2(n_395),
.B(n_451),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_766),
.A2(n_502),
.B(n_595),
.Y(n_927)
);

NAND2x1p5_ASAP7_75t_L g928 ( 
.A(n_744),
.B(n_391),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_698),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_655),
.B(n_502),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_713),
.A2(n_721),
.B(n_731),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_698),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_692),
.B(n_712),
.Y(n_933)
);

NAND2x1p5_ASAP7_75t_L g934 ( 
.A(n_716),
.B(n_391),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_722),
.A2(n_728),
.B(n_731),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_712),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_630),
.B(n_6),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_723),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_758),
.B(n_451),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_723),
.B(n_502),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_735),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_502),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_764),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_704),
.B(n_740),
.Y(n_944)
);

AOI22x1_ASAP7_75t_L g945 ( 
.A1(n_641),
.A2(n_395),
.B1(n_451),
.B2(n_452),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_612),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_704),
.B(n_6),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_742),
.B(n_9),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_729),
.A2(n_391),
.B(n_400),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_725),
.B(n_502),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_627),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_725),
.B(n_502),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_745),
.A2(n_395),
.B(n_452),
.C(n_432),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_747),
.A2(n_452),
.B(n_407),
.C(n_432),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_756),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_667),
.A2(n_391),
.B(n_400),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_725),
.B(n_502),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_725),
.B(n_595),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_646),
.A2(n_452),
.B(n_407),
.C(n_413),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_786),
.A2(n_673),
.B(n_719),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_804),
.A2(n_720),
.B1(n_702),
.B2(n_707),
.Y(n_961)
);

O2A1O1Ixp33_ASAP7_75t_L g962 ( 
.A1(n_937),
.A2(n_674),
.B(n_638),
.C(n_702),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_796),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_810),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_811),
.A2(n_720),
.B1(n_673),
.B2(n_707),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_955),
.B(n_775),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_822),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_837),
.Y(n_968)
);

BUFx8_ASAP7_75t_SL g969 ( 
.A(n_864),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_813),
.A2(n_719),
.B1(n_718),
.B2(n_641),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_825),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_793),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_902),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_848),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_775),
.B(n_761),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_843),
.Y(n_976)
);

OAI22xp5_ASAP7_75t_L g977 ( 
.A1(n_944),
.A2(n_718),
.B1(n_770),
.B2(n_753),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_871),
.B(n_637),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_790),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_790),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_877),
.Y(n_981)
);

O2A1O1Ixp5_ASAP7_75t_L g982 ( 
.A1(n_819),
.A2(n_762),
.B(n_750),
.C(n_759),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_876),
.B(n_653),
.Y(n_983)
);

INVx8_ASAP7_75t_L g984 ( 
.A(n_790),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_803),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_820),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_902),
.Y(n_987)
);

A2O1A1Ixp33_ASAP7_75t_SL g988 ( 
.A1(n_948),
.A2(n_774),
.B(n_869),
.C(n_944),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_876),
.B(n_653),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_800),
.A2(n_690),
.B(n_665),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_929),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_774),
.B(n_658),
.Y(n_992)
);

CKINVDCx11_ASAP7_75t_R g993 ( 
.A(n_902),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_790),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_891),
.Y(n_995)
);

AOI21x1_ASAP7_75t_L g996 ( 
.A1(n_824),
.A2(n_762),
.B(n_763),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_895),
.Y(n_997)
);

AOI21x1_ASAP7_75t_L g998 ( 
.A1(n_829),
.A2(n_734),
.B(n_660),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_773),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_833),
.B(n_650),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_841),
.B(n_799),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_866),
.B(n_705),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_841),
.B(n_705),
.Y(n_1003)
);

AOI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_937),
.A2(n_732),
.B1(n_595),
.B2(n_672),
.Y(n_1004)
);

BUFx2_ASAP7_75t_L g1005 ( 
.A(n_833),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_904),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_802),
.A2(n_676),
.B(n_648),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_SL g1008 ( 
.A(n_874),
.B(n_732),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_881),
.B(n_595),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_772),
.A2(n_432),
.B1(n_407),
.B2(n_444),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_908),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_806),
.A2(n_400),
.B(n_432),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_SL g1013 ( 
.A(n_818),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_948),
.A2(n_432),
.B(n_407),
.C(n_444),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_881),
.B(n_444),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_834),
.B(n_444),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_783),
.B(n_12),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_836),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_816),
.B(n_413),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_874),
.B(n_447),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_818),
.Y(n_1021)
);

O2A1O1Ixp5_ASAP7_75t_SL g1022 ( 
.A1(n_906),
.A2(n_400),
.B(n_14),
.C(n_15),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_R g1023 ( 
.A(n_862),
.B(n_63),
.Y(n_1023)
);

AND2x6_ASAP7_75t_L g1024 ( 
.A(n_787),
.B(n_444),
.Y(n_1024)
);

INVx3_ASAP7_75t_SL g1025 ( 
.A(n_858),
.Y(n_1025)
);

INVx1_ASAP7_75t_SL g1026 ( 
.A(n_849),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_912),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_869),
.A2(n_443),
.B1(n_413),
.B2(n_400),
.Y(n_1028)
);

CKINVDCx14_ASAP7_75t_R g1029 ( 
.A(n_857),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_919),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_R g1031 ( 
.A(n_902),
.B(n_60),
.Y(n_1031)
);

OR2x2_ASAP7_75t_L g1032 ( 
.A(n_828),
.B(n_443),
.Y(n_1032)
);

BUFx3_ASAP7_75t_L g1033 ( 
.A(n_828),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_808),
.A2(n_780),
.B(n_781),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_785),
.A2(n_443),
.B(n_413),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_947),
.A2(n_443),
.B(n_413),
.C(n_21),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_840),
.B(n_443),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_911),
.B(n_447),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_854),
.B(n_447),
.Y(n_1039)
);

HB1xp67_ASAP7_75t_L g1040 ( 
.A(n_836),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_788),
.A2(n_447),
.B1(n_445),
.B2(n_149),
.Y(n_1041)
);

AOI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_883),
.A2(n_447),
.B1(n_445),
.B2(n_148),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_797),
.A2(n_447),
.B1(n_445),
.B2(n_140),
.Y(n_1043)
);

OAI21xp33_ASAP7_75t_L g1044 ( 
.A1(n_830),
.A2(n_447),
.B(n_445),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_935),
.A2(n_447),
.B(n_445),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_932),
.Y(n_1046)
);

AOI33xp33_ASAP7_75t_L g1047 ( 
.A1(n_805),
.A2(n_13),
.A3(n_19),
.B1(n_22),
.B2(n_24),
.B3(n_28),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_931),
.A2(n_447),
.B(n_445),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_892),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_779),
.A2(n_445),
.B1(n_447),
.B2(n_139),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_947),
.B(n_22),
.Y(n_1051)
);

AO21x1_ASAP7_75t_L g1052 ( 
.A1(n_838),
.A2(n_29),
.B(n_30),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_936),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_911),
.B(n_445),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_807),
.A2(n_445),
.B(n_129),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_870),
.A2(n_29),
.B(n_33),
.C(n_34),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_836),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_817),
.A2(n_126),
.B(n_124),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_924),
.B(n_123),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_922),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_924),
.B(n_113),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_938),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_801),
.A2(n_33),
.B(n_39),
.C(n_41),
.Y(n_1063)
);

AND2x4_ASAP7_75t_L g1064 ( 
.A(n_883),
.B(n_99),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_836),
.B(n_93),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_842),
.A2(n_86),
.B(n_85),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_901),
.B(n_42),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_890),
.B(n_82),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_885),
.B(n_870),
.C(n_812),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_941),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_946),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_SL g1072 ( 
.A1(n_805),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_821),
.A2(n_75),
.B(n_71),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_873),
.B(n_44),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_782),
.B(n_46),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_830),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_943),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_850),
.A2(n_48),
.B(n_53),
.C(n_55),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_831),
.A2(n_69),
.B(n_55),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_SL g1080 ( 
.A1(n_795),
.A2(n_58),
.B1(n_939),
.B2(n_885),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_851),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_846),
.A2(n_878),
.B(n_865),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_851),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_899),
.A2(n_890),
.B1(n_939),
.B2(n_782),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_823),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_900),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_777),
.B(n_917),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_855),
.B(n_897),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_851),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_851),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_928),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_SL g1092 ( 
.A(n_815),
.B(n_791),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_928),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_927),
.A2(n_926),
.B(n_809),
.C(n_888),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_899),
.A2(n_915),
.B(n_905),
.C(n_860),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_933),
.B(n_792),
.Y(n_1096)
);

BUFx4f_ASAP7_75t_SL g1097 ( 
.A(n_815),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_794),
.B(n_861),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_951),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_879),
.B(n_814),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_776),
.A2(n_867),
.B1(n_863),
.B2(n_839),
.Y(n_1101)
);

AOI22xp5_ASAP7_75t_L g1102 ( 
.A1(n_894),
.A2(n_832),
.B1(n_872),
.B2(n_930),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_847),
.B(n_884),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_887),
.B(n_889),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_778),
.B(n_789),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_958),
.A2(n_950),
.B(n_957),
.Y(n_1106)
);

AO31x2_ASAP7_75t_L g1107 ( 
.A1(n_1082),
.A2(n_959),
.A3(n_896),
.B(n_856),
.Y(n_1107)
);

AOI221xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1074),
.A2(n_798),
.B1(n_907),
.B2(n_784),
.C(n_959),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_961),
.A2(n_956),
.A3(n_949),
.B(n_859),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1076),
.A2(n_1080),
.B(n_1051),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_976),
.B(n_903),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1034),
.A2(n_945),
.B(n_827),
.Y(n_1112)
);

OAI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1035),
.A2(n_827),
.B(n_868),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_978),
.B(n_893),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1048),
.A2(n_898),
.B(n_913),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_962),
.A2(n_925),
.B(n_916),
.C(n_909),
.Y(n_1116)
);

AO32x2_ASAP7_75t_L g1117 ( 
.A1(n_1072),
.A2(n_921),
.A3(n_954),
.B1(n_953),
.B2(n_914),
.Y(n_1117)
);

O2A1O1Ixp33_ASAP7_75t_L g1118 ( 
.A1(n_988),
.A2(n_914),
.B(n_844),
.C(n_835),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_965),
.A2(n_970),
.B(n_960),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1005),
.B(n_934),
.Y(n_1120)
);

AOI221xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1051),
.A2(n_1075),
.B1(n_1063),
.B2(n_1076),
.C(n_1001),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1098),
.B(n_920),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_990),
.A2(n_835),
.B(n_844),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1101),
.A2(n_942),
.B(n_940),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_966),
.B(n_934),
.Y(n_1125)
);

OAI21x1_ASAP7_75t_L g1126 ( 
.A1(n_1106),
.A2(n_918),
.B(n_910),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_983),
.A2(n_989),
.B(n_1088),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1055),
.A2(n_845),
.A3(n_852),
.B(n_923),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_963),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_964),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1098),
.B(n_882),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_979),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1017),
.A2(n_952),
.B1(n_880),
.B2(n_886),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_967),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_968),
.Y(n_1135)
);

AOI21x1_ASAP7_75t_L g1136 ( 
.A1(n_998),
.A2(n_880),
.B(n_853),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_971),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_SL g1138 ( 
.A1(n_977),
.A2(n_875),
.B(n_1104),
.Y(n_1138)
);

AOI221x1_ASAP7_75t_L g1139 ( 
.A1(n_1041),
.A2(n_1075),
.B1(n_992),
.B2(n_1050),
.C(n_1078),
.Y(n_1139)
);

OAI22x1_ASAP7_75t_L g1140 ( 
.A1(n_1017),
.A2(n_1025),
.B1(n_1084),
.B2(n_1064),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1086),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_999),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_979),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1007),
.A2(n_1105),
.B(n_1100),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_975),
.A2(n_1104),
.B(n_1103),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1103),
.A2(n_1095),
.B(n_1015),
.Y(n_1146)
);

BUFx10_ASAP7_75t_L g1147 ( 
.A(n_1013),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_974),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1045),
.A2(n_1012),
.B(n_996),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1070),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1066),
.A2(n_1094),
.B(n_982),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_988),
.A2(n_1102),
.B(n_1095),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1096),
.B(n_1087),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_999),
.Y(n_1154)
);

NAND2x1p5_ASAP7_75t_L g1155 ( 
.A(n_973),
.B(n_987),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1052),
.A2(n_1010),
.A3(n_1043),
.B(n_1014),
.Y(n_1156)
);

AO31x2_ASAP7_75t_L g1157 ( 
.A1(n_1087),
.A2(n_1009),
.A3(n_1079),
.B(n_1039),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1022),
.A2(n_1069),
.B(n_1037),
.Y(n_1158)
);

BUFx8_ASAP7_75t_L g1159 ( 
.A(n_1013),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_1003),
.A2(n_1058),
.A3(n_1073),
.B(n_1030),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_981),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1092),
.A2(n_1019),
.B(n_1020),
.Y(n_1162)
);

OR2x2_ASAP7_75t_L g1163 ( 
.A(n_1000),
.B(n_1032),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1033),
.B(n_1021),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1004),
.A2(n_1077),
.B1(n_973),
.B2(n_1064),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_995),
.A2(n_1053),
.A3(n_1011),
.B(n_1006),
.Y(n_1166)
);

NOR2xp67_ASAP7_75t_SL g1167 ( 
.A(n_1049),
.B(n_1085),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1020),
.A2(n_1054),
.B(n_1059),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_979),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1069),
.A2(n_1036),
.B(n_1056),
.C(n_1042),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1054),
.A2(n_1061),
.B(n_1059),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1061),
.A2(n_1044),
.B(n_1068),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_SL g1173 ( 
.A(n_1097),
.B(n_1025),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1046),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_972),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1068),
.A2(n_1038),
.B(n_1004),
.Y(n_1176)
);

INVx5_ASAP7_75t_L g1177 ( 
.A(n_984),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1067),
.B(n_1060),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_985),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_984),
.A2(n_1065),
.B(n_1062),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_1016),
.B(n_1093),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1099),
.B(n_1027),
.Y(n_1182)
);

CKINVDCx11_ASAP7_75t_R g1183 ( 
.A(n_1026),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_986),
.Y(n_1184)
);

OR2x6_ASAP7_75t_L g1185 ( 
.A(n_1016),
.B(n_1091),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_997),
.A2(n_991),
.A3(n_1071),
.B(n_1024),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_SL g1187 ( 
.A1(n_1018),
.A2(n_1090),
.B(n_1089),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1047),
.B(n_1008),
.Y(n_1188)
);

OAI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1028),
.A2(n_1024),
.B(n_1016),
.Y(n_1189)
);

INVx8_ASAP7_75t_L g1190 ( 
.A(n_980),
.Y(n_1190)
);

BUFx2_ASAP7_75t_L g1191 ( 
.A(n_1018),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1040),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1024),
.A2(n_1023),
.A3(n_1040),
.B(n_1089),
.Y(n_1193)
);

AOI22x1_ASAP7_75t_L g1194 ( 
.A1(n_1090),
.A2(n_1083),
.B1(n_1057),
.B2(n_1081),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_980),
.B(n_994),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1024),
.A2(n_1083),
.B(n_1081),
.Y(n_1196)
);

BUFx10_ASAP7_75t_L g1197 ( 
.A(n_1024),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1029),
.A2(n_1023),
.B1(n_1002),
.B2(n_1031),
.C(n_1057),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_1031),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_980),
.A2(n_994),
.B(n_1002),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_994),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_994),
.A2(n_1034),
.B(n_945),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_969),
.B(n_826),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_963),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1074),
.A2(n_412),
.B1(n_399),
.B2(n_937),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_988),
.A2(n_671),
.B(n_1051),
.C(n_439),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_1077),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_1086),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1101),
.A2(n_776),
.B(n_1102),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_961),
.A2(n_590),
.B(n_574),
.Y(n_1210)
);

INVxp67_ASAP7_75t_SL g1211 ( 
.A(n_999),
.Y(n_1211)
);

AO21x1_ASAP7_75t_L g1212 ( 
.A1(n_962),
.A2(n_1075),
.B(n_1041),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1034),
.A2(n_945),
.B(n_842),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_976),
.B(n_826),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_961),
.A2(n_590),
.B(n_574),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_963),
.Y(n_1216)
);

AOI221x1_ASAP7_75t_L g1217 ( 
.A1(n_1051),
.A2(n_1063),
.B1(n_961),
.B2(n_965),
.C(n_1041),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_993),
.Y(n_1218)
);

O2A1O1Ixp33_ASAP7_75t_SL g1219 ( 
.A1(n_988),
.A2(n_1063),
.B(n_1095),
.C(n_1001),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_976),
.B(n_871),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_993),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1034),
.A2(n_945),
.B(n_842),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_963),
.Y(n_1223)
);

A2O1A1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_962),
.A2(n_619),
.B(n_617),
.C(n_1075),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_988),
.A2(n_1063),
.B(n_1095),
.C(n_1001),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1074),
.A2(n_1051),
.B1(n_937),
.B2(n_1072),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1034),
.A2(n_945),
.B(n_842),
.Y(n_1227)
);

CKINVDCx8_ASAP7_75t_R g1228 ( 
.A(n_1086),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_1086),
.Y(n_1229)
);

AOI21x1_ASAP7_75t_L g1230 ( 
.A1(n_960),
.A2(n_888),
.B(n_935),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1082),
.A2(n_965),
.A3(n_961),
.B(n_970),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_961),
.A2(n_590),
.B(n_574),
.Y(n_1232)
);

AOI221x1_ASAP7_75t_L g1233 ( 
.A1(n_1051),
.A2(n_1063),
.B1(n_961),
.B2(n_965),
.C(n_1041),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_962),
.A2(n_619),
.B(n_617),
.C(n_1075),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_962),
.A2(n_619),
.B(n_617),
.C(n_1075),
.Y(n_1235)
);

CKINVDCx6p67_ASAP7_75t_R g1236 ( 
.A(n_993),
.Y(n_1236)
);

NOR4xp25_ASAP7_75t_L g1237 ( 
.A(n_1056),
.B(n_962),
.C(n_1074),
.D(n_1051),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_962),
.A2(n_619),
.B(n_617),
.C(n_1075),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_984),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_993),
.Y(n_1240)
);

CKINVDCx8_ASAP7_75t_R g1241 ( 
.A(n_1086),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_983),
.A2(n_619),
.B1(n_617),
.B2(n_671),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_963),
.Y(n_1243)
);

O2A1O1Ixp5_ASAP7_75t_L g1244 ( 
.A1(n_1082),
.A2(n_617),
.B(n_619),
.C(n_615),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_960),
.A2(n_888),
.B(n_935),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_963),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1226),
.A2(n_1110),
.B1(n_1212),
.B2(n_1205),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_SL g1248 ( 
.A1(n_1153),
.A2(n_1110),
.B1(n_1226),
.B2(n_1209),
.Y(n_1248)
);

BUFx8_ASAP7_75t_L g1249 ( 
.A(n_1218),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1224),
.A2(n_1234),
.B1(n_1235),
.B2(n_1238),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1159),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1183),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_1228),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1140),
.A2(n_1114),
.B1(n_1127),
.B2(n_1242),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1163),
.A2(n_1209),
.B1(n_1214),
.B2(n_1220),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1154),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1147),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1154),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1130),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1186),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1203),
.A2(n_1199),
.B1(n_1237),
.B2(n_1173),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1134),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1188),
.A2(n_1111),
.B1(n_1152),
.B2(n_1165),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1152),
.A2(n_1178),
.B1(n_1172),
.B2(n_1145),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1137),
.Y(n_1265)
);

BUFx2_ASAP7_75t_SL g1266 ( 
.A(n_1241),
.Y(n_1266)
);

BUFx2_ASAP7_75t_SL g1267 ( 
.A(n_1218),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1177),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1221),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1218),
.Y(n_1270)
);

BUFx2_ASAP7_75t_SL g1271 ( 
.A(n_1240),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1198),
.A2(n_1170),
.B1(n_1211),
.B2(n_1135),
.Y(n_1272)
);

BUFx8_ASAP7_75t_SL g1273 ( 
.A(n_1240),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1119),
.A2(n_1164),
.B1(n_1176),
.B2(n_1125),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1141),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1122),
.A2(n_1206),
.B1(n_1185),
.B2(n_1181),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_1208),
.Y(n_1277)
);

INVx6_ASAP7_75t_L g1278 ( 
.A(n_1177),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1148),
.Y(n_1279)
);

INVx6_ASAP7_75t_L g1280 ( 
.A(n_1239),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1190),
.Y(n_1281)
);

AOI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1164),
.A2(n_1181),
.B1(n_1185),
.B2(n_1142),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1150),
.Y(n_1283)
);

CKINVDCx11_ASAP7_75t_R g1284 ( 
.A(n_1240),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1237),
.A2(n_1189),
.B1(n_1121),
.B2(n_1159),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1147),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1204),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1190),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1216),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1181),
.A2(n_1185),
.B1(n_1189),
.B2(n_1131),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1190),
.Y(n_1291)
);

BUFx8_ASAP7_75t_SL g1292 ( 
.A(n_1229),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1120),
.A2(n_1182),
.B1(n_1243),
.B2(n_1223),
.Y(n_1293)
);

OAI21xp33_ASAP7_75t_L g1294 ( 
.A1(n_1173),
.A2(n_1158),
.B(n_1146),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1246),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1161),
.A2(n_1207),
.B1(n_1133),
.B2(n_1174),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1121),
.A2(n_1158),
.B1(n_1217),
.B2(n_1233),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1191),
.B(n_1167),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_SL g1299 ( 
.A1(n_1139),
.A2(n_1144),
.B1(n_1197),
.B2(n_1171),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1133),
.A2(n_1155),
.B1(n_1180),
.B2(n_1138),
.Y(n_1300)
);

AOI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1236),
.A2(n_1108),
.B1(n_1225),
.B2(n_1219),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1166),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1166),
.Y(n_1303)
);

BUFx8_ASAP7_75t_L g1304 ( 
.A(n_1192),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1175),
.A2(n_1179),
.B1(n_1184),
.B2(n_1124),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1124),
.A2(n_1162),
.B1(n_1194),
.B2(n_1168),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1166),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_1201),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1197),
.A2(n_1196),
.B1(n_1123),
.B2(n_1143),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1231),
.A2(n_1108),
.B1(n_1210),
.B2(n_1232),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1187),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1132),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1200),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1169),
.A2(n_1151),
.B1(n_1115),
.B2(n_1149),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1186),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1126),
.A2(n_1202),
.B1(n_1215),
.B2(n_1195),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1113),
.A2(n_1112),
.B1(n_1231),
.B2(n_1117),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1193),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1116),
.A2(n_1118),
.B1(n_1136),
.B2(n_1245),
.Y(n_1319)
);

INVx2_ASAP7_75t_SL g1320 ( 
.A(n_1193),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1186),
.B(n_1231),
.Y(n_1321)
);

CKINVDCx11_ASAP7_75t_R g1322 ( 
.A(n_1160),
.Y(n_1322)
);

CKINVDCx11_ASAP7_75t_R g1323 ( 
.A(n_1160),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_SL g1324 ( 
.A1(n_1244),
.A2(n_1156),
.B1(n_1227),
.B2(n_1222),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1160),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1213),
.A2(n_1156),
.B1(n_1157),
.B2(n_1107),
.Y(n_1326)
);

CKINVDCx6p67_ASAP7_75t_R g1327 ( 
.A(n_1157),
.Y(n_1327)
);

CKINVDCx20_ASAP7_75t_R g1328 ( 
.A(n_1157),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1230),
.B(n_1128),
.Y(n_1329)
);

INVx5_ASAP7_75t_L g1330 ( 
.A(n_1128),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1156),
.A2(n_1107),
.B1(n_1109),
.B2(n_1128),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1107),
.A2(n_1212),
.B1(n_1074),
.B2(n_1226),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1109),
.A2(n_1119),
.B(n_1210),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1109),
.A2(n_1074),
.B1(n_1072),
.B2(n_412),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1226),
.A2(n_1074),
.B1(n_1072),
.B2(n_1051),
.Y(n_1337)
);

INVx5_ASAP7_75t_L g1338 ( 
.A(n_1190),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1226),
.A2(n_1074),
.B1(n_1072),
.B2(n_1051),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1226),
.A2(n_1153),
.B1(n_671),
.B2(n_1110),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1147),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1183),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1129),
.Y(n_1344)
);

AOI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1226),
.A2(n_436),
.B1(n_336),
.B2(n_329),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1129),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1129),
.Y(n_1347)
);

INVx2_ASAP7_75t_SL g1348 ( 
.A(n_1147),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1183),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_1190),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1183),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1153),
.A2(n_1074),
.B1(n_1072),
.B2(n_412),
.Y(n_1354)
);

BUFx10_ASAP7_75t_L g1355 ( 
.A(n_1218),
.Y(n_1355)
);

BUFx12f_ASAP7_75t_L g1356 ( 
.A(n_1183),
.Y(n_1356)
);

OAI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1226),
.A2(n_1110),
.B1(n_1153),
.B2(n_1074),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1226),
.A2(n_1153),
.B1(n_671),
.B2(n_1110),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1207),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1183),
.Y(n_1360)
);

INVx4_ASAP7_75t_SL g1361 ( 
.A(n_1193),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1177),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1159),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1129),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1183),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1226),
.A2(n_1153),
.B1(n_671),
.B2(n_1110),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1226),
.A2(n_1110),
.B1(n_1153),
.B2(n_1074),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1226),
.A2(n_436),
.B1(n_336),
.B2(n_329),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_1211),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1159),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1212),
.A2(n_1074),
.B1(n_1226),
.B2(n_1205),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1153),
.A2(n_1074),
.B1(n_1072),
.B2(n_412),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1183),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1154),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1333),
.A2(n_1317),
.B(n_1325),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1333),
.A2(n_1319),
.B(n_1316),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1329),
.A2(n_1314),
.B(n_1306),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1302),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1303),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1307),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1260),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1311),
.Y(n_1383)
);

HB1xp67_ASAP7_75t_L g1384 ( 
.A(n_1370),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1318),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1370),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1260),
.Y(n_1387)
);

INVx2_ASAP7_75t_SL g1388 ( 
.A(n_1311),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1315),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1256),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1313),
.Y(n_1391)
);

HB1xp67_ASAP7_75t_L g1392 ( 
.A(n_1258),
.Y(n_1392)
);

OAI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1250),
.A2(n_1358),
.B(n_1341),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1300),
.A2(n_1317),
.B(n_1326),
.Y(n_1394)
);

AO21x1_ASAP7_75t_L g1395 ( 
.A1(n_1357),
.A2(n_1368),
.B(n_1247),
.Y(n_1395)
);

BUFx3_ASAP7_75t_L g1396 ( 
.A(n_1298),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1321),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1337),
.A2(n_1339),
.B1(n_1368),
.B2(n_1357),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1248),
.A2(n_1373),
.B1(n_1354),
.B2(n_1353),
.Y(n_1399)
);

AOI21xp33_ASAP7_75t_L g1400 ( 
.A1(n_1367),
.A2(n_1339),
.B(n_1337),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1331),
.A2(n_1309),
.B(n_1274),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1320),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1361),
.Y(n_1403)
);

OAI21x1_ASAP7_75t_L g1404 ( 
.A1(n_1296),
.A2(n_1264),
.B(n_1276),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1263),
.A2(n_1290),
.B(n_1305),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1361),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1299),
.A2(n_1248),
.B(n_1297),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1354),
.A2(n_1373),
.B(n_1336),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1330),
.B(n_1301),
.Y(n_1409)
);

INVx2_ASAP7_75t_SL g1410 ( 
.A(n_1311),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1335),
.A2(n_1364),
.B1(n_1340),
.B2(n_1372),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1330),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1294),
.A2(n_1254),
.B(n_1293),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1328),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1327),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1259),
.Y(n_1416)
);

NAND2x1_ASAP7_75t_L g1417 ( 
.A(n_1313),
.B(n_1278),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1352),
.A2(n_1285),
.B(n_1334),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1262),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1265),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1279),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1283),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1287),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1289),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1295),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1344),
.A2(n_1347),
.B(n_1346),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1365),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1322),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1332),
.B(n_1285),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1323),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1359),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1298),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1324),
.A2(n_1261),
.B(n_1310),
.Y(n_1433)
);

OA21x2_ASAP7_75t_L g1434 ( 
.A1(n_1255),
.A2(n_1324),
.B(n_1310),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1297),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1312),
.A2(n_1272),
.B(n_1299),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1375),
.Y(n_1437)
);

INVx3_ASAP7_75t_L g1438 ( 
.A(n_1313),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1308),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1334),
.A2(n_1345),
.B(n_1369),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1278),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1304),
.Y(n_1442)
);

INVx4_ASAP7_75t_L g1443 ( 
.A(n_1338),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1268),
.B(n_1282),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1304),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1280),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1362),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1362),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1291),
.B(n_1288),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1291),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1257),
.B(n_1348),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1342),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1281),
.A2(n_1350),
.B(n_1288),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1286),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1355),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1251),
.A2(n_1363),
.B1(n_1371),
.B2(n_1266),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1355),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1249),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1249),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1270),
.Y(n_1461)
);

BUFx12f_ASAP7_75t_L g1462 ( 
.A(n_1442),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_L g1463 ( 
.A(n_1396),
.B(n_1277),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1390),
.Y(n_1464)
);

NOR2x1_ASAP7_75t_SL g1465 ( 
.A(n_1436),
.B(n_1360),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1393),
.A2(n_1253),
.B(n_1275),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1396),
.B(n_1252),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1400),
.A2(n_1284),
.B1(n_1273),
.B2(n_1374),
.C(n_1366),
.Y(n_1468)
);

OR2x6_ASAP7_75t_L g1469 ( 
.A(n_1404),
.B(n_1349),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_SL g1470 ( 
.A1(n_1440),
.A2(n_1343),
.B(n_1351),
.C(n_1269),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1435),
.B(n_1292),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_SL g1472 ( 
.A1(n_1408),
.A2(n_1418),
.B(n_1428),
.C(n_1430),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1416),
.Y(n_1473)
);

OA21x2_ASAP7_75t_L g1474 ( 
.A1(n_1377),
.A2(n_1356),
.B(n_1404),
.Y(n_1474)
);

AO32x2_ASAP7_75t_L g1475 ( 
.A1(n_1383),
.A2(n_1410),
.A3(n_1388),
.B1(n_1441),
.B2(n_1397),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1407),
.A2(n_1398),
.B(n_1413),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1419),
.Y(n_1477)
);

NOR2x1_ASAP7_75t_SL g1478 ( 
.A(n_1436),
.B(n_1454),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1414),
.B(n_1397),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1396),
.B(n_1415),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_1451),
.Y(n_1481)
);

NOR2x1_ASAP7_75t_SL g1482 ( 
.A(n_1436),
.B(n_1454),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_L g1483 ( 
.A(n_1398),
.B(n_1399),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1439),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1411),
.A2(n_1429),
.B1(n_1385),
.B2(n_1428),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1397),
.B(n_1385),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1413),
.A2(n_1405),
.B(n_1429),
.C(n_1401),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1384),
.B(n_1386),
.Y(n_1488)
);

OA21x2_ASAP7_75t_L g1489 ( 
.A1(n_1394),
.A2(n_1378),
.B(n_1379),
.Y(n_1489)
);

O2A1O1Ixp5_ASAP7_75t_L g1490 ( 
.A1(n_1395),
.A2(n_1417),
.B(n_1430),
.C(n_1444),
.Y(n_1490)
);

BUFx4f_ASAP7_75t_L g1491 ( 
.A(n_1454),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1422),
.B(n_1424),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1439),
.A2(n_1437),
.B1(n_1392),
.B2(n_1445),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1424),
.B(n_1420),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1395),
.A2(n_1417),
.B(n_1432),
.C(n_1410),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1433),
.A2(n_1452),
.B1(n_1427),
.B2(n_1425),
.C(n_1423),
.Y(n_1496)
);

AOI221xp5_ASAP7_75t_L g1497 ( 
.A1(n_1433),
.A2(n_1452),
.B1(n_1427),
.B2(n_1425),
.C(n_1421),
.Y(n_1497)
);

AOI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1444),
.A2(n_1457),
.B1(n_1461),
.B2(n_1438),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1451),
.B(n_1461),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1426),
.B(n_1450),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1455),
.Y(n_1501)
);

OR2x6_ASAP7_75t_L g1502 ( 
.A(n_1409),
.B(n_1403),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1426),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1449),
.B(n_1431),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1459),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_SL g1506 ( 
.A1(n_1442),
.A2(n_1445),
.B1(n_1459),
.B2(n_1460),
.Y(n_1506)
);

NOR2x1_ASAP7_75t_SL g1507 ( 
.A(n_1454),
.B(n_1433),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_R g1508 ( 
.A(n_1460),
.B(n_1446),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1378),
.A2(n_1380),
.B(n_1381),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1434),
.A2(n_1391),
.B(n_1438),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1382),
.B(n_1387),
.Y(n_1511)
);

OR2x6_ASAP7_75t_L g1512 ( 
.A(n_1409),
.B(n_1406),
.Y(n_1512)
);

BUFx3_ASAP7_75t_L g1513 ( 
.A(n_1502),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1489),
.B(n_1376),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1476),
.A2(n_1434),
.B1(n_1459),
.B2(n_1458),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1492),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1486),
.B(n_1376),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1509),
.Y(n_1518)
);

INVx4_ASAP7_75t_L g1519 ( 
.A(n_1491),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1483),
.A2(n_1476),
.B1(n_1485),
.B2(n_1466),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1479),
.B(n_1376),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1503),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1509),
.B(n_1434),
.Y(n_1523)
);

AND2x4_ASAP7_75t_SL g1524 ( 
.A(n_1502),
.B(n_1412),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1511),
.B(n_1484),
.Y(n_1525)
);

OR2x2_ASAP7_75t_SL g1526 ( 
.A(n_1474),
.B(n_1434),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1488),
.B(n_1389),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1500),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1485),
.A2(n_1391),
.B1(n_1456),
.B2(n_1448),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1473),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1477),
.Y(n_1531)
);

BUFx3_ASAP7_75t_L g1532 ( 
.A(n_1512),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1494),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1507),
.B(n_1381),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1475),
.B(n_1389),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1493),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1494),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1475),
.B(n_1389),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1475),
.B(n_1402),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1466),
.A2(n_1391),
.B1(n_1456),
.B2(n_1447),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1530),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1530),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1535),
.B(n_1478),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1513),
.B(n_1482),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1513),
.B(n_1532),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1513),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1517),
.B(n_1488),
.Y(n_1547)
);

INVx5_ASAP7_75t_L g1548 ( 
.A(n_1523),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1535),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1518),
.A2(n_1487),
.B(n_1465),
.Y(n_1550)
);

AOI33xp33_ASAP7_75t_L g1551 ( 
.A1(n_1520),
.A2(n_1472),
.A3(n_1497),
.B1(n_1496),
.B2(n_1470),
.B3(n_1481),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1530),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1522),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1537),
.B(n_1496),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1519),
.B(n_1469),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1520),
.A2(n_1490),
.B(n_1495),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1535),
.B(n_1497),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1537),
.B(n_1510),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1531),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1538),
.B(n_1474),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1561)
);

INVx1_ASAP7_75t_SL g1562 ( 
.A(n_1525),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1513),
.B(n_1532),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1519),
.Y(n_1564)
);

NAND2x1_ASAP7_75t_L g1565 ( 
.A(n_1538),
.B(n_1480),
.Y(n_1565)
);

OAI222xp33_ASAP7_75t_L g1566 ( 
.A1(n_1529),
.A2(n_1463),
.B1(n_1536),
.B2(n_1498),
.C1(n_1515),
.C2(n_1540),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1536),
.B(n_1508),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

NOR2x1_ASAP7_75t_L g1569 ( 
.A(n_1515),
.B(n_1527),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1523),
.B(n_1504),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1554),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1549),
.B(n_1521),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.B(n_1523),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1557),
.B(n_1537),
.Y(n_1574)
);

AND4x1_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1468),
.C(n_1540),
.D(n_1529),
.Y(n_1575)
);

INVxp67_ASAP7_75t_SL g1576 ( 
.A(n_1558),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1541),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1541),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1553),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1553),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1557),
.B(n_1554),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1543),
.B(n_1539),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1543),
.B(n_1539),
.Y(n_1583)
);

INVxp67_ASAP7_75t_SL g1584 ( 
.A(n_1558),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1542),
.Y(n_1585)
);

INVx6_ASAP7_75t_L g1586 ( 
.A(n_1548),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1539),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1542),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1553),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1552),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1560),
.B(n_1534),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1560),
.B(n_1548),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1568),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1560),
.B(n_1534),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1548),
.B(n_1534),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1548),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1548),
.B(n_1524),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1548),
.B(n_1514),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1548),
.B(n_1514),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1557),
.B(n_1533),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1562),
.B(n_1533),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1562),
.B(n_1516),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1559),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1590),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1590),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1577),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1576),
.B(n_1547),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1571),
.B(n_1569),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1563),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1577),
.Y(n_1612)
);

NOR2x1p5_ASAP7_75t_L g1613 ( 
.A(n_1581),
.B(n_1564),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1577),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1592),
.B(n_1545),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1578),
.Y(n_1616)
);

OR2x6_ASAP7_75t_L g1617 ( 
.A(n_1586),
.B(n_1556),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1571),
.B(n_1581),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1578),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1578),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1575),
.B(n_1462),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1582),
.B(n_1545),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1585),
.Y(n_1625)
);

HB1xp67_ASAP7_75t_L g1626 ( 
.A(n_1600),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1576),
.B(n_1569),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1579),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1575),
.B(n_1471),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1597),
.B(n_1544),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1582),
.B(n_1583),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1584),
.B(n_1600),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1584),
.B(n_1556),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1585),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1579),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1588),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1579),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1574),
.B(n_1561),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1574),
.A2(n_1555),
.B1(n_1564),
.B2(n_1545),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1602),
.B(n_1561),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1588),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1583),
.B(n_1545),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1591),
.B(n_1546),
.Y(n_1646)
);

INVxp33_ASAP7_75t_SL g1647 ( 
.A(n_1622),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1607),
.B(n_1591),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1591),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1608),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1607),
.B(n_1594),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1594),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1608),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1633),
.B(n_1594),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1618),
.B(n_1471),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1612),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1617),
.B(n_1467),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1546),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1619),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1595),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1640),
.B(n_1601),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1613),
.B(n_1596),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1595),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1612),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1614),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1467),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1617),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1614),
.Y(n_1670)
);

OAI21xp33_ASAP7_75t_L g1671 ( 
.A1(n_1617),
.A2(n_1599),
.B(n_1598),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1632),
.B(n_1601),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1617),
.B(n_1499),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1642),
.B(n_1572),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1624),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1626),
.B(n_1570),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1631),
.B(n_1595),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1627),
.B(n_1570),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1631),
.B(n_1587),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1609),
.B(n_1645),
.Y(n_1681)
);

AOI222xp33_ASAP7_75t_L g1682 ( 
.A1(n_1647),
.A2(n_1566),
.B1(n_1468),
.B2(n_1641),
.C1(n_1615),
.C2(n_1587),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1656),
.B(n_1646),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_SL g1684 ( 
.A(n_1647),
.B(n_1566),
.Y(n_1684)
);

NAND2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1649),
.B(n_1565),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

AOI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1659),
.A2(n_1615),
.B1(n_1630),
.B2(n_1550),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1668),
.B(n_1623),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1673),
.A2(n_1526),
.B1(n_1586),
.B2(n_1630),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_L g1690 ( 
.A1(n_1669),
.A2(n_1606),
.B1(n_1605),
.B2(n_1609),
.C(n_1464),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1660),
.B(n_1506),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1648),
.B(n_1646),
.Y(n_1692)
);

AOI221xp5_ASAP7_75t_L g1693 ( 
.A1(n_1671),
.A2(n_1606),
.B1(n_1605),
.B2(n_1643),
.C(n_1638),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1662),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1681),
.B(n_1623),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1674),
.Y(n_1698)
);

NAND2x1_ASAP7_75t_SL g1699 ( 
.A(n_1661),
.B(n_1596),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1676),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1681),
.B(n_1644),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1653),
.Y(n_1702)
);

AOI22xp5_ASAP7_75t_L g1703 ( 
.A1(n_1655),
.A2(n_1630),
.B1(n_1550),
.B2(n_1544),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1658),
.Y(n_1704)
);

AOI21xp33_ASAP7_75t_L g1705 ( 
.A1(n_1661),
.A2(n_1619),
.B(n_1550),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1655),
.B(n_1564),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1684),
.A2(n_1664),
.B1(n_1655),
.B2(n_1676),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1700),
.Y(n_1708)
);

NAND4xp25_ASAP7_75t_SL g1709 ( 
.A(n_1682),
.B(n_1654),
.C(n_1662),
.D(n_1678),
.Y(n_1709)
);

AO22x1_ASAP7_75t_L g1710 ( 
.A1(n_1691),
.A2(n_1661),
.B1(n_1664),
.B2(n_1596),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1690),
.B(n_1648),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1686),
.Y(n_1712)
);

AOI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_1685),
.A2(n_1664),
.B1(n_1630),
.B2(n_1679),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1694),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1690),
.B(n_1683),
.Y(n_1715)
);

OAI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1697),
.A2(n_1586),
.B1(n_1619),
.B2(n_1651),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1706),
.A2(n_1586),
.B1(n_1678),
.B2(n_1665),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1696),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1644),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1698),
.Y(n_1720)
);

NAND4xp25_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1672),
.C(n_1675),
.D(n_1665),
.Y(n_1721)
);

INVx2_ASAP7_75t_SL g1722 ( 
.A(n_1699),
.Y(n_1722)
);

OAI22xp5_ASAP7_75t_L g1723 ( 
.A1(n_1701),
.A2(n_1586),
.B1(n_1651),
.B2(n_1652),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_L g1724 ( 
.A1(n_1693),
.A2(n_1550),
.B1(n_1652),
.B2(n_1666),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1702),
.Y(n_1725)
);

BUFx2_ASAP7_75t_L g1726 ( 
.A(n_1722),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1718),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1718),
.Y(n_1728)
);

OAI21xp33_ASAP7_75t_L g1729 ( 
.A1(n_1715),
.A2(n_1695),
.B(n_1692),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1724),
.B(n_1687),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1708),
.Y(n_1731)
);

OAI21xp33_ASAP7_75t_L g1732 ( 
.A1(n_1707),
.A2(n_1703),
.B(n_1704),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1712),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1714),
.Y(n_1734)
);

NOR4xp25_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1696),
.C(n_1705),
.D(n_1689),
.Y(n_1735)
);

AOI32xp33_ASAP7_75t_L g1736 ( 
.A1(n_1711),
.A2(n_1680),
.A3(n_1667),
.B1(n_1670),
.B2(n_1599),
.Y(n_1736)
);

NAND2xp33_ASAP7_75t_SL g1737 ( 
.A(n_1725),
.B(n_1657),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1720),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1726),
.Y(n_1739)
);

NAND3xp33_ASAP7_75t_SL g1740 ( 
.A(n_1735),
.B(n_1717),
.C(n_1713),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1727),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1737),
.B(n_1736),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1743)
);

INVxp33_ASAP7_75t_L g1744 ( 
.A(n_1732),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1737),
.A2(n_1721),
.B(n_1716),
.C(n_1723),
.Y(n_1745)
);

INVx3_ASAP7_75t_L g1746 ( 
.A(n_1731),
.Y(n_1746)
);

OAI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1730),
.A2(n_1719),
.B(n_1672),
.Y(n_1747)
);

CKINVDCx6p67_ASAP7_75t_R g1748 ( 
.A(n_1741),
.Y(n_1748)
);

AOI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1740),
.A2(n_1730),
.B1(n_1710),
.B2(n_1734),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_SL g1750 ( 
.A1(n_1745),
.A2(n_1733),
.B1(n_1663),
.B2(n_1657),
.C(n_1675),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1739),
.B(n_1680),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1744),
.A2(n_1663),
.B1(n_1677),
.B2(n_1637),
.C(n_1639),
.Y(n_1752)
);

AOI222xp33_ASAP7_75t_L g1753 ( 
.A1(n_1752),
.A2(n_1742),
.B1(n_1743),
.B2(n_1747),
.C1(n_1738),
.C2(n_1746),
.Y(n_1753)
);

OAI311xp33_ASAP7_75t_L g1754 ( 
.A1(n_1749),
.A2(n_1746),
.A3(n_1572),
.B1(n_1501),
.C1(n_1599),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1750),
.A2(n_1586),
.B1(n_1555),
.B2(n_1639),
.C(n_1628),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1748),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1751),
.A2(n_1643),
.B(n_1638),
.Y(n_1757)
);

AO22x2_ASAP7_75t_L g1758 ( 
.A1(n_1751),
.A2(n_1620),
.B1(n_1636),
.B2(n_1635),
.Y(n_1758)
);

AOI22x1_ASAP7_75t_L g1759 ( 
.A1(n_1753),
.A2(n_1637),
.B1(n_1628),
.B2(n_1635),
.Y(n_1759)
);

INVx5_ASAP7_75t_L g1760 ( 
.A(n_1756),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1755),
.B(n_1572),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1757),
.B(n_1616),
.Y(n_1762)
);

AOI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1758),
.A2(n_1586),
.B1(n_1597),
.B2(n_1621),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1761),
.B(n_1754),
.Y(n_1764)
);

NOR3xp33_ASAP7_75t_L g1765 ( 
.A(n_1760),
.B(n_1637),
.C(n_1567),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1762),
.A2(n_1636),
.B1(n_1634),
.B2(n_1620),
.C(n_1625),
.Y(n_1766)
);

NAND2x1p5_ASAP7_75t_L g1767 ( 
.A(n_1764),
.B(n_1759),
.Y(n_1767)
);

AOI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1767),
.A2(n_1765),
.B1(n_1763),
.B2(n_1766),
.Y(n_1768)
);

OAI22x1_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1634),
.B1(n_1625),
.B2(n_1621),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1768),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1770),
.A2(n_1598),
.B1(n_1597),
.B2(n_1573),
.Y(n_1771)
);

AOI22x1_ASAP7_75t_L g1772 ( 
.A1(n_1769),
.A2(n_1598),
.B1(n_1589),
.B2(n_1593),
.Y(n_1772)
);

AOI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1573),
.B(n_1589),
.Y(n_1773)
);

AO22x2_ASAP7_75t_L g1774 ( 
.A1(n_1771),
.A2(n_1589),
.B1(n_1580),
.B2(n_1579),
.Y(n_1774)
);

OAI21xp5_ASAP7_75t_L g1775 ( 
.A1(n_1773),
.A2(n_1573),
.B(n_1603),
.Y(n_1775)
);

OAI222xp33_ASAP7_75t_SL g1776 ( 
.A1(n_1775),
.A2(n_1774),
.B1(n_1519),
.B2(n_1443),
.C1(n_1603),
.C2(n_1604),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1580),
.B1(n_1589),
.B2(n_1593),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_R g1778 ( 
.A1(n_1777),
.A2(n_1580),
.B1(n_1593),
.B2(n_1587),
.C(n_1597),
.Y(n_1778)
);

AOI211xp5_ASAP7_75t_L g1779 ( 
.A1(n_1778),
.A2(n_1453),
.B(n_1505),
.C(n_1441),
.Y(n_1779)
);


endmodule