module fake_netlist_1_3088_n_43 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_43);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_43;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_6), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_5), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_1), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_10), .Y(n_21) );
BUFx4f_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
CKINVDCx5p33_ASAP7_75t_R g23 ( .A(n_16), .Y(n_23) );
O2A1O1Ixp33_ASAP7_75t_L g24 ( .A1(n_20), .A2(n_1), .B(n_2), .C(n_3), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_19), .Y(n_25) );
INVx3_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
OAI21x1_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_21), .B(n_15), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_23), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_27), .Y(n_33) );
AOI21xp33_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_30), .B(n_27), .Y(n_34) );
OAI221xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_22), .B1(n_18), .B2(n_17), .C(n_2), .Y(n_35) );
AOI22xp33_ASAP7_75t_L g36 ( .A1(n_32), .A2(n_22), .B1(n_18), .B2(n_3), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
NAND3xp33_ASAP7_75t_L g38 ( .A(n_36), .B(n_4), .C(n_7), .Y(n_38) );
INVxp67_ASAP7_75t_L g39 ( .A(n_34), .Y(n_39) );
OR4x1_ASAP7_75t_L g40 ( .A(n_39), .B(n_8), .C(n_11), .D(n_12), .Y(n_40) );
XNOR2xp5_ASAP7_75t_L g41 ( .A(n_37), .B(n_13), .Y(n_41) );
OAI22xp5_ASAP7_75t_L g42 ( .A1(n_41), .A2(n_38), .B1(n_40), .B2(n_14), .Y(n_42) );
BUFx2_ASAP7_75t_L g43 ( .A(n_42), .Y(n_43) );
endmodule