module fake_jpeg_29466_n_239 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_20),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_34),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_28),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_29),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_53),
.Y(n_81)
);

O2A1O1Ixp33_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_31),
.B(n_17),
.C(n_19),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_52),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_29),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_31),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_33),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_31),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_19),
.B1(n_14),
.B2(n_23),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_63),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_35),
.A2(n_15),
.B(n_26),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_42),
.A2(n_14),
.B1(n_23),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_24),
.B1(n_44),
.B2(n_21),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_36),
.A2(n_19),
.B1(n_21),
.B2(n_18),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_35),
.B1(n_26),
.B2(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_75),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_42),
.B1(n_43),
.B2(n_40),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_79),
.B1(n_84),
.B2(n_86),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_87),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_23),
.B1(n_14),
.B2(n_24),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_23),
.B1(n_14),
.B2(n_24),
.Y(n_86)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_27),
.C(n_25),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_51),
.C(n_63),
.Y(n_111)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_54),
.B(n_25),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_103),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_95),
.Y(n_120)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_44),
.B1(n_31),
.B2(n_16),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_102),
.B1(n_105),
.B2(n_48),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_60),
.A2(n_44),
.B1(n_22),
.B2(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_104),
.Y(n_112)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_62),
.A2(n_22),
.B1(n_16),
.B2(n_44),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_31),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_67),
.B(n_1),
.C(n_2),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_111),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_127),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_115),
.A2(n_105),
.B1(n_77),
.B2(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_124),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_82),
.B(n_10),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_122),
.B(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_92),
.B(n_50),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_125),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_73),
.B(n_104),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_59),
.Y(n_127)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR3xp33_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_59),
.C(n_8),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_96),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_76),
.B(n_100),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_147),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_138),
.A2(n_156),
.B1(n_159),
.B2(n_108),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_144),
.B(n_149),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_101),
.C(n_87),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_152),
.C(n_158),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_95),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_68),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_130),
.A2(n_74),
.B(n_93),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_153),
.A2(n_120),
.B(n_125),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_72),
.B1(n_91),
.B2(n_98),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_130),
.A2(n_58),
.B1(n_93),
.B2(n_56),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_157),
.A2(n_109),
.B1(n_136),
.B2(n_107),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_80),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_160),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_58),
.B1(n_48),
.B2(n_80),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_59),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_122),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_168),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_143),
.B(n_133),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_164),
.B(n_154),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_109),
.B1(n_108),
.B2(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_165),
.A2(n_170),
.B1(n_175),
.B2(n_178),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_160),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_113),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_174),
.C(n_179),
.Y(n_180)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_140),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_153),
.B(n_149),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_173),
.A2(n_159),
.B1(n_139),
.B2(n_155),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_113),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_131),
.B1(n_119),
.B2(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_144),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_131),
.B1(n_119),
.B2(n_123),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_134),
.C(n_121),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_166),
.B(n_169),
.C(n_173),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g182 ( 
.A1(n_166),
.A2(n_146),
.B(n_139),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_129),
.B1(n_128),
.B2(n_121),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_187),
.C(n_193),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_194),
.B1(n_178),
.B2(n_170),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_142),
.C(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_142),
.A3(n_147),
.B1(n_137),
.B2(n_157),
.C1(n_120),
.C2(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_190),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_164),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_154),
.Y(n_193)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_167),
.A2(n_120),
.B1(n_151),
.B2(n_129),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_151),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_179),
.C(n_174),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_180),
.C(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_183),
.C(n_198),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_206),
.B(n_207),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_176),
.Y(n_202)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_203),
.A2(n_208),
.B1(n_184),
.B2(n_186),
.Y(n_214)
);

AO22x1_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_175),
.B1(n_120),
.B2(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_204),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_131),
.Y(n_205)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_205),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_192),
.B(n_74),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_128),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_210),
.C(n_199),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_198),
.B(n_180),
.C(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_215),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_214),
.A2(n_212),
.B1(n_204),
.B2(n_211),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_201),
.B(n_194),
.C(n_185),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_218),
.A2(n_221),
.B1(n_10),
.B2(n_9),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_217),
.A2(n_200),
.B1(n_196),
.B2(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

OAI21x1_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_222),
.B(n_224),
.Y(n_228)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_202),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_200),
.B(n_11),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_200),
.B(n_48),
.Y(n_225)
);

AOI21x1_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_229),
.B(n_228),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_221),
.C(n_218),
.Y(n_232)
);

AOI31xp67_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_10),
.A3(n_8),
.B(n_2),
.Y(n_229)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_220),
.C(n_224),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_232),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_48),
.B(n_1),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g237 ( 
.A1(n_234),
.A2(n_4),
.B(n_5),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g236 ( 
.A1(n_235),
.A2(n_0),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_237),
.B(n_233),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_6),
.B(n_7),
.Y(n_239)
);


endmodule