module fake_jpeg_26940_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_32),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_35),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_22),
.B(n_9),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_41),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_27),
.B1(n_25),
.B2(n_28),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_50),
.B1(n_33),
.B2(n_19),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_34),
.A2(n_27),
.B1(n_17),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_58),
.B1(n_18),
.B2(n_31),
.Y(n_60)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_17),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_27),
.B1(n_25),
.B2(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_24),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_33),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_32),
.B1(n_30),
.B2(n_16),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_63),
.B1(n_59),
.B2(n_44),
.Y(n_99)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_64),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_29),
.B1(n_30),
.B2(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_20),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_57),
.Y(n_65)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_20),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_75),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_69),
.B(n_55),
.Y(n_117)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_37),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_54),
.B(n_51),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_30),
.B1(n_16),
.B2(n_23),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_48),
.B1(n_55),
.B2(n_3),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_30),
.B2(n_23),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_76),
.B1(n_55),
.B2(n_54),
.Y(n_107)
);

NOR4xp25_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_12),
.C(n_15),
.D(n_14),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_85),
.Y(n_95)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_74),
.A2(n_82),
.B1(n_91),
.B2(n_55),
.Y(n_102)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_42),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_21),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_79),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_81),
.Y(n_116)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_21),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

OA22x2_ASAP7_75t_SL g89 ( 
.A1(n_42),
.A2(n_41),
.B1(n_21),
.B2(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_9),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_52),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_89),
.B1(n_81),
.B2(n_87),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_95),
.B1(n_76),
.B2(n_94),
.Y(n_143)
);

A2O1A1Ixp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_79),
.B(n_70),
.C(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_104),
.B(n_109),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_106),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_117),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_69),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_70),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_89),
.B(n_61),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_92),
.A2(n_62),
.B1(n_109),
.B2(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_119),
.A2(n_127),
.B1(n_129),
.B2(n_144),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_118),
.B(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_135),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_92),
.A2(n_80),
.B1(n_70),
.B2(n_66),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_107),
.B1(n_106),
.B2(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_134),
.Y(n_166)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_98),
.B(n_93),
.Y(n_172)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_61),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_108),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_139),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_99),
.A2(n_89),
.B1(n_73),
.B2(n_75),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_138),
.A2(n_143),
.B1(n_107),
.B2(n_101),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_97),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_142),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_111),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_83),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_96),
.B(n_77),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_93),
.Y(n_173)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_148),
.A2(n_171),
.B(n_172),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_101),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_149),
.B(n_157),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_150),
.A2(n_153),
.B1(n_138),
.B2(n_122),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_103),
.B1(n_110),
.B2(n_100),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_130),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_173),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_83),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_83),
.B(n_6),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_158),
.B(n_159),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_125),
.B(n_103),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_162),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_100),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_122),
.C(n_129),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_100),
.B1(n_98),
.B2(n_67),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_167),
.A2(n_120),
.B1(n_139),
.B2(n_126),
.Y(n_196)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_170),
.Y(n_199)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_147),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_133),
.A2(n_98),
.B(n_112),
.Y(n_171)
);

OA21x2_ASAP7_75t_SL g174 ( 
.A1(n_140),
.A2(n_12),
.B(n_14),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_11),
.B(n_15),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_1),
.B(n_2),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_175),
.A2(n_142),
.B(n_134),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_132),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g193 ( 
.A(n_176),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_122),
.B(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_180),
.Y(n_201)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_162),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_181),
.B(n_182),
.Y(n_217)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_186),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_122),
.B(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_187),
.A2(n_195),
.B1(n_197),
.B2(n_175),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_200),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_121),
.B1(n_128),
.B2(n_123),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_189),
.A2(n_196),
.B1(n_150),
.B2(n_153),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_149),
.C(n_164),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_126),
.B1(n_74),
.B2(n_120),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_205),
.B(n_209),
.Y(n_230)
);

AOI22x1_ASAP7_75t_L g206 ( 
.A1(n_190),
.A2(n_171),
.B1(n_164),
.B2(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_206),
.A2(n_218),
.B1(n_181),
.B2(n_180),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_193),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_179),
.B(n_187),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_196),
.A2(n_169),
.B1(n_159),
.B2(n_155),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_166),
.B1(n_170),
.B2(n_138),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_151),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_214),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_151),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_161),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_199),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_183),
.B(n_174),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_177),
.C(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_225),
.Y(n_238)
);

NOR2x1_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_227),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_226),
.A2(n_112),
.B1(n_93),
.B2(n_54),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_208),
.B(n_212),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_179),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_203),
.C(n_213),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_233),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_198),
.Y(n_233)
);

A2O1A1O1Ixp25_ASAP7_75t_L g234 ( 
.A1(n_219),
.A2(n_186),
.B(n_184),
.C(n_185),
.D(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_200),
.Y(n_244)
);

FAx1_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_5),
.CI(n_6),
.CON(n_256),
.SN(n_256)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_223),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_228),
.B(n_214),
.C(n_215),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_242),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_207),
.B1(n_204),
.B2(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_245),
.B1(n_246),
.B2(n_230),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_185),
.C(n_202),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_244),
.A2(n_5),
.B(n_6),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_229),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_220),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_251),
.B(n_253),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_243),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_248),
.B(n_238),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_256),
.B1(n_246),
.B2(n_245),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_225),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_250),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_231),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_255),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_240),
.A2(n_234),
.B(n_4),
.C(n_5),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_236),
.B(n_238),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_259),
.C(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_237),
.C(n_239),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_247),
.Y(n_265)
);

INVxp33_ASAP7_75t_SL g264 ( 
.A(n_258),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_264),
.A2(n_266),
.B(n_260),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_263),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_259),
.B(n_10),
.Y(n_267)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_267),
.A2(n_260),
.A3(n_258),
.B1(n_11),
.B2(n_15),
.C1(n_10),
.C2(n_1),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_269),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_270),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_268),
.Y(n_272)
);

AOI321xp33_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_271),
.A3(n_274),
.B1(n_272),
.B2(n_10),
.C(n_51),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_275),
.B(n_1),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_51),
.B(n_200),
.Y(n_277)
);


endmodule