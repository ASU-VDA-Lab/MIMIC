module real_jpeg_20703_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_277, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_277;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_1),
.A2(n_2),
.B1(n_18),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_1),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_61),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_61),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_1),
.A2(n_61),
.B1(n_72),
.B2(n_73),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_2),
.A2(n_4),
.B1(n_17),
.B2(n_18),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_2),
.A2(n_8),
.B1(n_18),
.B2(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_7),
.B1(n_18),
.B2(n_57),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_2),
.A2(n_26),
.B(n_57),
.C(n_164),
.Y(n_163)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_3),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_3),
.A2(n_153),
.B(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_4),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_17),
.B1(n_46),
.B2(n_47),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_4),
.A2(n_17),
.B1(n_72),
.B2(n_73),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_5),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_57),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_7),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_7),
.A2(n_24),
.B(n_25),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_7),
.B(n_33),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_10),
.B(n_73),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_SL g214 ( 
.A1(n_7),
.A2(n_47),
.B(n_48),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_8),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_8),
.A2(n_31),
.B1(n_72),
.B2(n_73),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_18),
.B(n_21),
.C(n_22),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_18),
.Y(n_21)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_70),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_10),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_10),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

BUFx3_ASAP7_75t_SL g47 ( 
.A(n_11),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_36),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_34),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_27),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_19),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_22),
.Y(n_19)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_22),
.A2(n_30),
.B(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_23),
.A2(n_45),
.B(n_48),
.C(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_23),
.B(n_48),
.Y(n_52)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_24),
.A2(n_49),
.B(n_57),
.C(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_28),
.B(n_38),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_32),
.A2(n_33),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_33),
.A2(n_55),
.B(n_60),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_75),
.B(n_275),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_39),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_39),
.B(n_273),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_53),
.CI(n_58),
.CON(n_39),
.SN(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_44),
.B1(n_50),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_43),
.B(n_101),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_44),
.A2(n_100),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_45),
.A2(n_51),
.B1(n_99),
.B2(n_101),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_45),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_45),
.B(n_57),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_47),
.A2(n_57),
.B(n_70),
.C(n_191),
.Y(n_190)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_101),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_57),
.B(n_86),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_57),
.B(n_71),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_65),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_106),
.C(n_111),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_59),
.A2(n_98),
.B1(n_133),
.B2(n_160),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_59),
.B(n_160),
.C(n_161),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_59),
.A2(n_111),
.B1(n_133),
.B2(n_171),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_65),
.B1(n_119),
.B2(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_63),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_64),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_65),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_74),
.Y(n_65)
);

INVxp33_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_68),
.B(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_68),
.A2(n_71),
.B1(n_74),
.B2(n_93),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_68),
.A2(n_71),
.B1(n_96),
.B2(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_72),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_72),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_73),
.B(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_272),
.B(n_274),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_128),
.A3(n_139),
.B1(n_270),
.B2(n_271),
.C(n_277),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_113),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_78),
.B(n_113),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_97),
.C(n_104),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_79),
.B(n_97),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_81),
.A2(n_82),
.B1(n_92),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_82),
.A2(n_89),
.B(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

INVxp33_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_84),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_85),
.A2(n_86),
.B1(n_154),
.B2(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_86),
.A2(n_108),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_92),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_95),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_103),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_102),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_98),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_98),
.B(n_176),
.C(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_98),
.A2(n_160),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_103),
.B(n_115),
.C(n_125),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_104),
.A2(n_105),
.B1(n_267),
.B2(n_268),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_106),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_107),
.A2(n_109),
.B1(n_206),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_107),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_109),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_109),
.B(n_165),
.C(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_109),
.A2(n_206),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_109),
.B(n_224),
.C(n_229),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_110),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_116),
.C(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_156),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_111),
.A2(n_146),
.B1(n_147),
.B2(n_171),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_111),
.B(n_147),
.C(n_212),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_114),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_124),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_116),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_124),
.B1(n_132),
.B2(n_137),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_116),
.A2(n_124),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_116),
.A2(n_124),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_116),
.B(n_245),
.C(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_124),
.B(n_137),
.C(n_138),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_129),
.B(n_130),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_138),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_264),
.B(n_269),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_252),
.B(n_263),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_181),
.B(n_237),
.C(n_251),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_167),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_143),
.B(n_167),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_158),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_145),
.B(n_155),
.C(n_158),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_147),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_146),
.B(n_151),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_147),
.B(n_190),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_154),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_165),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

NOR2x1_ASAP7_75t_R g196 ( 
.A(n_165),
.B(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_197),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_165),
.A2(n_174),
.B1(n_203),
.B2(n_207),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_166),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.C(n_175),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_168),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_173),
.B(n_175),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_188),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_236),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_231),
.B(n_235),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_221),
.B(n_230),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_209),
.B(n_220),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_200),
.B(n_208),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_192),
.B(n_199),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_196),
.B(n_198),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_215),
.B(n_218),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_228),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_232),
.B(n_233),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_239),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_249),
.B2(n_250),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_242),
.B(n_244),
.C(n_250),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_249),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_262),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_256),
.B(n_260),
.C(n_262),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_266),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);


endmodule