module fake_jpeg_4819_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_3),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_41),
.B(n_47),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_52),
.Y(n_74)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_15),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_55),
.B1(n_29),
.B2(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_56),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_19),
.B(n_8),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_57),
.B(n_58),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_8),
.Y(n_60)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_62),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_28),
.B(n_1),
.C(n_2),
.Y(n_62)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_21),
.B1(n_39),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_67),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_34),
.B1(n_29),
.B2(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_68),
.A2(n_90),
.B1(n_94),
.B2(n_100),
.Y(n_132)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_70),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_41),
.A2(n_26),
.B1(n_21),
.B2(n_34),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_71),
.B(n_73),
.Y(n_115)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_36),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_76),
.B(n_78),
.Y(n_131)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_79),
.B(n_83),
.Y(n_133)
);

AOI21xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_30),
.B(n_33),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_80),
.A2(n_4),
.B(n_11),
.Y(n_127)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_86),
.Y(n_136)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_29),
.B1(n_28),
.B2(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_48),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_43),
.A2(n_31),
.B1(n_50),
.B2(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_46),
.A2(n_32),
.B1(n_37),
.B2(n_20),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_92),
.B(n_93),
.Y(n_138)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_62),
.A2(n_37),
.B1(n_33),
.B2(n_30),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_33),
.B1(n_22),
.B2(n_17),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_42),
.A2(n_18),
.B1(n_22),
.B2(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_10),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_4),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_112),
.Y(n_114)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_55),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_106),
.B(n_110),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_51),
.A2(n_9),
.B1(n_13),
.B2(n_5),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_108),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_10),
.B1(n_12),
.B2(n_7),
.Y(n_109)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_7),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_51),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_112)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_122),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_3),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_123),
.B(n_87),
.Y(n_170)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_125),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_127),
.A2(n_126),
.B(n_114),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_81),
.B(n_14),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_137),
.Y(n_179)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_95),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_141),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_72),
.B(n_68),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_85),
.Y(n_155)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_95),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_143),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_69),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_97),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_148),
.Y(n_206)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_150),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_121),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_153),
.Y(n_193)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_140),
.A2(n_72),
.B1(n_70),
.B2(n_96),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_154),
.A2(n_155),
.B1(n_159),
.B2(n_177),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_179),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_107),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_156),
.B(n_162),
.Y(n_191)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_103),
.B(n_76),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_159),
.A2(n_115),
.B(n_137),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_116),
.A2(n_98),
.B1(n_82),
.B2(n_99),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_167),
.B1(n_175),
.B2(n_66),
.Y(n_198)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_163),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_120),
.B(n_128),
.Y(n_189)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_166),
.B(n_172),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_132),
.A2(n_113),
.B1(n_114),
.B2(n_127),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_87),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_174),
.B(n_130),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_132),
.A2(n_92),
.B1(n_111),
.B2(n_66),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_125),
.B(n_65),
.Y(n_177)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_178),
.Y(n_181)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_188),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_187),
.B(n_157),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_165),
.A2(n_167),
.B(n_173),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_203),
.B(n_211),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_212),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_170),
.A2(n_119),
.B(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_187),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_194),
.A2(n_204),
.B1(n_161),
.B2(n_176),
.Y(n_223)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_78),
.C(n_86),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_198),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_205),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_207),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_105),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_162),
.A2(n_73),
.B1(n_79),
.B2(n_111),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_104),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_149),
.B(n_143),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_210),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_151),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_209),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_166),
.B(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_180),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_180),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_150),
.B(n_153),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_218),
.B(n_222),
.Y(n_245)
);

NAND2xp33_ASAP7_75t_SL g218 ( 
.A(n_189),
.B(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_230),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_223),
.A2(n_229),
.B1(n_181),
.B2(n_183),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_152),
.B1(n_186),
.B2(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_203),
.B1(n_184),
.B2(n_191),
.Y(n_243)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_203),
.Y(n_242)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_234),
.Y(n_241)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_235),
.B(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_209),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_186),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_224),
.Y(n_271)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_239),
.B(n_231),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_257),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_215),
.Y(n_246)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_246),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_201),
.B1(n_188),
.B2(n_181),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_247),
.A2(n_253),
.B1(n_256),
.B2(n_226),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_250),
.Y(n_275)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_182),
.B1(n_190),
.B2(n_212),
.Y(n_251)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_206),
.B1(n_213),
.B2(n_199),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_255),
.B(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_218),
.A2(n_196),
.B1(n_199),
.B2(n_225),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_199),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_223),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_235),
.B(n_229),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_252),
.B(n_245),
.Y(n_276)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_241),
.B(n_216),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_255),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_238),
.C(n_221),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_267),
.C(n_252),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_221),
.C(n_222),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_268),
.A2(n_249),
.B(n_255),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_240),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_270),
.B(n_247),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_251),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_273),
.B1(n_242),
.B2(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_259),
.A2(n_224),
.B1(n_220),
.B2(n_219),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_237),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_280),
.B(n_283),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_286),
.C(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_242),
.B(n_245),
.C(n_243),
.D(n_256),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_261),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_272),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_270),
.B(n_233),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_282),
.B(n_288),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_268),
.A2(n_226),
.B(n_253),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_266),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_240),
.C(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_274),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_264),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_293),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_291),
.B(n_295),
.Y(n_309)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_267),
.C(n_271),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_292),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_280),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_261),
.C(n_264),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_296),
.B(n_300),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_303),
.A2(n_306),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_254),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_304),
.B(n_284),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_297),
.A2(n_283),
.B1(n_269),
.B2(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_295),
.B1(n_301),
.B2(n_269),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_250),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_312),
.B(n_313),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_299),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_254),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_314),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_294),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_286),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_293),
.C(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_317),
.A2(n_314),
.B(n_311),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_321),
.Y(n_322)
);

O2A1O1Ixp33_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_306),
.B(n_320),
.C(n_230),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_302),
.B(n_246),
.Y(n_324)
);


endmodule