module fake_jpeg_16340_n_359 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_359);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_359;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_34),
.B(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_33),
.Y(n_72)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_32),
.B1(n_35),
.B2(n_19),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_59),
.A2(n_71),
.B1(n_47),
.B2(n_29),
.Y(n_107)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_32),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_78),
.Y(n_84)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_39),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_SL g76 ( 
.A(n_46),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_54),
.C(n_49),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_0),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_89),
.B(n_38),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_47),
.B1(n_46),
.B2(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_98),
.B1(n_101),
.B2(n_64),
.Y(n_113)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_24),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_92),
.B(n_87),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_94),
.Y(n_121)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_65),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_103),
.Y(n_135)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_66),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_55),
.B1(n_40),
.B2(n_41),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_67),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_49),
.B1(n_24),
.B2(n_37),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_107),
.A2(n_64),
.B1(n_66),
.B2(n_77),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_125),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_113),
.A2(n_44),
.B1(n_55),
.B2(n_58),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_83),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_84),
.A2(n_54),
.B1(n_40),
.B2(n_41),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_74),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_128),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_88),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_100),
.A2(n_39),
.B1(n_34),
.B2(n_30),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_123),
.A2(n_124),
.B1(n_20),
.B2(n_18),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_30),
.B1(n_38),
.B2(n_62),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_101),
.A2(n_54),
.B1(n_41),
.B2(n_44),
.Y(n_125)
);

XNOR2x1_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_82),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_74),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_60),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_138),
.B(n_109),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_140),
.B(n_26),
.Y(n_142)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_81),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_166),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_112),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_148),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_158),
.B(n_160),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_132),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_45),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_48),
.C(n_28),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_55),
.B1(n_44),
.B2(n_27),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_157),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_140),
.B(n_31),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_126),
.B(n_31),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_165),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_164),
.B(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_113),
.B(n_114),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_93),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_60),
.B1(n_80),
.B2(n_11),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_97),
.B1(n_85),
.B2(n_108),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_168),
.A2(n_131),
.B1(n_133),
.B2(n_116),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_135),
.B(n_31),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_115),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_175),
.Y(n_211)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_142),
.B(n_137),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_147),
.A2(n_143),
.B(n_150),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_176),
.A2(n_188),
.B1(n_191),
.B2(n_48),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_127),
.B(n_121),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_178),
.A2(n_195),
.B(n_0),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_149),
.B(n_130),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_179),
.B(n_183),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_130),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_143),
.B(n_133),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_131),
.B1(n_116),
.B2(n_20),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_45),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_190),
.B(n_193),
.C(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_136),
.B1(n_109),
.B2(n_108),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_31),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_146),
.A2(n_120),
.B1(n_28),
.B2(n_18),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_167),
.B1(n_160),
.B2(n_144),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_162),
.A2(n_120),
.B(n_22),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_28),
.Y(n_198)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_146),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_199),
.A2(n_217),
.B(n_220),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_200),
.A2(n_203),
.B1(n_204),
.B2(n_212),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_156),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_202),
.C(n_208),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_189),
.A2(n_150),
.B1(n_145),
.B2(n_166),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_145),
.B1(n_164),
.B2(n_148),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_213),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_196),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_182),
.A2(n_129),
.B1(n_112),
.B2(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_214),
.A2(n_215),
.B1(n_227),
.B2(n_198),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_129),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_45),
.C(n_28),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_226),
.C(n_197),
.Y(n_240)
);

AOI221xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.C(n_23),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_185),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_190),
.B(n_45),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_181),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_233),
.C(n_239),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_226),
.B(n_173),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_245),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_193),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_36),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_193),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_242),
.C(n_243),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_181),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_186),
.C(n_184),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_216),
.C(n_222),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_249),
.C(n_252),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_170),
.B1(n_191),
.B2(n_194),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_247),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_180),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_206),
.A2(n_187),
.B1(n_184),
.B2(n_175),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_250),
.A2(n_218),
.B1(n_222),
.B2(n_195),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_214),
.A2(n_187),
.B1(n_179),
.B2(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_195),
.Y(n_252)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_192),
.Y(n_255)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_216),
.B1(n_211),
.B2(n_200),
.Y(n_256)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_221),
.B1(n_172),
.B2(n_203),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_260),
.A2(n_266),
.B1(n_272),
.B2(n_249),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_270),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_172),
.CI(n_227),
.CON(n_262),
.SN(n_262)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_244),
.A2(n_18),
.B1(n_20),
.B2(n_23),
.Y(n_263)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

INVxp33_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_13),
.B(n_16),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_265),
.A2(n_16),
.B(n_15),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_243),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_248),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_45),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_280),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_232),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_14),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_276),
.B(n_235),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_22),
.Y(n_280)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_286),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_264),
.B(n_237),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_299),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_277),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_293),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_260),
.A2(n_252),
.B(n_238),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_292),
.A2(n_257),
.B(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_263),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_258),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_294),
.B(n_295),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_258),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_298),
.B1(n_266),
.B2(n_262),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_239),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_295),
.C(n_294),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_242),
.B1(n_240),
.B2(n_245),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_261),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_281),
.A2(n_278),
.B1(n_275),
.B2(n_269),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_301),
.A2(n_306),
.B1(n_314),
.B2(n_305),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_279),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_307),
.C(n_308),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_290),
.B(n_282),
.Y(n_303)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_303),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_283),
.A2(n_272),
.B(n_270),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_304),
.A2(n_23),
.B(n_26),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_273),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_285),
.A2(n_262),
.B(n_231),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_309),
.A2(n_15),
.B(n_9),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_312),
.B(n_313),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_271),
.C(n_280),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_285),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_306),
.A2(n_287),
.B(n_299),
.Y(n_316)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_316),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_289),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_317),
.B(n_320),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_300),
.B(n_291),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_287),
.B1(n_296),
.B2(n_7),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_321),
.B1(n_326),
.B2(n_328),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_309),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_325),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_301),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_313),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_331),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_307),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_337),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_320),
.A2(n_308),
.B1(n_302),
.B2(n_311),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_335),
.B(n_338),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_319),
.B(n_20),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_333),
.A2(n_327),
.B(n_325),
.Y(n_341)
);

OAI321xp33_ASAP7_75t_L g349 ( 
.A1(n_341),
.A2(n_334),
.A3(n_12),
.B1(n_14),
.B2(n_11),
.C(n_26),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_345),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_SL g343 ( 
.A(n_339),
.B(n_329),
.Y(n_343)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_343),
.A2(n_14),
.B(n_23),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_338),
.B(n_326),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_330),
.A2(n_321),
.B(n_317),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_346),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_334),
.C(n_336),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_348),
.B(n_349),
.Y(n_354)
);

NAND4xp25_ASAP7_75t_SL g353 ( 
.A(n_350),
.B(n_36),
.C(n_81),
.D(n_22),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_353),
.A2(n_340),
.B(n_351),
.Y(n_355)
);

BUFx24_ASAP7_75t_SL g356 ( 
.A(n_355),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_354),
.B(n_352),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_357),
.A2(n_344),
.B(n_36),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_358),
.A2(n_22),
.B(n_352),
.Y(n_359)
);


endmodule