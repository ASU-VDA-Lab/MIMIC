module fake_jpeg_22220_n_306 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_306);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_306;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_305;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_42),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_31),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_31),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_40),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_22),
.B1(n_38),
.B2(n_19),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_51),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_49),
.B1(n_43),
.B2(n_22),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_69),
.B1(n_28),
.B2(n_23),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_57),
.B(n_62),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_22),
.B1(n_30),
.B2(n_24),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_63),
.B1(n_75),
.B2(n_78),
.Y(n_106)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_30),
.B1(n_34),
.B2(n_26),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_24),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_69),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_26),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_49),
.A2(n_42),
.B1(n_45),
.B2(n_29),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_71),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g72 ( 
.A1(n_42),
.A2(n_36),
.B(n_35),
.C(n_32),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_76),
.B(n_36),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_26),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_49),
.A2(n_18),
.B1(n_21),
.B2(n_34),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_24),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_0),
.B(n_1),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_33),
.C(n_0),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_18),
.B1(n_21),
.B2(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_79),
.B(n_88),
.Y(n_145)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_82),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_32),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_32),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_90),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_86),
.A2(n_91),
.B1(n_102),
.B2(n_107),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_87),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_19),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_37),
.Y(n_89)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_28),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_29),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_79),
.C(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_37),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_53),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_96),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_108),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_103),
.B1(n_109),
.B2(n_70),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_68),
.B(n_14),
.Y(n_126)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_46),
.B1(n_44),
.B2(n_33),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_66),
.A2(n_52),
.B1(n_54),
.B2(n_70),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_13),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_77),
.A2(n_46),
.B1(n_44),
.B2(n_36),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_66),
.A2(n_70),
.B1(n_54),
.B2(n_58),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_50),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_115),
.B(n_83),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_66),
.A2(n_32),
.B1(n_36),
.B2(n_35),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_61),
.B(n_65),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_35),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_0),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_128),
.B1(n_132),
.B2(n_144),
.Y(n_157)
);

CKINVDCx9p33_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_118),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_55),
.B(n_73),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_129),
.B(n_137),
.Y(n_150)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_142),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_149),
.B(n_112),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_54),
.B1(n_50),
.B2(n_61),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_55),
.B(n_40),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_12),
.Y(n_131)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_133),
.C(n_134),
.Y(n_155)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_10),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g137 ( 
.A1(n_91),
.A2(n_40),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_86),
.Y(n_170)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_106),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_144)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_147),
.Y(n_158)
);

INVx13_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

CKINVDCx11_ASAP7_75t_R g151 ( 
.A(n_142),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_148),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_167),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_99),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_162),
.C(n_164),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_119),
.A2(n_82),
.B1(n_121),
.B2(n_133),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_135),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_159),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_122),
.A2(n_84),
.B(n_81),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_160),
.A2(n_174),
.B(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_168),
.B(n_170),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_120),
.B(n_80),
.C(n_102),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_100),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_80),
.C(n_104),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_119),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_123),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_98),
.B(n_94),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_88),
.B(n_104),
.Y(n_174)
);

AO22x1_ASAP7_75t_L g175 ( 
.A1(n_137),
.A2(n_88),
.B1(n_101),
.B2(n_116),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_92),
.Y(n_176)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_176),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_114),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_137),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_147),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_6),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_126),
.C(n_125),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_150),
.B(n_174),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_139),
.Y(n_189)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_127),
.B1(n_118),
.B2(n_143),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_190),
.A2(n_201),
.B1(n_208),
.B2(n_182),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_127),
.C(n_136),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_192),
.B(n_181),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_195),
.B(n_197),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_177),
.B(n_136),
.Y(n_196)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_159),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_143),
.B1(n_125),
.B2(n_141),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_141),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_9),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_124),
.Y(n_205)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_124),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_208),
.B(n_6),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_92),
.C(n_130),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_179),
.C(n_160),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_210),
.B(n_231),
.C(n_209),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_172),
.Y(n_211)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_211),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_212),
.B(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_227),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_223),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_194),
.A2(n_150),
.B(n_175),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_191),
.B(n_190),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_170),
.B1(n_157),
.B2(n_155),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_218),
.A2(n_220),
.B1(n_224),
.B2(n_226),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_207),
.A2(n_180),
.B1(n_166),
.B2(n_152),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_165),
.B(n_158),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_194),
.A2(n_165),
.B1(n_167),
.B2(n_178),
.Y(n_224)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_230),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_189),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_169),
.C(n_130),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_187),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_239),
.C(n_240),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_184),
.C(n_210),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_242),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_217),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_245),
.C(n_248),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_196),
.C(n_185),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_246),
.B(n_224),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_201),
.B1(n_202),
.B2(n_195),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_222),
.B1(n_214),
.B2(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_203),
.C(n_192),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_197),
.C(n_183),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_216),
.C(n_220),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_254),
.B(n_259),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_216),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_227),
.Y(n_257)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_215),
.B(n_223),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_260),
.A2(n_240),
.B(n_10),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_206),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_264),
.C(n_245),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_213),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_265),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_204),
.B1(n_229),
.B2(n_169),
.Y(n_265)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_249),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_266),
.B(n_9),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_269),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_239),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_271),
.B(n_272),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_248),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_276),
.A2(n_278),
.B(n_267),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_169),
.C(n_114),
.Y(n_278)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_263),
.A3(n_252),
.B1(n_266),
.B2(n_257),
.C1(n_265),
.C2(n_267),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_270),
.B(n_268),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_275),
.A2(n_262),
.B(n_260),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_281),
.A2(n_276),
.B(n_277),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_258),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_273),
.A2(n_256),
.B1(n_258),
.B2(n_252),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_271),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_288),
.A2(n_292),
.B1(n_280),
.B2(n_282),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_269),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_287),
.B(n_281),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_11),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_294),
.B(n_11),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_297),
.B(n_13),
.Y(n_300)
);

AOI322xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_284),
.A3(n_283),
.B1(n_294),
.B2(n_289),
.C1(n_16),
.C2(n_11),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_300),
.B1(n_297),
.B2(n_14),
.C(n_15),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_302),
.A2(n_303),
.B1(n_13),
.B2(n_15),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_301),
.B(n_298),
.C(n_15),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_16),
.C(n_17),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_298),
.Y(n_306)
);


endmodule