module fake_jpeg_12432_n_41 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_41);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_41;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_7),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_9),
.B(n_8),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_2),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_2),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_3),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_19),
.C(n_6),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_34),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_38),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_36),
.C(n_26),
.Y(n_41)
);


endmodule