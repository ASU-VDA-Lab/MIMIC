module fake_jpeg_17635_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_SL g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_46),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_47),
.Y(n_54)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_48),
.A2(n_16),
.B1(n_33),
.B2(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_21),
.B1(n_33),
.B2(n_16),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_50),
.A2(n_52),
.B1(n_59),
.B2(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_47),
.B1(n_39),
.B2(n_40),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_62),
.B1(n_32),
.B2(n_44),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_33),
.B1(n_27),
.B2(n_25),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_55),
.A2(n_57),
.B1(n_34),
.B2(n_22),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_32),
.B1(n_28),
.B2(n_26),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_32),
.B1(n_28),
.B2(n_23),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_19),
.B1(n_13),
.B2(n_15),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_34),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_91),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_44),
.B1(n_18),
.B2(n_24),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_70),
.A2(n_83),
.B1(n_90),
.B2(n_96),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_74),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_37),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_81),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_54),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_80),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_53),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_86),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_59),
.B1(n_65),
.B2(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_85),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_87),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_19),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_62),
.A2(n_38),
.B1(n_32),
.B2(n_48),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_64),
.B1(n_38),
.B2(n_63),
.Y(n_109)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_63),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_117),
.B1(n_119),
.B2(n_92),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_111),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_55),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_64),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_95),
.B1(n_91),
.B2(n_86),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_76),
.A2(n_52),
.B1(n_58),
.B2(n_42),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_63),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_122),
.B(n_111),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_82),
.B1(n_81),
.B2(n_72),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_131),
.B(n_141),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_58),
.B1(n_79),
.B2(n_78),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_110),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_76),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_136),
.C(n_139),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_89),
.B1(n_88),
.B2(n_93),
.Y(n_130)
);

FAx1_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_89),
.CI(n_69),
.CON(n_131),
.SN(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_89),
.B1(n_69),
.B2(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_96),
.B1(n_99),
.B2(n_87),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_107),
.B1(n_112),
.B2(n_119),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_138),
.B1(n_114),
.B2(n_121),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_75),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_142),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_37),
.C(n_56),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_103),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_144),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_56),
.C(n_35),
.Y(n_139)
);

HAxp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_35),
.CON(n_140),
.SN(n_140)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_123),
.B1(n_104),
.B2(n_118),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_98),
.B(n_42),
.C(n_58),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_56),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_109),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_29),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_145),
.B(n_105),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_125),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_147),
.A2(n_154),
.B1(n_165),
.B2(n_130),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_106),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_148),
.A2(n_153),
.B(n_158),
.Y(n_170)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_124),
.A3(n_101),
.B1(n_102),
.B2(n_100),
.C(n_105),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_157),
.B(n_159),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_146),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_104),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_104),
.Y(n_163)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_118),
.B(n_1),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_29),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_168),
.C(n_29),
.Y(n_183)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_56),
.C(n_35),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_115),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_0),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_173),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_134),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_183),
.C(n_186),
.Y(n_193)
);

OA21x2_ASAP7_75t_SL g175 ( 
.A1(n_157),
.A2(n_135),
.B(n_136),
.Y(n_175)
);

AOI321xp33_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_177),
.A3(n_189),
.B1(n_6),
.B2(n_14),
.C(n_13),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_154),
.B1(n_162),
.B2(n_158),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_131),
.B(n_141),
.C(n_132),
.D(n_133),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_138),
.B1(n_145),
.B2(n_139),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_178),
.A2(n_148),
.B1(n_9),
.B2(n_10),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_181),
.B(n_184),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_115),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_85),
.C(n_110),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_85),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_187),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_8),
.C(n_14),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_8),
.C(n_14),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_167),
.C(n_9),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_165),
.B1(n_164),
.B2(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_194),
.B1(n_197),
.B2(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_168),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_200),
.Y(n_212)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_148),
.A3(n_155),
.B1(n_151),
.B2(n_156),
.C1(n_160),
.C2(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_196),
.B(n_201),
.Y(n_214)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_182),
.Y(n_198)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_198),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_171),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_182),
.Y(n_203)
);

FAx1_ASAP7_75t_SL g211 ( 
.A(n_204),
.B(n_189),
.CI(n_177),
.CON(n_211),
.SN(n_211)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_185),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_205),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_206),
.B(n_190),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_186),
.C(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_208),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_178),
.C(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_187),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_216),
.Y(n_223)
);

FAx1_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_171),
.CI(n_180),
.CON(n_216),
.SN(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_181),
.C(n_179),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_220),
.B1(n_201),
.B2(n_192),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_179),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_218),
.B(n_5),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_5),
.B(n_11),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_230),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_217),
.A2(n_206),
.B(n_203),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_198),
.B1(n_202),
.B2(n_192),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_222),
.Y(n_237)
);

NAND4xp25_ASAP7_75t_SL g225 ( 
.A(n_209),
.B(n_202),
.C(n_197),
.D(n_2),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_226),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_209),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_215),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_232),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_208),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_231),
.A2(n_219),
.B(n_216),
.Y(n_233)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_230),
.B(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_237),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_241),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_207),
.C(n_212),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_213),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_248),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_SL g245 ( 
.A(n_234),
.B(n_216),
.C(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_232),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_238),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_223),
.Y(n_248)
);

OA22x2_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_223),
.B1(n_239),
.B2(n_210),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_243),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_228),
.C(n_212),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_211),
.C(n_7),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_7),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_249),
.C(n_250),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_258),
.B(n_251),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_244),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_15),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_261),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_211),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);


endmodule