module fake_jpeg_15475_n_77 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_24),
.A2(n_13),
.B(n_6),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_51),
.B(n_52),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_54),
.B(n_55),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_23),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_30),
.B(n_7),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_36),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_56),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.C(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_59),
.B(n_56),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_43),
.B2(n_45),
.Y(n_64)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_60),
.A2(n_24),
.B(n_29),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_44),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_47),
.B(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_25),
.C(n_26),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_70),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_42),
.B(n_47),
.Y(n_70)
);

NOR3xp33_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_27),
.C(n_39),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_37),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_71),
.B(n_28),
.Y(n_73)
);

AOI322xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_74),
.A3(n_22),
.B1(n_34),
.B2(n_42),
.C1(n_33),
.C2(n_41),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_33),
.C(n_46),
.Y(n_76)
);

AOI221xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_31),
.B1(n_50),
.B2(n_53),
.C(n_46),
.Y(n_77)
);


endmodule