module fake_jpeg_29182_n_123 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_123);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_123;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_53),
.C(n_40),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_57),
.A2(n_41),
.B1(n_53),
.B2(n_49),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_64),
.A2(n_54),
.B1(n_50),
.B2(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_49),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_51),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_41),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_42),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_62),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_87),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_14),
.B1(n_37),
.B2(n_34),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_68),
.B1(n_74),
.B2(n_65),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_6),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_13),
.B(n_33),
.C(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_15),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_6),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_73),
.A2(n_12),
.B1(n_29),
.B2(n_27),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_5),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_93),
.A2(n_102),
.B1(n_10),
.B2(n_76),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_96),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_97),
.B(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_5),
.Y(n_96)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_7),
.Y(n_100)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_7),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_104),
.B1(n_39),
.B2(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_8),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_79),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_23),
.B(n_24),
.C(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_108),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_17),
.B1(n_18),
.B2(n_21),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_112),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_99),
.Y(n_113)
);

NOR2xp67_ASAP7_75t_SL g118 ( 
.A(n_113),
.B(n_115),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_92),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_114),
.A2(n_103),
.B(n_110),
.Y(n_117)
);

OA21x2_ASAP7_75t_SL g119 ( 
.A1(n_117),
.A2(n_110),
.B(n_116),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_113),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_120),
.B(n_118),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_109),
.Y(n_122)
);

AOI221xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_111),
.B1(n_91),
.B2(n_106),
.C(n_90),
.Y(n_123)
);


endmodule