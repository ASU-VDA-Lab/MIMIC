module fake_jpeg_2205_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_241;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_13),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_49),
.B(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_25),
.B(n_1),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_35),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_60),
.B1(n_49),
.B2(n_54),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_63),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_72),
.Y(n_114)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_65),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_38),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_69),
.A2(n_12),
.B(n_10),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_21),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_40),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_75),
.A2(n_77),
.B1(n_79),
.B2(n_86),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_40),
.A2(n_35),
.B1(n_32),
.B2(n_31),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_27),
.B1(n_30),
.B2(n_28),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_83),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_29),
.B1(n_23),
.B2(n_22),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_94),
.B1(n_11),
.B2(n_78),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_20),
.B1(n_18),
.B2(n_16),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_88),
.B(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_39),
.B(n_20),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_39),
.B(n_18),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_39),
.A2(n_57),
.B1(n_51),
.B2(n_41),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_19),
.C(n_4),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_19),
.C(n_5),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_44),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_7),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_2),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_4),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_109),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_120),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_72),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_6),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_6),
.Y(n_124)
);

OR2x4_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_19),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_107),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_131),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_8),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_67),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_10),
.B(n_11),
.C(n_96),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_136),
.A2(n_137),
.B(n_78),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_144),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_101),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_143),
.B(n_149),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_62),
.A3(n_68),
.B1(n_89),
.B2(n_70),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_68),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_73),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_69),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_155),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_103),
.B1(n_66),
.B2(n_97),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_153),
.A2(n_159),
.B(n_136),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_129),
.A2(n_76),
.B1(n_100),
.B2(n_66),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_154),
.A2(n_119),
.B1(n_127),
.B2(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_111),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_156),
.B(n_157),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_110),
.B(n_84),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_123),
.B(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_163),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_162),
.Y(n_184)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_116),
.B(n_67),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_99),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_129),
.A2(n_76),
.B1(n_84),
.B2(n_104),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_164),
.A2(n_165),
.B1(n_113),
.B2(n_130),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_112),
.A2(n_104),
.B1(n_103),
.B2(n_74),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_167),
.B(n_118),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_171),
.B1(n_175),
.B2(n_153),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_115),
.B1(n_126),
.B2(n_121),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_120),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_115),
.B1(n_121),
.B2(n_133),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_176),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_138),
.B1(n_161),
.B2(n_142),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_156),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_183),
.B(n_189),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_164),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_140),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_144),
.B(n_117),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_141),
.Y(n_202)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_159),
.B(n_147),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_205),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_195),
.B1(n_201),
.B2(n_190),
.Y(n_214)
);

AOI221xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_159),
.B1(n_141),
.B2(n_157),
.C(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_146),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_198),
.B(n_204),
.Y(n_216)
);

OAI21x1_ASAP7_75t_L g224 ( 
.A1(n_202),
.A2(n_210),
.B(n_173),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_146),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_153),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_206),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_150),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_166),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_150),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_210),
.A2(n_188),
.A3(n_182),
.B1(n_187),
.B2(n_172),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_181),
.B(n_178),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_223),
.B(n_205),
.C(n_201),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_185),
.B1(n_184),
.B2(n_182),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_170),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_171),
.B(n_172),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_224),
.B(n_198),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_180),
.C(n_187),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_225),
.B(n_203),
.C(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_235),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_234),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_237),
.B(n_221),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_199),
.B1(n_207),
.B2(n_206),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_204),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_223),
.C(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_246),
.C(n_237),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_236),
.A2(n_222),
.B1(n_226),
.B2(n_199),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_228),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_216),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_233),
.Y(n_248)
);

AO21x2_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_217),
.B(n_221),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_244),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_250),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_245),
.B1(n_220),
.B2(n_219),
.Y(n_258)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_216),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_241),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_246),
.C(n_244),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g257 ( 
.A1(n_249),
.A2(n_244),
.A3(n_245),
.B1(n_231),
.B2(n_232),
.C1(n_219),
.C2(n_220),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_253),
.A2(n_244),
.B1(n_231),
.B2(n_211),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_169),
.C(n_174),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_254),
.A2(n_253),
.B(n_209),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_262),
.A2(n_263),
.B1(n_256),
.B2(n_259),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_264),
.B(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_260),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_261),
.B(n_168),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_149),
.C(n_168),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_145),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_268),
.Y(n_270)
);


endmodule