module real_jpeg_2955_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_139;
wire n_33;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_64),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_64),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_35),
.B1(n_63),
.B2(n_65),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_4),
.A2(n_35),
.B1(n_59),
.B2(n_61),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_9),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_9),
.A2(n_39),
.B1(n_59),
.B2(n_61),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_57),
.C(n_59),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_9),
.A2(n_23),
.B1(n_24),
.B2(n_39),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_9),
.A2(n_39),
.B1(n_63),
.B2(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_9),
.B(n_55),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_9),
.B(n_40),
.C(n_73),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_24),
.C(n_46),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_71),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_9),
.B(n_31),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_9),
.B(n_51),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_134),
.B1(n_252),
.B2(n_253),
.Y(n_13)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_133),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_108),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_17),
.B(n_108),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_81),
.C(n_99),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_18),
.A2(n_19),
.B1(n_99),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_52),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_20),
.B(n_70),
.C(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_21),
.B(n_36),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_32),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_22),
.A2(n_30),
.B(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_23),
.A2(n_24),
.B1(n_45),
.B2(n_46),
.Y(n_48)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_24),
.B(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_34),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_29),
.A2(n_30),
.B(n_107),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_29),
.B(n_107),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_29),
.B(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_30),
.B(n_216),
.Y(n_230)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_31),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_32),
.B(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_33),
.B(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_49),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_37),
.B(n_201),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_43),
.Y(n_37)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_38),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_38),
.B(n_51),
.Y(n_187)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_40),
.A2(n_42),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_40),
.B(n_210),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_43),
.B(n_50),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_43),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_43),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI21x1_ASAP7_75t_R g130 ( 
.A1(n_49),
.A2(n_102),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_49),
.B(n_188),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_51),
.B(n_189),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_70),
.B1(n_79),
.B2(n_80),
.Y(n_52)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_66),
.Y(n_53)
);

INVxp33_ASAP7_75t_L g146 ( 
.A(n_54),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_62),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_55),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_57),
.B1(n_63),
.B2(n_65),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_61),
.B1(n_73),
.B2(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_59),
.B(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_67),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_78),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_78),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_92),
.Y(n_155)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_73),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_75),
.B(n_78),
.Y(n_125)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_76),
.B(n_123),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_81),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_93),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_85),
.B(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_90),
.B(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_98),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B(n_103),
.Y(n_100)
);

AOI21x1_ASAP7_75t_SL g150 ( 
.A1(n_101),
.A2(n_131),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_103),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_105),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_126),
.B2(n_127),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_124),
.Y(n_121)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_132),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_128),
.A2(n_129),
.B1(n_182),
.B2(n_183),
.Y(n_203)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_130),
.Y(n_132)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_134),
.Y(n_253)
);

OAI21x1_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_156),
.B(n_249),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_136),
.A2(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_137),
.B(n_140),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.C(n_144),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_144),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_174),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_158),
.B(n_160),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_161),
.A2(n_162),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.C(n_170),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_173),
.B(n_230),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_193),
.B(n_248),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_190),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_185),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_177),
.A2(n_178),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_181),
.A2(n_185),
.B1(n_186),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21x1_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_204),
.B(n_247),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_199),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_202),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_203),
.B(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_242),
.B(n_246),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_224),
.B(n_241),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_208),
.A2(n_209),
.B1(n_211),
.B2(n_227),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_212)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_219),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_221),
.C(n_223),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_231),
.B(n_240),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_228),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_236),
.B(n_239),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_243),
.B(n_244),
.Y(n_246)
);


endmodule