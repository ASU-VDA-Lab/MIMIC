module fake_jpeg_10568_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

HAxp5_ASAP7_75t_SL g65 ( 
.A(n_39),
.B(n_30),
.CON(n_65),
.SN(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_1),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_17),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_52),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_48),
.A2(n_65),
.B1(n_32),
.B2(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_36),
.B2(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_61),
.B1(n_63),
.B2(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_23),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_57),
.B(n_64),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_37),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_23),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_20),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_32),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_22),
.B(n_21),
.C(n_16),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_32),
.B1(n_22),
.B2(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_40),
.B(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_69),
.Y(n_89)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_82),
.Y(n_105)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_75),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_71),
.A2(n_76),
.B1(n_16),
.B2(n_27),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_77),
.A2(n_79),
.B1(n_84),
.B2(n_58),
.Y(n_86)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_19),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_63),
.A2(n_19),
.B1(n_20),
.B2(n_17),
.Y(n_84)
);

HAxp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_49),
.CON(n_85),
.SN(n_85)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_102),
.B(n_45),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_67),
.B1(n_51),
.B2(n_19),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_92),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_74),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_52),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_99),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_46),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_84),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_60),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_62),
.Y(n_102)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_62),
.B(n_59),
.Y(n_106)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_111),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_77),
.B1(n_78),
.B2(n_81),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_107),
.A2(n_112),
.B1(n_118),
.B2(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_50),
.B1(n_62),
.B2(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_102),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_24),
.A3(n_31),
.B1(n_28),
.B2(n_34),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g129 ( 
.A1(n_115),
.A2(n_101),
.B(n_94),
.C(n_102),
.D(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_34),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_121),
.C(n_108),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_104),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_124),
.C(n_114),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_134),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_141),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_112),
.A2(n_95),
.B(n_87),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_106),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_133),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_136),
.B1(n_112),
.B2(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_138),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_88),
.B1(n_98),
.B2(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_88),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_140),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_107),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_142),
.A2(n_143),
.B1(n_108),
.B2(n_116),
.Y(n_144)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_90),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_129),
.B(n_141),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_147),
.A2(n_148),
.B(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_128),
.A2(n_126),
.B(n_135),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_155),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_151),
.C(n_154),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_131),
.C(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_123),
.C(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_143),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_157),
.B(n_132),
.C(n_140),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_119),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_168),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_162),
.A2(n_164),
.B(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_163),
.B(n_165),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_158),
.A2(n_17),
.B(n_27),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_159),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_170),
.B(n_146),
.Y(n_181)
);

AOI21x1_ASAP7_75t_SL g171 ( 
.A1(n_148),
.A2(n_24),
.B(n_31),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_171),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_151),
.B(n_147),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_178),
.A2(n_181),
.B1(n_160),
.B2(n_28),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_180),
.Y(n_188)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_149),
.B1(n_169),
.B2(n_152),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_161),
.C(n_157),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_187),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_189),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_160),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_24),
.A3(n_14),
.B1(n_12),
.B2(n_11),
.C1(n_10),
.C2(n_6),
.Y(n_190)
);

AOI322xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_183),
.A3(n_185),
.B1(n_12),
.B2(n_189),
.C1(n_5),
.C2(n_1),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_173),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_195),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_176),
.B(n_179),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_1),
.B(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_11),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_3),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_197),
.A2(n_198),
.B1(n_193),
.B2(n_7),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_191),
.A2(n_4),
.B(n_5),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_201),
.B(n_7),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_200),
.A2(n_4),
.B(n_8),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_204),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_199),
.B(n_8),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_206),
.Y(n_208)
);


endmodule