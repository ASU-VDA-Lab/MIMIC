module fake_jpeg_29133_n_101 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_101);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_101;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_6),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_1),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx6p67_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g38 ( 
.A1(n_14),
.A2(n_3),
.B(n_7),
.C(n_8),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_9),
.Y(n_42)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_50),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_28),
.A2(n_19),
.B1(n_12),
.B2(n_20),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_17),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_57),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_29),
.B1(n_19),
.B2(n_16),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_54),
.A2(n_21),
.B1(n_23),
.B2(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_16),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_21),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_65),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_20),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_64),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_52),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_47),
.C(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_68),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_69),
.B(n_72),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_48),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_63),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_79),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_48),
.B(n_43),
.C(n_47),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_82),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_78),
.A2(n_61),
.B(n_60),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_45),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_81),
.B1(n_77),
.B2(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_89),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_90),
.A2(n_83),
.B(n_84),
.Y(n_95)
);

AO221x1_ASAP7_75t_L g91 ( 
.A1(n_85),
.A2(n_73),
.B1(n_82),
.B2(n_79),
.C(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_96),
.B1(n_93),
.B2(n_92),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_87),
.B1(n_84),
.B2(n_88),
.Y(n_96)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_94),
.B(n_96),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_49),
.B(n_55),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_45),
.C(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_100),
.Y(n_101)
);


endmodule