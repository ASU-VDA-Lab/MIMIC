module fake_jpeg_1204_n_450 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_450);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_450;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_58),
.B(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_38),
.A2(n_1),
.B(n_2),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g173 ( 
.A(n_62),
.B(n_2),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_67),
.Y(n_122)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_66),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_7),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_68),
.B(n_69),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_70),
.Y(n_115)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_71),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_20),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_72),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_21),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_74),
.B(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_75),
.Y(n_180)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_78),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_36),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_83),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_41),
.B(n_1),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_84),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_87),
.Y(n_163)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_88),
.B(n_90),
.Y(n_144)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_92),
.B(n_98),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_24),
.B(n_15),
.Y(n_98)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_14),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_107),
.Y(n_174)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_37),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_111),
.Y(n_161)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_108),
.Y(n_147)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_40),
.B(n_1),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_27),
.B(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_109),
.B(n_110),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_47),
.B(n_10),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_34),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_112),
.B(n_22),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_34),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_102),
.A2(n_31),
.B1(n_50),
.B2(n_54),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_117),
.A2(n_120),
.B1(n_126),
.B2(n_138),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_62),
.A2(n_31),
.B1(n_50),
.B2(n_29),
.Y(n_119)
);

AOI22x1_ASAP7_75t_L g221 ( 
.A1(n_119),
.A2(n_160),
.B1(n_172),
.B2(n_151),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_56),
.A2(n_54),
.B1(n_29),
.B2(n_28),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_56),
.A2(n_54),
.B1(n_44),
.B2(n_52),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_68),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_128),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_134),
.B(n_124),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_82),
.A2(n_77),
.B1(n_86),
.B2(n_59),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_136),
.A2(n_154),
.B1(n_156),
.B2(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_44),
.B1(n_52),
.B2(n_48),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_153),
.B1(n_4),
.B2(n_140),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_66),
.A2(n_76),
.B1(n_96),
.B2(n_73),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_108),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_100),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_106),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_104),
.A2(n_48),
.B1(n_42),
.B2(n_35),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_149),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_173),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_65),
.A2(n_53),
.B1(n_42),
.B2(n_35),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_94),
.A2(n_95),
.B1(n_103),
.B2(n_89),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_91),
.A2(n_99),
.B1(n_97),
.B2(n_57),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_180),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_78),
.A2(n_34),
.B1(n_39),
.B2(n_26),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_79),
.A2(n_93),
.B1(n_84),
.B2(n_71),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_113),
.A2(n_34),
.B1(n_53),
.B2(n_39),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_176),
.B1(n_177),
.B2(n_182),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_93),
.A2(n_53),
.B1(n_26),
.B2(n_9),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_70),
.A2(n_53),
.B1(n_25),
.B2(n_5),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_87),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_87),
.A2(n_4),
.B1(n_6),
.B2(n_105),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_183),
.A2(n_115),
.B1(n_163),
.B2(n_133),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_185),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_153),
.B1(n_127),
.B2(n_121),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_186),
.A2(n_218),
.B1(n_215),
.B2(n_225),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_187),
.A2(n_224),
.B1(n_188),
.B2(n_211),
.Y(n_259)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_188),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_190),
.B(n_193),
.Y(n_249)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_192),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_114),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_4),
.C(n_174),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_194),
.B(n_196),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_158),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_123),
.B(n_122),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_197),
.B(n_198),
.Y(n_254)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_179),
.B(n_181),
.C(n_137),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g261 ( 
.A1(n_199),
.A2(n_221),
.B1(n_189),
.B2(n_219),
.Y(n_261)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g274 ( 
.A(n_200),
.Y(n_274)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_129),
.Y(n_201)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_201),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_131),
.B(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_206),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_148),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_116),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_208),
.B(n_210),
.Y(n_272)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_181),
.Y(n_209)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_211),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_121),
.B(n_164),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_116),
.B(n_145),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_213),
.B(n_228),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_133),
.Y(n_214)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_145),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_215),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_216),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_127),
.B(n_164),
.C(n_147),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_222),
.C(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_136),
.B(n_129),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_225),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_152),
.C(n_151),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_223),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_226),
.B(n_227),
.Y(n_282)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_130),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_166),
.B(n_130),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_229),
.B(n_230),
.Y(n_276)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_125),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_152),
.B(n_150),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_232),
.B(n_233),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_150),
.B(n_125),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_132),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_171),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_135),
.Y(n_238)
);

CKINVDCx11_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_141),
.B(n_155),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_141),
.A2(n_115),
.B1(n_159),
.B2(n_155),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_159),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_133),
.Y(n_242)
);

INVx13_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_SL g243 ( 
.A(n_207),
.B(n_205),
.C(n_184),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_263),
.C(n_277),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_240),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_207),
.Y(n_247)
);

A2O1A1O1Ixp25_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_236),
.B(n_235),
.C(n_234),
.D(n_230),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_259),
.A2(n_269),
.B1(n_192),
.B2(n_195),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_261),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_222),
.C(n_212),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_239),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_199),
.B(n_187),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_202),
.B(n_226),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_284),
.Y(n_305)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_215),
.B(n_241),
.Y(n_277)
);

OR2x2_ASAP7_75t_SL g280 ( 
.A(n_219),
.B(n_200),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_L g308 ( 
.A(n_280),
.B(n_231),
.C(n_216),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_201),
.B(n_227),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_284),
.Y(n_288)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_242),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_289),
.B(n_294),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_246),
.B(n_204),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_296),
.C(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_292),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_255),
.Y(n_293)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_293),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_250),
.B(n_214),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_260),
.Y(n_295)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_295),
.Y(n_340)
);

BUFx8_ASAP7_75t_L g297 ( 
.A(n_262),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_297),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_298),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_303),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_249),
.B(n_185),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_255),
.Y(n_301)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_301),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_283),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_304),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_310),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_308),
.A2(n_316),
.B(n_317),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_265),
.A2(n_216),
.B1(n_223),
.B2(n_268),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_309),
.A2(n_313),
.B1(n_266),
.B2(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_287),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_312),
.Y(n_349)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_265),
.A2(n_259),
.B1(n_247),
.B2(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_315),
.B1(n_320),
.B2(n_321),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_277),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_318),
.A2(n_271),
.B(n_281),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_248),
.B(n_263),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_319),
.B(n_253),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_275),
.B(n_270),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_264),
.B(n_273),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_322),
.A2(n_298),
.B1(n_290),
.B2(n_305),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_248),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_346),
.C(n_291),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_307),
.A2(n_265),
.B(n_261),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_325),
.A2(n_327),
.B(n_317),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_307),
.A2(n_261),
.B(n_271),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_328),
.B(n_331),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_330),
.A2(n_339),
.B(n_297),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_290),
.A2(n_252),
.B1(n_251),
.B2(n_245),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_347),
.Y(n_362)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_313),
.A2(n_251),
.B(n_253),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g370 ( 
.A(n_336),
.B(n_293),
.C(n_318),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_309),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_302),
.B(n_266),
.C(n_245),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_288),
.A2(n_252),
.B1(n_256),
.B2(n_276),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_350),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_348),
.B(n_305),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_352),
.C(n_353),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_348),
.B(n_310),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_315),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_365),
.B(n_368),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_323),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_355),
.B(n_357),
.Y(n_389)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_356),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_323),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_358),
.B(n_364),
.C(n_346),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_333),
.B(n_301),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_359),
.B(n_367),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_360),
.A2(n_366),
.B1(n_370),
.B2(n_344),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_361),
.B(n_363),
.Y(n_380)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_342),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_SL g364 ( 
.A(n_331),
.B(n_302),
.C(n_296),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_299),
.B(n_316),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_344),
.B(n_293),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_341),
.B(n_321),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_371),
.A2(n_329),
.B1(n_347),
.B2(n_338),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_360),
.A2(n_343),
.B1(n_325),
.B2(n_336),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_372),
.A2(n_373),
.B1(n_379),
.B2(n_381),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_375),
.B(n_377),
.C(n_382),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_364),
.B(n_358),
.C(n_369),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_368),
.A2(n_343),
.B1(n_336),
.B2(n_339),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_343),
.B1(n_326),
.B2(n_334),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_324),
.C(n_328),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_383),
.A2(n_371),
.B(n_354),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_326),
.C(n_341),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_384),
.B(n_387),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_369),
.B(n_329),
.C(n_332),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_353),
.A2(n_352),
.B1(n_351),
.B2(n_359),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_340),
.C(n_335),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_267),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_390),
.B(n_350),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_384),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_393),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_365),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_378),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_394),
.B(n_398),
.Y(n_407)
);

BUFx12f_ASAP7_75t_SL g395 ( 
.A(n_376),
.Y(n_395)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_400),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_399),
.Y(n_417)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_385),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_389),
.A2(n_363),
.B1(n_356),
.B2(n_297),
.Y(n_399)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_386),
.B(n_370),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_402),
.B(n_366),
.Y(n_409)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_380),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_404),
.A2(n_367),
.B1(n_363),
.B2(n_381),
.Y(n_406)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_403),
.A2(n_374),
.B1(n_372),
.B2(n_379),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_408),
.A2(n_404),
.B1(n_391),
.B2(n_394),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_410),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_375),
.C(n_387),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_383),
.C(n_335),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_413),
.B(n_415),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_340),
.C(n_267),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_337),
.B1(n_244),
.B2(n_304),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_416),
.A2(n_412),
.B1(n_407),
.B2(n_413),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_412),
.A2(n_397),
.B(n_400),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_418),
.A2(n_411),
.B(n_410),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_419),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_414),
.A2(n_393),
.B1(n_395),
.B2(n_396),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_420),
.A2(n_424),
.B1(n_423),
.B2(n_417),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_408),
.A2(n_396),
.B1(n_337),
.B2(n_244),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_422),
.B(n_423),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_415),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_432),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_429),
.A2(n_430),
.B(n_431),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_418),
.A2(n_411),
.B(n_274),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_421),
.A2(n_285),
.B(n_257),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_283),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_279),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_433),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_427),
.A2(n_420),
.B(n_434),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_437),
.B(n_438),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_431),
.Y(n_438)
);

AOI21xp33_ASAP7_75t_SL g440 ( 
.A1(n_427),
.A2(n_422),
.B(n_425),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_440),
.A2(n_425),
.B(n_257),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_439),
.Y(n_441)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_441),
.A2(n_443),
.B(n_436),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_282),
.C(n_279),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_444),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_446),
.A2(n_442),
.B(n_262),
.Y(n_447)
);

NAND2xp33_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_448),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_445),
.A2(n_258),
.B(n_286),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_449),
.B(n_286),
.Y(n_450)
);


endmodule