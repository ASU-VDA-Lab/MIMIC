module fake_jpeg_7274_n_228 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_228);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_228;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_20),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx2_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_38),
.Y(n_50)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_40),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_16),
.B1(n_26),
.B2(n_18),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_26),
.B1(n_18),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_25),
.B1(n_18),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_16),
.B1(n_41),
.B2(n_36),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_15),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_16),
.B1(n_24),
.B2(n_23),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_55),
.Y(n_61)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_15),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_57),
.B1(n_34),
.B2(n_21),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_17),
.B1(n_27),
.B2(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_59),
.Y(n_65)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_33),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_62),
.A2(n_66),
.B(n_71),
.C(n_46),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_81),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_33),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_74),
.Y(n_88)
);

AND2x4_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_37),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_77),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_80),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g102 ( 
.A1(n_76),
.A2(n_60),
.B1(n_59),
.B2(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_58),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_79),
.A2(n_42),
.B1(n_48),
.B2(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_47),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_22),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_51),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_82),
.A2(n_49),
.B1(n_36),
.B2(n_46),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_91),
.B(n_62),
.Y(n_111)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_84),
.Y(n_108)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_13),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_87),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_90),
.B1(n_93),
.B2(n_102),
.Y(n_120)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_48),
.A3(n_39),
.B1(n_29),
.B2(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_39),
.B1(n_34),
.B2(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_92),
.B(n_95),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_82),
.A2(n_39),
.B1(n_31),
.B2(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_96),
.B(n_65),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_71),
.A2(n_46),
.B(n_35),
.C(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_74),
.B(n_13),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_68),
.B(n_13),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_79),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_38),
.B1(n_35),
.B2(n_40),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_66),
.B1(n_36),
.B2(n_59),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_71),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_107),
.A2(n_111),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_64),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_113),
.C(n_86),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_78),
.C(n_64),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_89),
.B(n_81),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_117),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_98),
.A2(n_69),
.B1(n_77),
.B2(n_62),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_100),
.B1(n_98),
.B2(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_65),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_93),
.B1(n_90),
.B2(n_127),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_60),
.Y(n_127)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_136),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_105),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_135),
.C(n_145),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_141),
.B(n_143),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_87),
.B(n_85),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_66),
.B(n_97),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_101),
.B1(n_97),
.B2(n_92),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_144),
.A2(n_147),
.B(n_126),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_54),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_55),
.C(n_36),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_106),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_0),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_151),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_116),
.Y(n_151)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_154),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_157),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_148),
.B(n_111),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_115),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_160),
.B(n_162),
.Y(n_176)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_109),
.C(n_117),
.D(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_122),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_121),
.C(n_124),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_108),
.B1(n_84),
.B2(n_139),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_164),
.A2(n_140),
.B1(n_143),
.B2(n_120),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_146),
.C(n_131),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_159),
.B(n_145),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_171),
.C(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_135),
.C(n_148),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_133),
.C(n_128),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_175),
.B(n_179),
.C(n_180),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_177),
.B(n_176),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_120),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_150),
.C(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_114),
.C(n_139),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_29),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_163),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_186),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_152),
.B1(n_165),
.B2(n_157),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_138),
.B(n_172),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_181),
.B(n_158),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_141),
.A3(n_115),
.B1(n_155),
.B2(n_152),
.C(n_122),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_171),
.B(n_167),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_173),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_153),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_138),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_189),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_184),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_203),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_29),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_197),
.B(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_84),
.C(n_27),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_199),
.C(n_191),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_27),
.C(n_28),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_192),
.Y(n_204)
);

BUFx24_ASAP7_75t_SL g203 ( 
.A(n_193),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_201),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_198),
.A2(n_192),
.B(n_190),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_208),
.B(n_210),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_191),
.B(n_8),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_9),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_214),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_204),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_202),
.B1(n_199),
.B2(n_2),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_205),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_215),
.A2(n_9),
.B(n_14),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_217),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_206),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g222 ( 
.A1(n_219),
.A2(n_220),
.A3(n_216),
.B1(n_215),
.B2(n_212),
.C1(n_4),
.C2(n_5),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_223),
.A3(n_7),
.B1(n_11),
.B2(n_5),
.C1(n_6),
.C2(n_12),
.Y(n_224)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_7),
.A3(n_12),
.B1(n_3),
.B2(n_5),
.C1(n_6),
.C2(n_14),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_224),
.A2(n_225),
.B(n_10),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_226),
.B(n_0),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_SL g228 ( 
.A(n_227),
.B(n_1),
.Y(n_228)
);


endmodule