module fake_jpeg_295_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_7),
.B(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_41),
.Y(n_101)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_46),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_44),
.B(n_50),
.Y(n_87)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_15),
.B(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_67),
.Y(n_108)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_3),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_57),
.B(n_63),
.Y(n_91)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_66),
.Y(n_92)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_18),
.B(n_3),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_36),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_68),
.B(n_69),
.Y(n_107)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

NOR2xp67_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_4),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_73),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_18),
.B(n_5),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_74),
.B(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_75),
.B(n_77),
.Y(n_105)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_38),
.Y(n_104)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_78),
.B(n_113),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_21),
.B1(n_37),
.B2(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_81),
.A2(n_103),
.B1(n_112),
.B2(n_8),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_19),
.B1(n_37),
.B2(n_29),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_86),
.A2(n_88),
.B1(n_117),
.B2(n_40),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_25),
.B1(n_34),
.B2(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_42),
.B(n_25),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_98),
.B(n_111),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_54),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_76),
.B(n_30),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g112 ( 
.A1(n_55),
.A2(n_38),
.B1(n_6),
.B2(n_7),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_59),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_69),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_71),
.A2(n_73),
.B1(n_56),
.B2(n_52),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_73),
.B1(n_53),
.B2(n_58),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_SL g164 ( 
.A1(n_118),
.A2(n_122),
.B(n_127),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_119),
.Y(n_155)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_107),
.A2(n_62),
.B1(n_61),
.B2(n_72),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_123),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_91),
.A2(n_108),
.B(n_99),
.C(n_90),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_139),
.B(n_145),
.Y(n_158)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_128),
.A2(n_134),
.B1(n_144),
.B2(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_131),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_137),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_92),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_136),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_40),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_101),
.A2(n_82),
.B1(n_114),
.B2(n_80),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_112),
.A2(n_101),
.B1(n_109),
.B2(n_116),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_134),
.Y(n_176)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_80),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_110),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_109),
.B1(n_83),
.B2(n_79),
.Y(n_144)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_85),
.B(n_110),
.C(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_149),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_85),
.A2(n_102),
.B1(n_93),
.B2(n_97),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_152),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_85),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g198 ( 
.A(n_157),
.Y(n_198)
);

FAx1_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_97),
.CI(n_121),
.CON(n_161),
.SN(n_161)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_161),
.A2(n_145),
.B(n_126),
.C(n_132),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_151),
.B(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_125),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_178),
.Y(n_187)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_130),
.B1(n_131),
.B2(n_119),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_139),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_120),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_165),
.Y(n_180)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_166),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_194),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_182),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_191),
.C(n_158),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_184),
.B(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_149),
.B1(n_150),
.B2(n_141),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_160),
.B(n_129),
.C(n_123),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_170),
.C(n_171),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_174),
.B1(n_173),
.B2(n_159),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_190),
.B(n_193),
.Y(n_199)
);

AO22x1_ASAP7_75t_L g190 ( 
.A1(n_161),
.A2(n_156),
.B1(n_172),
.B2(n_160),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_166),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_192),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_148),
.B(n_176),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_156),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_196),
.B(n_197),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_178),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_158),
.B(n_175),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_200),
.B(n_207),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_154),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_201),
.B(n_208),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_208),
.B(n_209),
.C(n_171),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_164),
.C(n_170),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_169),
.B(n_159),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_212),
.B1(n_196),
.B2(n_189),
.Y(n_223)
);

AOI322xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_187),
.A3(n_198),
.B1(n_182),
.B2(n_180),
.C1(n_179),
.C2(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_219),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_201),
.B(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_217),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_190),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_218),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_205),
.A2(n_188),
.B1(n_189),
.B2(n_186),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_205),
.B1(n_189),
.B2(n_199),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_209),
.B(n_194),
.Y(n_222)
);

AOI321xp33_ASAP7_75t_L g230 ( 
.A1(n_222),
.A2(n_213),
.A3(n_211),
.B1(n_203),
.B2(n_210),
.C(n_189),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_223),
.A2(n_224),
.B(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_228),
.A2(n_206),
.B1(n_212),
.B2(n_177),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_215),
.A2(n_199),
.B1(n_200),
.B2(n_213),
.Y(n_229)
);

A2O1A1Ixp33_ASAP7_75t_SL g236 ( 
.A1(n_229),
.A2(n_217),
.B(n_216),
.C(n_222),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_231),
.B(n_226),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_232),
.B(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_234),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_224),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_173),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_236),
.A2(n_225),
.B1(n_153),
.B2(n_177),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_206),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_174),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_238),
.A2(n_229),
.B1(n_230),
.B2(n_228),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_242),
.B(n_243),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_238),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_241),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_250),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_239),
.B(n_243),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_249),
.B(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_155),
.C(n_153),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_253),
.A2(n_251),
.B(n_245),
.Y(n_254)
);


endmodule