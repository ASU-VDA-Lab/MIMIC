module fake_jpeg_39_n_220 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_220);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_220;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_50),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_3),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_1),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_0),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_84),
.B(n_60),
.Y(n_98)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_58),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_95),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_59),
.B1(n_67),
.B2(n_74),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_74),
.B1(n_62),
.B2(n_68),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_89),
.A2(n_83),
.B1(n_81),
.B2(n_85),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g92 ( 
.A(n_80),
.B(n_73),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_66),
.B1(n_82),
.B2(n_24),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_106),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_65),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_85),
.B1(n_62),
.B2(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_110),
.A2(n_115),
.B1(n_70),
.B2(n_57),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_53),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_116),
.Y(n_133)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_99),
.Y(n_112)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_112),
.Y(n_126)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_63),
.B1(n_57),
.B2(n_71),
.Y(n_115)
);

FAx1_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_83),
.CI(n_81),
.CON(n_116),
.SN(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_22),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_121),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_56),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_123),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_54),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_128),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_64),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_130),
.B(n_134),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_90),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_108),
.A2(n_96),
.B1(n_71),
.B2(n_70),
.Y(n_135)
);

AO22x1_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_19),
.B1(n_41),
.B2(n_38),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_52),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_2),
.Y(n_146)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_25),
.B1(n_46),
.B2(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_140),
.B(n_18),
.Y(n_162)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_145),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_2),
.B(n_3),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_146),
.A2(n_157),
.B1(n_8),
.B2(n_12),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_149),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_21),
.C(n_44),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_27),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_123),
.A2(n_139),
.B1(n_134),
.B2(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_4),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_28),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_153),
.Y(n_173)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_136),
.Y(n_154)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_124),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_5),
.C(n_6),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_183),
.B1(n_13),
.B2(n_14),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_147),
.Y(n_170)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_148),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_144),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_178),
.A2(n_179),
.B(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_195),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_181),
.B(n_160),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_187),
.B(n_194),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_191),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_181),
.A2(n_151),
.B(n_158),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_30),
.C(n_35),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_196),
.B(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_180),
.B1(n_177),
.B2(n_172),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_197),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_180),
.B1(n_193),
.B2(n_187),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_176),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_173),
.C(n_165),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_173),
.B(n_184),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_174),
.B(n_171),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_206),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_194),
.C(n_15),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_201),
.C(n_198),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_182),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_199),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_211),
.B(n_212),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_210),
.A2(n_204),
.B1(n_208),
.B2(n_14),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_16),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_215),
.Y(n_216)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_214),
.B(n_26),
.C(n_32),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_17),
.C(n_33),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_51),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_219),
.B(n_34),
.Y(n_220)
);


endmodule