module real_jpeg_29156_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_4),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_61),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_7),
.A2(n_28),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_20),
.B1(n_22),
.B2(n_28),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_7),
.A2(n_28),
.B1(n_81),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_9),
.A2(n_31),
.B1(n_45),
.B2(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_20),
.B1(n_22),
.B2(n_31),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_20),
.B(n_70),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_9),
.A2(n_25),
.B(n_38),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_9),
.A2(n_31),
.B1(n_81),
.B2(n_88),
.Y(n_90)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_9),
.A2(n_46),
.B(n_60),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_9),
.B(n_19),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_105),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_103),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_74),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_57),
.C(n_65),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_14),
.A2(n_15),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_33),
.B1(n_55),
.B2(n_56),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_34),
.C(n_40),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_18),
.B(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_20),
.A2(n_22),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_20),
.A2(n_31),
.B(n_61),
.C(n_122),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_21),
.A2(n_25),
.B(n_31),
.C(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_27),
.A2(n_32),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_31),
.A2(n_37),
.B(n_80),
.C(n_81),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_31),
.B(n_43),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_31),
.B(n_62),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_33),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_36),
.B(n_92),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_37),
.A2(n_38),
.B1(n_81),
.B2(n_88),
.Y(n_92)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_39),
.B(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_39),
.B(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_40),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_48),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_54),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_45),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_53),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_51),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_65),
.B1(n_66),
.B2(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_57),
.A2(n_116),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_57),
.B(n_83),
.C(n_126),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_58),
.B(n_62),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_58),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.Y(n_58)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_67),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_84),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_77),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_82),
.B2(n_83),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_83),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_138),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B1(n_101),
.B2(n_102),
.Y(n_84)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B(n_89),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_108),
.C(n_112),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_98),
.A2(n_99),
.B1(n_108),
.B2(n_132),
.Y(n_145)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_117),
.B(n_147),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_113),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_121),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_108),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B(n_111),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_142),
.B(n_146),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_128),
.B(n_141),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_123),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_124),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_125),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B(n_140),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_137),
.B(n_139),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_143),
.B(n_144),
.Y(n_146)
);


endmodule