module fake_ariane_58_n_107 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_16, n_5, n_12, n_15, n_10, n_107);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_107;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx5p33_ASAP7_75t_R g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx2_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_0),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

CKINVDCx5p33_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_R g43 ( 
.A(n_27),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_24),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_21),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_30),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_23),
.B1(n_31),
.B2(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR3xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_20),
.C(n_26),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_42),
.B(n_45),
.C(n_41),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_47),
.B(n_44),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_45),
.B(n_42),
.C(n_44),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_47),
.B(n_44),
.C(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_57),
.B(n_58),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_54),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_53),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

OAI21x1_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_55),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_R g69 ( 
.A(n_65),
.B(n_46),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_R g70 ( 
.A(n_65),
.B(n_48),
.Y(n_70)
);

OAI21x1_ASAP7_75t_SL g71 ( 
.A1(n_63),
.A2(n_54),
.B(n_2),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

AND2x4_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

AOI211xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_63),
.B(n_43),
.C(n_67),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_54),
.B1(n_64),
.B2(n_66),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_54),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_81),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_67),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_67),
.B1(n_73),
.B2(n_66),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_83),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_86),
.Y(n_92)
);

OAI221xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_83),
.B1(n_84),
.B2(n_34),
.C(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_88),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_84),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_71),
.B1(n_34),
.B2(n_84),
.C(n_49),
.Y(n_97)
);

AOI211xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_85),
.B(n_2),
.C(n_3),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_96),
.A2(n_73),
.B(n_6),
.C(n_7),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_92),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_92),
.B(n_94),
.C(n_68),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_94),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_97),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_101),
.B1(n_6),
.B2(n_8),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_68),
.B2(n_49),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_49),
.B1(n_8),
.B2(n_9),
.Y(n_107)
);


endmodule