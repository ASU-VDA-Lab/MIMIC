module real_aes_6504_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_310;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_602;
wire n_552;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_293;
wire n_358;
wire n_397;
wire n_275;
wire n_385;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_498;
wire n_481;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp5_ASAP7_75t_SL g712 ( .A1(n_0), .A2(n_192), .B1(n_314), .B2(n_599), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_1), .B(n_277), .Y(n_276) );
AOI22xp5_ASAP7_75t_SL g660 ( .A1(n_2), .A2(n_50), .B1(n_343), .B2(n_516), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_3), .A2(n_19), .B1(n_508), .B2(n_573), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_4), .A2(n_220), .B1(n_358), .B2(n_360), .C(n_362), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_5), .A2(n_143), .B1(n_306), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_6), .A2(n_107), .B1(n_359), .B2(n_360), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_7), .A2(n_18), .B1(n_445), .B2(n_446), .Y(n_444) );
AOI22xp33_ASAP7_75t_SL g305 ( .A1(n_8), .A2(n_100), .B1(n_306), .B2(n_308), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_9), .Y(n_242) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_10), .A2(n_106), .B1(n_137), .B2(n_373), .C1(n_376), .C2(n_377), .Y(n_372) );
CKINVDCx20_ASAP7_75t_R g429 ( .A(n_11), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_12), .A2(n_120), .B1(n_290), .B2(n_314), .Y(n_682) );
OA22x2_ASAP7_75t_L g419 ( .A1(n_13), .A2(n_420), .B1(n_421), .B2(n_454), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_13), .Y(n_420) );
AOI22xp33_ASAP7_75t_SL g289 ( .A1(n_14), .A2(n_158), .B1(n_290), .B2(n_294), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_15), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_16), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g448 ( .A1(n_17), .A2(n_194), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_20), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_21), .A2(n_211), .B1(n_396), .B2(n_522), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_22), .A2(n_149), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_SL g658 ( .A1(n_23), .A2(n_216), .B1(n_593), .B2(n_659), .Y(n_658) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_24), .A2(n_70), .B1(n_247), .B2(n_248), .Y(n_246) );
INVx1_ASAP7_75t_L g675 ( .A(n_24), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_25), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_26), .A2(n_30), .B1(n_258), .B2(n_263), .Y(n_257) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_27), .A2(n_197), .B1(n_347), .B2(n_504), .C(n_601), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g719 ( .A1(n_28), .A2(n_170), .B1(n_477), .B2(n_649), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_29), .A2(n_89), .B1(n_136), .B2(n_377), .C1(n_614), .C2(n_615), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_31), .Y(n_597) );
AOI22xp5_ASAP7_75t_SL g652 ( .A1(n_32), .A2(n_119), .B1(n_581), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_33), .A2(n_48), .B1(n_562), .B2(n_563), .Y(n_561) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_34), .A2(n_108), .B1(n_165), .B2(n_562), .C1(n_563), .C2(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_35), .A2(n_214), .B1(n_284), .B2(n_376), .Y(n_691) );
AO22x2_ASAP7_75t_L g250 ( .A1(n_36), .A2(n_71), .B1(n_247), .B2(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g676 ( .A(n_36), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_37), .Y(n_353) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_38), .A2(n_196), .B1(n_303), .B2(n_498), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_39), .A2(n_160), .B1(n_343), .B2(n_494), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g489 ( .A1(n_40), .A2(n_84), .B1(n_446), .B2(n_490), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_41), .A2(n_54), .B1(n_520), .B2(n_522), .Y(n_519) );
AOI222xp33_ASAP7_75t_L g523 ( .A1(n_42), .A2(n_134), .B1(n_177), .B2(n_377), .C1(n_524), .C2(n_525), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_43), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_44), .A2(n_135), .B1(n_581), .B2(n_593), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_45), .A2(n_221), .B1(n_495), .B2(n_599), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_46), .Y(n_611) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_47), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_49), .A2(n_198), .B1(n_581), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_SL g628 ( .A1(n_51), .A2(n_116), .B1(n_284), .B2(n_522), .Y(n_628) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_52), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_53), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_55), .A2(n_159), .B1(n_294), .B2(n_299), .Y(n_544) );
AOI22xp5_ASAP7_75t_SL g710 ( .A1(n_56), .A2(n_128), .B1(n_352), .B2(n_405), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_57), .B(n_359), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_58), .A2(n_121), .B1(n_486), .B2(n_591), .C(n_594), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_59), .A2(n_123), .B1(n_607), .B2(n_609), .C(n_610), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_60), .A2(n_185), .B1(n_352), .B2(n_452), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_61), .A2(n_207), .B1(n_649), .B2(n_650), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_62), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g311 ( .A1(n_63), .A2(n_132), .B1(n_312), .B2(n_314), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g319 ( .A1(n_64), .A2(n_320), .B1(n_378), .B2(n_379), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g378 ( .A(n_64), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_65), .A2(n_589), .B1(n_616), .B2(n_617), .Y(n_588) );
INVx1_ASAP7_75t_L g616 ( .A(n_65), .Y(n_616) );
AOI22xp5_ASAP7_75t_SL g708 ( .A1(n_66), .A2(n_115), .B1(n_508), .B2(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_67), .A2(n_179), .B1(n_277), .B2(n_359), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g397 ( .A(n_68), .Y(n_397) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_69), .Y(n_435) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_72), .Y(n_327) );
AOI22xp33_ASAP7_75t_SL g412 ( .A1(n_73), .A2(n_174), .B1(n_294), .B2(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_74), .A2(n_153), .B1(n_486), .B2(n_488), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_75), .B(n_358), .Y(n_647) );
INVx1_ASAP7_75t_L g230 ( .A(n_76), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_77), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_78), .Y(n_603) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_79), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_80), .A2(n_180), .B1(n_392), .B2(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_81), .A2(n_157), .B1(n_312), .B2(n_314), .Y(n_533) );
INVx1_ASAP7_75t_L g226 ( .A(n_82), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_83), .A2(n_95), .B1(n_506), .B2(n_571), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_85), .A2(n_223), .B(n_231), .C(n_677), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_86), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_87), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g557 ( .A(n_88), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_90), .A2(n_142), .B1(n_359), .B2(n_402), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_91), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g399 ( .A1(n_92), .A2(n_113), .B1(n_263), .B2(n_400), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_93), .A2(n_122), .B1(n_446), .B2(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_94), .A2(n_112), .B1(n_280), .B2(n_284), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_96), .A2(n_178), .B1(n_415), .B2(n_571), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g393 ( .A(n_97), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_98), .A2(n_105), .B1(n_504), .B2(n_506), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_99), .A2(n_146), .B1(n_258), .B2(n_642), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_101), .A2(n_140), .B1(n_290), .B2(n_624), .Y(n_623) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_102), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g532 ( .A1(n_103), .A2(n_182), .B1(n_307), .B2(n_491), .Y(n_532) );
AOI22xp33_ASAP7_75t_SL g414 ( .A1(n_104), .A2(n_152), .B1(n_325), .B2(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_109), .A2(n_147), .B1(n_258), .B2(n_264), .Y(n_717) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_110), .A2(n_184), .B1(n_405), .B2(n_406), .Y(n_404) );
XOR2x2_ASAP7_75t_L g460 ( .A(n_111), .B(n_461), .Y(n_460) );
XNOR2x2_ASAP7_75t_L g500 ( .A(n_114), .B(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_117), .Y(n_640) );
AND2x2_ASAP7_75t_L g229 ( .A(n_118), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g316 ( .A(n_124), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_125), .B(n_277), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_126), .A2(n_215), .B1(n_490), .B2(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_127), .B(n_608), .Y(n_689) );
AND2x6_ASAP7_75t_L g225 ( .A(n_129), .B(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_129), .Y(n_669) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_130), .A2(n_189), .B1(n_247), .B2(n_251), .Y(n_254) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_131), .A2(n_172), .B1(n_290), .B2(n_347), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_133), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_138), .A2(n_208), .B1(n_396), .B2(n_522), .Y(n_687) );
AOI22xp5_ASAP7_75t_SL g654 ( .A1(n_139), .A2(n_188), .B1(n_655), .B2(n_656), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g602 ( .A(n_141), .Y(n_602) );
CKINVDCx20_ASAP7_75t_R g350 ( .A(n_144), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_145), .A2(n_176), .B1(n_281), .B2(n_284), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_148), .B(n_269), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_150), .Y(n_595) );
AO22x2_ASAP7_75t_L g256 ( .A1(n_151), .A2(n_200), .B1(n_247), .B2(n_248), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_154), .A2(n_219), .B1(n_299), .B2(n_508), .Y(n_695) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_155), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_156), .A2(n_186), .B1(n_299), .B2(n_301), .Y(n_298) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_161), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_162), .A2(n_181), .B1(n_515), .B2(n_516), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_163), .Y(n_626) );
INVx1_ASAP7_75t_L g661 ( .A(n_164), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_166), .Y(n_481) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_167), .A2(n_171), .B1(n_336), .B2(n_409), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g425 ( .A(n_168), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_169), .A2(n_217), .B1(n_306), .B2(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_173), .B(n_277), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g345 ( .A(n_175), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_183), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_187), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_189), .B(n_674), .Y(n_673) );
OA22x2_ASAP7_75t_L g385 ( .A1(n_190), .A2(n_386), .B1(n_387), .B2(n_417), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_190), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_191), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g363 ( .A(n_193), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g686 ( .A(n_195), .Y(n_686) );
CKINVDCx20_ASAP7_75t_R g536 ( .A(n_199), .Y(n_536) );
INVx1_ASAP7_75t_L g672 ( .A(n_200), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_201), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_202), .B(n_477), .Y(n_476) );
OA22x2_ASAP7_75t_L g547 ( .A1(n_203), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_547) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_203), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_204), .B(n_358), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_205), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g678 ( .A1(n_206), .A2(n_679), .B1(n_680), .B2(n_696), .Y(n_678) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_206), .Y(n_696) );
INVx1_ASAP7_75t_L g247 ( .A(n_209), .Y(n_247) );
INVx1_ASAP7_75t_L g249 ( .A(n_209), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_210), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_212), .B(n_646), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_213), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g390 ( .A(n_218), .Y(n_390) );
INVx1_ASAP7_75t_SL g223 ( .A(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_226), .Y(n_668) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_227), .A2(n_667), .B(n_704), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_228), .Y(n_227) );
INVxp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_585), .B1(n_586), .B2(n_663), .C(n_664), .Y(n_231) );
INVx1_ASAP7_75t_L g663 ( .A(n_232), .Y(n_663) );
XOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_455), .Y(n_232) );
OAI22xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_235), .B1(n_381), .B2(n_382), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_317), .B1(n_318), .B2(n_380), .Y(n_235) );
INVx1_ASAP7_75t_L g380 ( .A(n_236), .Y(n_380) );
INVx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
XOR2x2_ASAP7_75t_L g238 ( .A(n_239), .B(n_316), .Y(n_238) );
NAND2x1p5_ASAP7_75t_L g239 ( .A(n_240), .B(n_287), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_267), .Y(n_240) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_257), .Y(n_241) );
OAI21xp33_ASAP7_75t_L g428 ( .A1(n_243), .A2(n_429), .B(n_430), .Y(n_428) );
OAI221xp5_ASAP7_75t_L g471 ( .A1(n_243), .A2(n_472), .B1(n_473), .B2(n_475), .C(n_476), .Y(n_471) );
OAI21xp5_ASAP7_75t_L g715 ( .A1(n_243), .A2(n_716), .B(n_717), .Y(n_715) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx4_ASAP7_75t_L g375 ( .A(n_244), .Y(n_375) );
BUFx3_ASAP7_75t_L g524 ( .A(n_244), .Y(n_524) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_244), .Y(n_634) );
AND2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_252), .Y(n_244) );
AND2x4_ASAP7_75t_L g264 ( .A(n_245), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g370 ( .A(n_245), .Y(n_370) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_250), .Y(n_245) );
AND2x2_ASAP7_75t_L g262 ( .A(n_246), .B(n_254), .Y(n_262) );
INVx2_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g251 ( .A(n_249), .Y(n_251) );
OR2x2_ASAP7_75t_L g274 ( .A(n_250), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g278 ( .A(n_250), .B(n_275), .Y(n_278) );
INVx2_ASAP7_75t_L g283 ( .A(n_250), .Y(n_283) );
INVx1_ASAP7_75t_L g286 ( .A(n_250), .Y(n_286) );
AND2x2_ASAP7_75t_L g300 ( .A(n_252), .B(n_293), .Y(n_300) );
AND2x6_ASAP7_75t_L g303 ( .A(n_252), .B(n_273), .Y(n_303) );
AND2x4_ASAP7_75t_L g307 ( .A(n_252), .B(n_278), .Y(n_307) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_255), .Y(n_252) );
AND2x2_ASAP7_75t_L g272 ( .A(n_253), .B(n_256), .Y(n_272) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g292 ( .A(n_254), .B(n_266), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_254), .B(n_256), .Y(n_297) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g261 ( .A(n_256), .Y(n_261) );
INVx1_ASAP7_75t_L g266 ( .A(n_256), .Y(n_266) );
BUFx4f_ASAP7_75t_SL g377 ( .A(n_258), .Y(n_377) );
INVx2_ASAP7_75t_L g564 ( .A(n_258), .Y(n_564) );
BUFx12f_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_259), .Y(n_396) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_259), .Y(n_433) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_261), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g281 ( .A(n_262), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g284 ( .A(n_262), .B(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_L g366 ( .A(n_262), .B(n_315), .Y(n_366) );
BUFx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_264), .Y(n_522) );
BUFx2_ASAP7_75t_SL g650 ( .A(n_264), .Y(n_650) );
INVx1_ASAP7_75t_L g371 ( .A(n_265), .Y(n_371) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_268), .B(n_276), .C(n_279), .Y(n_267) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx5_ASAP7_75t_L g359 ( .A(n_270), .Y(n_359) );
INVx2_ASAP7_75t_L g608 ( .A(n_270), .Y(n_608) );
INVx4_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x6_ASAP7_75t_L g277 ( .A(n_272), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g313 ( .A(n_272), .B(n_293), .Y(n_313) );
INVx1_ASAP7_75t_L g438 ( .A(n_272), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_272), .B(n_278), .Y(n_442) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g437 ( .A(n_274), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g293 ( .A(n_275), .B(n_283), .Y(n_293) );
INVx1_ASAP7_75t_SL g361 ( .A(n_277), .Y(n_361) );
BUFx2_ASAP7_75t_L g402 ( .A(n_277), .Y(n_402) );
BUFx4f_ASAP7_75t_L g609 ( .A(n_277), .Y(n_609) );
AND2x2_ASAP7_75t_L g310 ( .A(n_278), .B(n_292), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_278), .B(n_292), .Y(n_333) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_280), .Y(n_615) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx4f_ASAP7_75t_SL g376 ( .A(n_281), .Y(n_376) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_281), .Y(n_392) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_281), .Y(n_477) );
BUFx2_ASAP7_75t_L g525 ( .A(n_281), .Y(n_525) );
INVx1_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
BUFx2_ASAP7_75t_L g400 ( .A(n_284), .Y(n_400) );
INVx1_ASAP7_75t_L g521 ( .A(n_284), .Y(n_521) );
BUFx3_ASAP7_75t_L g649 ( .A(n_284), .Y(n_649) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x6_ASAP7_75t_L g338 ( .A(n_286), .B(n_297), .Y(n_338) );
NOR2x1_ASAP7_75t_L g287 ( .A(n_288), .B(n_304), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_298), .Y(n_288) );
BUFx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
BUFx3_ASAP7_75t_L g407 ( .A(n_291), .Y(n_407) );
BUFx3_ASAP7_75t_L g498 ( .A(n_291), .Y(n_498) );
BUFx3_ASAP7_75t_L g593 ( .A(n_291), .Y(n_593) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_292), .B(n_293), .Y(n_356) );
AND2x4_ASAP7_75t_L g295 ( .A(n_293), .B(n_296), .Y(n_295) );
BUFx3_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx3_ASAP7_75t_L g329 ( .A(n_295), .Y(n_329) );
BUFx2_ASAP7_75t_SL g450 ( .A(n_295), .Y(n_450) );
BUFx2_ASAP7_75t_SL g488 ( .A(n_295), .Y(n_488) );
BUFx3_ASAP7_75t_L g506 ( .A(n_295), .Y(n_506) );
INVx1_ASAP7_75t_L g583 ( .A(n_295), .Y(n_583) );
BUFx3_ASAP7_75t_L g599 ( .A(n_295), .Y(n_599) );
BUFx2_ASAP7_75t_L g659 ( .A(n_295), .Y(n_659) );
AND2x2_ASAP7_75t_L g314 ( .A(n_296), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx3_ASAP7_75t_L g487 ( .A(n_299), .Y(n_487) );
BUFx3_ASAP7_75t_L g511 ( .A(n_299), .Y(n_511) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx2_ASAP7_75t_SL g352 ( .A(n_300), .Y(n_352) );
INVx2_ASAP7_75t_L g416 ( .A(n_300), .Y(n_416) );
BUFx2_ASAP7_75t_SL g653 ( .A(n_300), .Y(n_653) );
INVx5_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g413 ( .A(n_302), .Y(n_413) );
INVx4_ASAP7_75t_L g515 ( .A(n_302), .Y(n_515) );
INVx2_ASAP7_75t_L g571 ( .A(n_302), .Y(n_571) );
INVx2_ASAP7_75t_SL g694 ( .A(n_302), .Y(n_694) );
INVx11_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx11_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_311), .Y(n_304) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx6_ASAP7_75t_L g348 ( .A(n_307), .Y(n_348) );
BUFx3_ASAP7_75t_L g405 ( .A(n_307), .Y(n_405) );
BUFx2_ASAP7_75t_L g445 ( .A(n_308), .Y(n_445) );
INVx5_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g410 ( .A(n_309), .Y(n_410) );
INVx4_ASAP7_75t_L g491 ( .A(n_309), .Y(n_491) );
INVx3_ASAP7_75t_L g508 ( .A(n_309), .Y(n_508) );
INVx8_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx4_ASAP7_75t_L g505 ( .A(n_312), .Y(n_505) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
BUFx3_ASAP7_75t_L g326 ( .A(n_313), .Y(n_326) );
INVx2_ASAP7_75t_L g453 ( .A(n_313), .Y(n_453) );
BUFx3_ASAP7_75t_L g495 ( .A(n_313), .Y(n_495) );
BUFx3_ASAP7_75t_L g581 ( .A(n_313), .Y(n_581) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g379 ( .A(n_320), .Y(n_379) );
AND4x1_ASAP7_75t_L g320 ( .A(n_321), .B(n_339), .C(n_357), .D(n_372), .Y(n_320) );
NOR2xp33_ASAP7_75t_SL g321 ( .A(n_322), .B(n_330), .Y(n_321) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_327), .B2(n_328), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_332), .B1(n_334), .B2(n_335), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_332), .A2(n_602), .B1(n_603), .B2(n_604), .Y(n_601) );
BUFx2_ASAP7_75t_R g332 ( .A(n_333), .Y(n_332) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g573 ( .A(n_337), .Y(n_573) );
BUFx2_ASAP7_75t_L g605 ( .A(n_337), .Y(n_605) );
BUFx2_ASAP7_75t_L g656 ( .A(n_337), .Y(n_656) );
INVx6_ASAP7_75t_SL g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g446 ( .A(n_338), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_349), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_345), .B2(n_346), .Y(n_340) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx4_ASAP7_75t_L g449 ( .A(n_344), .Y(n_449) );
INVx3_ASAP7_75t_L g709 ( .A(n_344), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_346), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g516 ( .A(n_348), .Y(n_516) );
INVx3_ASAP7_75t_L g631 ( .A(n_348), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_353), .B2(n_354), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g577 ( .A(n_355), .Y(n_577) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g646 ( .A(n_361), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_367), .B2(n_368), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_364), .A2(n_368), .B1(n_611), .B2(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx4_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_366), .A2(n_424), .B1(n_425), .B2(n_426), .Y(n_423) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_366), .Y(n_480) );
OAI22xp33_ASAP7_75t_SL g565 ( .A1(n_366), .A2(n_482), .B1(n_566), .B2(n_567), .Y(n_565) );
BUFx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_369), .Y(n_427) );
OR2x6_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI222xp33_ASAP7_75t_L g389 ( .A1(n_374), .A2(n_390), .B1(n_391), .B2(n_393), .C1(n_394), .C2(n_397), .Y(n_389) );
BUFx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g535 ( .A1(n_375), .A2(n_536), .B(n_537), .Y(n_535) );
INVx4_ASAP7_75t_L g614 ( .A(n_375), .Y(n_614) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_375), .A2(n_640), .B(n_641), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g685 ( .A1(n_375), .A2(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B1(n_418), .B2(n_419), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_403), .C(n_411), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_398), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx4f_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_399), .B(n_401), .Y(n_398) );
AND2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_408), .Y(n_403) );
BUFx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx3_ASAP7_75t_L g624 ( .A(n_416), .Y(n_624) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g454 ( .A(n_421), .Y(n_454) );
NAND2x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_443), .Y(n_421) );
NOR3xp33_ASAP7_75t_SL g422 ( .A(n_423), .B(n_428), .C(n_434), .Y(n_422) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g482 ( .A(n_427), .Y(n_482) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g474 ( .A(n_433), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_436), .B1(n_439), .B2(n_440), .Y(n_434) );
INVx1_ASAP7_75t_L g554 ( .A(n_436), .Y(n_554) );
BUFx6f_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g466 ( .A(n_437), .Y(n_466) );
OA211x2_ASAP7_75t_L g625 ( .A1(n_440), .A2(n_626), .B(n_627), .C(n_628), .Y(n_625) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx3_ASAP7_75t_L g470 ( .A(n_442), .Y(n_470) );
AND4x1_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .C(n_448), .D(n_451), .Y(n_443) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_456), .A2(n_457), .B1(n_526), .B2(n_527), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_460), .B1(n_499), .B2(n_500), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_462), .B(n_483), .Y(n_461) );
NOR3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_471), .C(n_478), .Y(n_462) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_465), .B1(n_467), .B2(n_468), .Y(n_463) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g556 ( .A(n_470), .Y(n_556) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g562 ( .A(n_477), .Y(n_562) );
INVx4_ASAP7_75t_L g643 ( .A(n_477), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_480), .B1(n_481), .B2(n_482), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_492), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_489), .Y(n_484) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
BUFx2_ASAP7_75t_L g655 ( .A(n_491), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .Y(n_492) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx4f_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g513 ( .A(n_498), .Y(n_513) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND4xp75_ASAP7_75t_L g501 ( .A(n_502), .B(n_509), .C(n_517), .D(n_523), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_507), .Y(n_502) );
INVx4_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_SL g596 ( .A(n_515), .Y(n_596) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx3_ASAP7_75t_L g559 ( .A(n_524), .Y(n_559) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_546), .B1(n_547), .B2(n_584), .Y(n_528) );
INVx3_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
XOR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_545), .Y(n_529) );
NAND3x1_ASAP7_75t_SL g530 ( .A(n_531), .B(n_534), .C(n_542), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NOR2x1_ASAP7_75t_L g534 ( .A(n_535), .B(n_538), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .C(n_541), .Y(n_538) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_568), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_558), .C(n_565), .Y(n_551) );
OAI22xp5_ASAP7_75t_SL g552 ( .A1(n_553), .A2(n_555), .B1(n_556), .B2(n_557), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI21xp33_ASAP7_75t_SL g558 ( .A1(n_559), .A2(n_560), .B(n_561), .Y(n_558) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_569), .B(n_574), .C(n_578), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_580), .B1(n_582), .B2(n_583), .Y(n_578) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
CKINVDCx14_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B1(n_618), .B2(n_662), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g617 ( .A(n_589), .Y(n_617) );
AND4x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_600), .C(n_606), .D(n_613), .Y(n_589) );
INVx2_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_594) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g662 ( .A(n_618), .Y(n_662) );
XNOR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_636), .Y(n_618) );
XOR2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_635), .Y(n_619) );
NAND4xp75_ASAP7_75t_L g620 ( .A(n_621), .B(n_625), .C(n_629), .D(n_633), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_661), .Y(n_636) );
NAND3x1_ASAP7_75t_L g637 ( .A(n_638), .B(n_651), .C(n_657), .Y(n_637) );
NOR2x1_ASAP7_75t_L g638 ( .A(n_639), .B(n_644), .Y(n_638) );
INVx3_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .C(n_648), .Y(n_644) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_670), .Y(n_665) );
OR2x2_ASAP7_75t_SL g723 ( .A(n_666), .B(n_671), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_668), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_668), .B(n_701), .Y(n_704) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_669), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_697), .A3(n_698), .B1(n_702), .B2(n_705), .C1(n_706), .C2(n_721), .Y(n_677) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
NAND3x1_ASAP7_75t_L g680 ( .A(n_681), .B(n_684), .C(n_692), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
NOR2x1_ASAP7_75t_L g684 ( .A(n_685), .B(n_688), .Y(n_684) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .C(n_691), .Y(n_688) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
BUFx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
XOR2x2_ASAP7_75t_L g706 ( .A(n_705), .B(n_707), .Y(n_706) );
NAND4xp75_ASAP7_75t_SL g707 ( .A(n_708), .B(n_710), .C(n_711), .D(n_714), .Y(n_707) );
AND2x2_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_719), .B(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
endmodule