module fake_jpeg_10114_n_299 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_299);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_299;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_36),
.Y(n_48)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_16),
.B1(n_32),
.B2(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_31),
.B1(n_27),
.B2(n_32),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_66),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_23),
.C(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_51),
.Y(n_84)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_53),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_56),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_17),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_40),
.A2(n_30),
.B1(n_17),
.B2(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_30),
.B1(n_38),
.B2(n_37),
.Y(n_78)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_30),
.B1(n_16),
.B2(n_18),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_21),
.B1(n_28),
.B2(n_25),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_34),
.C(n_38),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_89),
.C(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_53),
.A2(n_19),
.B1(n_24),
.B2(n_20),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_81),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_30),
.B1(n_17),
.B2(n_28),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_55),
.A2(n_37),
.B1(n_38),
.B2(n_34),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_78),
.B1(n_87),
.B2(n_62),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_42),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_10),
.B1(n_9),
.B2(n_11),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_62),
.B1(n_60),
.B2(n_46),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_25),
.B(n_33),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_91),
.B(n_25),
.C(n_28),
.Y(n_114)
);

NAND2x1_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_115),
.B1(n_68),
.B2(n_91),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_61),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_94),
.B(n_110),
.C(n_113),
.Y(n_143)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_102),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_105),
.B1(n_107),
.B2(n_69),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_99),
.B(n_103),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_74),
.B1(n_78),
.B2(n_71),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_88),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_91),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_64),
.B1(n_47),
.B2(n_54),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_112),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_45),
.C(n_64),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_91),
.B(n_21),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_74),
.A2(n_49),
.B1(n_51),
.B2(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_67),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

CKINVDCx12_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_14),
.C(n_13),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_112),
.A2(n_73),
.B1(n_85),
.B2(n_87),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_131),
.B(n_68),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_123),
.B1(n_80),
.B2(n_83),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_69),
.B1(n_80),
.B2(n_83),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_125),
.A2(n_96),
.B1(n_105),
.B2(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_127),
.Y(n_151)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_137),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_129),
.B(n_45),
.Y(n_169)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_80),
.B(n_45),
.C(n_43),
.Y(n_137)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_140),
.Y(n_149)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_141),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_167),
.B1(n_119),
.B2(n_138),
.Y(n_176)
);

INVx2_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_146),
.B(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_152),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_143),
.B(n_124),
.C(n_129),
.D(n_94),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_169),
.Y(n_180)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_160),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_104),
.C(n_110),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_122),
.C(n_134),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_126),
.B(n_99),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_101),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_168),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_146),
.B(n_148),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_166),
.B1(n_135),
.B2(n_72),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_100),
.B1(n_93),
.B2(n_45),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_100),
.B1(n_45),
.B2(n_65),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_135),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_136),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_175),
.C(n_186),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_142),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_185),
.B(n_153),
.Y(n_200)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_138),
.B(n_122),
.C(n_43),
.D(n_63),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_168),
.A2(n_144),
.B1(n_160),
.B2(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_195),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_63),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_162),
.A2(n_145),
.B1(n_167),
.B2(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_140),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_134),
.C(n_141),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_SL g197 ( 
.A1(n_192),
.A2(n_166),
.B(n_161),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_72),
.B1(n_28),
.B2(n_21),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_152),
.B(n_33),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_196),
.A2(n_197),
.B1(n_211),
.B2(n_213),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_164),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_155),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_185),
.A2(n_149),
.B(n_170),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_149),
.Y(n_209)
);

OAI31xp33_ASAP7_75t_L g221 ( 
.A1(n_209),
.A2(n_177),
.A3(n_172),
.B(n_188),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_157),
.B1(n_72),
.B2(n_3),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_1),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_215),
.B1(n_173),
.B2(n_181),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_171),
.A2(n_72),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_33),
.B1(n_22),
.B2(n_12),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_184),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_184),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_216),
.A2(n_10),
.B1(n_2),
.B2(n_4),
.Y(n_237)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_33),
.Y(n_217)
);

XNOR2x1_ASAP7_75t_L g228 ( 
.A(n_217),
.B(n_194),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_9),
.B(n_14),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_11),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_186),
.C(n_174),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_227),
.C(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_180),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_231),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_214),
.C(n_180),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_228),
.B(n_235),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_187),
.C(n_175),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_176),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_33),
.C(n_22),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_236),
.C(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_213),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_22),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_217),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_202),
.C(n_199),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_212),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_215),
.B(n_199),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_210),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_201),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_201),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_249),
.B(n_218),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_229),
.A2(n_198),
.B(n_206),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_222),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_228),
.A2(n_198),
.B1(n_203),
.B2(n_217),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_235),
.B1(n_234),
.B2(n_210),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_232),
.C(n_220),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_241),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_244),
.A2(n_231),
.B1(n_203),
.B2(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_241),
.C(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_239),
.B(n_216),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_263),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_252),
.A2(n_227),
.B(n_230),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_211),
.B1(n_223),
.B2(n_4),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_264),
.B(n_242),
.Y(n_269)
);

AO221x1_ASAP7_75t_L g265 ( 
.A1(n_251),
.A2(n_10),
.B1(n_2),
.B2(n_5),
.C(n_6),
.Y(n_265)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_265),
.Y(n_276)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_258),
.A2(n_245),
.B(n_247),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_1),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_269),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_256),
.A2(n_247),
.B(n_238),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_259),
.B(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_273),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_22),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_276),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_254),
.B1(n_258),
.B2(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_277),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_276),
.B1(n_270),
.B2(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_271),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_6),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_282),
.B(n_7),
.Y(n_290)
);

OAI21xp33_ASAP7_75t_L g287 ( 
.A1(n_283),
.A2(n_1),
.B(n_5),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_272),
.B(n_266),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_290),
.B(n_283),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_280),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.C(n_7),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_281),
.C(n_278),
.Y(n_293)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_8),
.B(n_291),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_8),
.C(n_293),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_298),
.B(n_8),
.Y(n_299)
);


endmodule