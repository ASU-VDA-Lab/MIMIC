module fake_jpeg_17629_n_246 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_36),
.Y(n_46)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_26),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_28),
.B1(n_21),
.B2(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_22),
.B1(n_23),
.B2(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_59),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_21),
.B1(n_28),
.B2(n_17),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_57),
.B1(n_22),
.B2(n_23),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_19),
.Y(n_52)
);

OR2x2_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_53),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_19),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_19),
.Y(n_54)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_32),
.C(n_27),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_28),
.B1(n_17),
.B2(n_27),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_18),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_26),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_65),
.B1(n_24),
.B2(n_32),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_54),
.B1(n_53),
.B2(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_66),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_41),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_74),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_73),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_41),
.Y(n_75)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_53),
.B(n_42),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_61),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_23),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_16),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_18),
.Y(n_98)
);

AND2x6_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_54),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_91),
.B1(n_96),
.B2(n_102),
.Y(n_130)
);

NOR4xp25_ASAP7_75t_SL g91 ( 
.A(n_71),
.B(n_0),
.C(n_1),
.D(n_2),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_64),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_97),
.B1(n_107),
.B2(n_70),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_40),
.B1(n_51),
.B2(n_63),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_29),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_66),
.B(n_0),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_110),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_40),
.B1(n_26),
.B2(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_63),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_109),
.B(n_85),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_89),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_109),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_119),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_122),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_121),
.B(n_124),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_100),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_72),
.A3(n_84),
.B1(n_69),
.B2(n_78),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_82),
.B1(n_70),
.B2(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_123),
.A2(n_130),
.B1(n_132),
.B2(n_108),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_76),
.B(n_20),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_76),
.B(n_20),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_87),
.B(n_97),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_69),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_127),
.B(n_101),
.Y(n_136)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_131),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_77),
.B1(n_45),
.B2(n_63),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_73),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_134),
.C(n_93),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_55),
.C(n_47),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_136),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_141),
.A2(n_151),
.B(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_90),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_145),
.Y(n_167)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_96),
.Y(n_145)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_93),
.B(n_101),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_120),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_155),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_91),
.B(n_103),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_105),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_139),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_161),
.B(n_168),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_163),
.Y(n_184)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_170),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_115),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_129),
.B1(n_122),
.B2(n_119),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_178),
.B1(n_144),
.B2(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_126),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_173),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_147),
.B(n_118),
.Y(n_174)
);

NAND3xp33_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_138),
.C(n_98),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_129),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_150),
.Y(n_183)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_192),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_178),
.A2(n_156),
.B1(n_145),
.B2(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_186),
.A2(n_189),
.B1(n_191),
.B2(n_176),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_142),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_194),
.C(n_175),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_160),
.A2(n_152),
.B1(n_157),
.B2(n_137),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_150),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_171),
.B(n_173),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_161),
.A2(n_141),
.B1(n_154),
.B2(n_132),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_168),
.A2(n_26),
.B1(n_51),
.B2(n_25),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_20),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_164),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_51),
.C(n_20),
.Y(n_194)
);

BUFx12f_ASAP7_75t_SL g197 ( 
.A(n_196),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_180),
.B(n_175),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_162),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_0),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_179),
.B(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_207),
.B(n_209),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_163),
.C(n_171),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_193),
.C(n_183),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_202),
.A2(n_187),
.B1(n_176),
.B2(n_190),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_200),
.Y(n_227)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_212),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_194),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_216),
.A2(n_210),
.B(n_218),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_201),
.C(n_208),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_1),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_227),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_198),
.C(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_225),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_224),
.B(n_226),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_197),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_203),
.B(n_213),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_230),
.B(n_231),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_25),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_25),
.Y(n_235)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_232),
.A2(n_222),
.B(n_229),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g239 ( 
.A1(n_234),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_239)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_237),
.A3(n_238),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_SL g237 ( 
.A(n_231),
.B(n_1),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_228),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_3),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_20),
.C(n_9),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_8),
.Y(n_244)
);

OAI32xp33_ASAP7_75t_L g245 ( 
.A1(n_244),
.A2(n_243),
.A3(n_11),
.B1(n_13),
.B2(n_10),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_10),
.Y(n_246)
);


endmodule