module real_jpeg_30505_n_11 (n_108, n_8, n_0, n_2, n_10, n_9, n_107, n_6, n_104, n_100, n_106, n_7, n_3, n_99, n_5, n_4, n_102, n_105, n_101, n_1, n_103, n_11);

input n_108;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_107;
input n_6;
input n_104;
input n_100;
input n_106;
input n_7;
input n_3;
input n_99;
input n_5;
input n_4;
input n_102;
input n_105;
input n_101;
input n_1;
input n_103;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_0),
.B(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_0),
.Y(n_96)
);

AOI221xp5_ASAP7_75t_L g56 ( 
.A1(n_1),
.A2(n_10),
.B1(n_57),
.B2(n_61),
.C(n_62),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_3),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_5),
.Y(n_76)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_6),
.B(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_8),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_86),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_9),
.B(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_10),
.B(n_57),
.C(n_61),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_21),
.Y(n_11)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_99),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_28),
.B(n_94),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_23),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_26),
.B(n_105),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_37),
.B(n_92),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_85),
.B(n_91),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_47),
.B(n_83),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_76),
.C(n_77),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_66),
.B(n_75),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_56),
.B1(n_64),
.B2(n_65),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_58),
.B(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_74),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_74),
.Y(n_75)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_100),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_101),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_102),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_103),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_104),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_106),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_107),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_108),
.Y(n_87)
);


endmodule