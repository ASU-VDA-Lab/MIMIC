module fake_ariane_2792_n_1954 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1954);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1954;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1920;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_1901;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_887;
wire n_729;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1937;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_1),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_45),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_40),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_77),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_106),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_14),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_59),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_39),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_86),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_156),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_94),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_76),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_124),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_55),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_36),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_16),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_51),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_171),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_52),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_154),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_83),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_131),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_148),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_174),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_181),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_0),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_4),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_44),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_99),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_36),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_125),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_190),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_92),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_109),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_44),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_62),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_98),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_50),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_139),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_31),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_25),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_8),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_6),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_64),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_13),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_69),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_71),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_169),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_48),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_23),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_8),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_185),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_82),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_2),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_194),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_9),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_165),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_111),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_87),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_147),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_136),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_123),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_186),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_70),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_66),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_97),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_189),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_129),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_164),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_153),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_20),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_85),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_184),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_27),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_102),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_158),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_45),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_90),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_93),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_31),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_161),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_67),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_26),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_127),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_101),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_29),
.Y(n_307)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_17),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_193),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_37),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_37),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_57),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_57),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_121),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_105),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_5),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_24),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_73),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_66),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_49),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_3),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_146),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_62),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_15),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_21),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_80),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_32),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_72),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_68),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_157),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_187),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_34),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_107),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_138),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_50),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_115),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_177),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_38),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_119),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_43),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_29),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_0),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_75),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_26),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_195),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_79),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_166),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_176),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_2),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_3),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_17),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_30),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_137),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_63),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_52),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_56),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_54),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_150),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_24),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_16),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_6),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_168),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_149),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_33),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_18),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_141),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_100),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_65),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_35),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_23),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_30),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_27),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_114),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_160),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_126),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_21),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_18),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_56),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_132),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_32),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_63),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_122),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_188),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_155),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_53),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_60),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_28),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_34),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_49),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_219),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_200),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_263),
.B(n_5),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_228),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_200),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_253),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_267),
.Y(n_398)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_318),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_328),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_275),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_241),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_267),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_361),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_203),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_203),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_220),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_329),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_308),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_256),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_223),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_349),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_227),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_251),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_327),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_272),
.Y(n_417)
);

INVxp67_ASAP7_75t_SL g418 ( 
.A(n_329),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_281),
.B(n_254),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_203),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_349),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_279),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_197),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_198),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_257),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_286),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_261),
.Y(n_429)
);

INVxp33_ASAP7_75t_SL g430 ( 
.A(n_197),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_294),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_309),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_198),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_311),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_314),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_202),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_296),
.Y(n_437)
);

INVxp33_ASAP7_75t_SL g438 ( 
.A(n_205),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_383),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_302),
.Y(n_440)
);

INVxp33_ASAP7_75t_SL g441 ( 
.A(n_205),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_202),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_206),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_196),
.B(n_212),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_210),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_320),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_324),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_322),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_254),
.B(n_7),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_206),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_323),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_217),
.B(n_7),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_210),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_337),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_R g457 ( 
.A(n_347),
.B(n_74),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_239),
.B(n_207),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_211),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_207),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_362),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_373),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_374),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_387),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_211),
.Y(n_466)
);

INVxp33_ASAP7_75t_SL g467 ( 
.A(n_209),
.Y(n_467)
);

INVxp67_ASAP7_75t_SL g468 ( 
.A(n_329),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_329),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_369),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_381),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_199),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_359),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_213),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_359),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_204),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_359),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_359),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_213),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_214),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_359),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_372),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_214),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_239),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_215),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_258),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_372),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_283),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_215),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_303),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_307),
.Y(n_491)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_372),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_372),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_372),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_413),
.B(n_349),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_409),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_421),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_421),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_418),
.B(n_221),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_459),
.B(n_316),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_230),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_413),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_469),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_394),
.B(n_405),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_423),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_459),
.B(n_316),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_423),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_232),
.Y(n_516)
);

INVxp33_ASAP7_75t_SL g517 ( 
.A(n_392),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_451),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_451),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_423),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_475),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_475),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_393),
.B(n_355),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_494),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_478),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_481),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_396),
.B(n_355),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g529 ( 
.A(n_482),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_405),
.B(n_231),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_492),
.B(n_233),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_392),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_395),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_487),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_407),
.B(n_231),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_444),
.B(n_237),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_450),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_408),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_414),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_461),
.B(n_244),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_398),
.B(n_239),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_415),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_461),
.B(n_276),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_427),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_429),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_403),
.B(n_216),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_426),
.B(n_433),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_434),
.Y(n_551)
);

NOR3xp33_ASAP7_75t_L g552 ( 
.A(n_453),
.B(n_249),
.C(n_224),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_435),
.A2(n_341),
.B(n_276),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_446),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_448),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_404),
.B(n_245),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_449),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_452),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_456),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_458),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_406),
.B(n_247),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_462),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_463),
.Y(n_564)
);

CKINVDCx14_ASAP7_75t_R g565 ( 
.A(n_407),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_420),
.B(n_341),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_464),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_410),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_419),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_419),
.Y(n_571)
);

NOR2x1_ASAP7_75t_L g572 ( 
.A(n_410),
.B(n_201),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_439),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_416),
.B(n_216),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_535),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_549),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

INVx2_ASAP7_75t_SL g578 ( 
.A(n_503),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_535),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_L g580 ( 
.A(n_549),
.B(n_433),
.C(n_426),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_512),
.B(n_484),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_535),
.Y(n_582)
);

NAND2xp33_ASAP7_75t_SL g583 ( 
.A(n_509),
.B(n_457),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_532),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_552),
.A2(n_416),
.B1(n_401),
.B2(n_430),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_499),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_499),
.Y(n_588)
);

NOR2x1p5_ASAP7_75t_L g589 ( 
.A(n_574),
.B(n_395),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_512),
.B(n_422),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_500),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_509),
.B(n_397),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_530),
.B(n_536),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_543),
.B(n_436),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_503),
.B(n_422),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_543),
.B(n_442),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_535),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_564),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_564),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_500),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_500),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_557),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_521),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_521),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_512),
.B(n_442),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_563),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_518),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_537),
.B(n_208),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_530),
.A2(n_536),
.B1(n_552),
.B2(n_572),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_532),
.Y(n_611)
);

INVx4_ASAP7_75t_SL g612 ( 
.A(n_498),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_537),
.B(n_454),
.C(n_445),
.Y(n_614)
);

AOI21x1_ASAP7_75t_L g615 ( 
.A1(n_553),
.A2(n_287),
.B(n_270),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_563),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_521),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_564),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_505),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_564),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

INVxp67_ASAP7_75t_SL g622 ( 
.A(n_502),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_557),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_548),
.B(n_445),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_454),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_512),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_564),
.Y(n_627)
);

NOR2x1p5_ASAP7_75t_L g628 ( 
.A(n_574),
.B(n_397),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_564),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_503),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_570),
.B(n_400),
.Y(n_631)
);

AND2x6_ASAP7_75t_L g632 ( 
.A(n_512),
.B(n_349),
.Y(n_632)
);

INVx6_ASAP7_75t_L g633 ( 
.A(n_545),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_523),
.B(n_425),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_557),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_545),
.A2(n_401),
.B1(n_441),
.B2(n_438),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_534),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_570),
.B(n_400),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_534),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_534),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_508),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_508),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_548),
.B(n_460),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_460),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_564),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_508),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_569),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_513),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_564),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_513),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_568),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_513),
.Y(n_653)
);

AND2x2_ASAP7_75t_SL g654 ( 
.A(n_532),
.B(n_399),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_524),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_568),
.B(n_208),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_548),
.B(n_466),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_545),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_523),
.B(n_466),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_524),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_570),
.B(n_474),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_524),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_563),
.B(n_474),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_496),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_568),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_570),
.B(n_479),
.Y(n_667)
);

CKINVDCx6p67_ASAP7_75t_R g668 ( 
.A(n_533),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_563),
.B(n_479),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_496),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_574),
.A2(n_273),
.B1(n_377),
.B2(n_299),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_568),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_571),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_568),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_557),
.B(n_480),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_568),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_568),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_568),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_571),
.A2(n_489),
.B1(n_485),
.B2(n_483),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_571),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_571),
.B(n_480),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_501),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_501),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_568),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_502),
.B(n_483),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_526),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_545),
.A2(n_443),
.B1(n_467),
.B2(n_485),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_515),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_504),
.B(n_489),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_573),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_525),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_R g692 ( 
.A(n_517),
.B(n_402),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_526),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_504),
.B(n_360),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_517),
.B(n_222),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_516),
.B(n_411),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_526),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_527),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_533),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_525),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_533),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_525),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_525),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_527),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_527),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_566),
.B(n_209),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_539),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_553),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_518),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_516),
.B(n_417),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_545),
.B(n_349),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_525),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

AND2x6_ASAP7_75t_L g717 ( 
.A(n_545),
.B(n_300),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_525),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_573),
.Y(n_719)
);

OR2x6_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_305),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_531),
.B(n_424),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_566),
.B(n_315),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_525),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_531),
.B(n_428),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_626),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_622),
.B(n_690),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_707),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_690),
.B(n_565),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_719),
.B(n_565),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_673),
.A2(n_539),
.B(n_541),
.C(n_540),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_584),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_692),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_671),
.A2(n_553),
.B1(n_547),
.B2(n_551),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_659),
.B(n_519),
.Y(n_734)
);

INVx8_ASAP7_75t_L g735 ( 
.A(n_632),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_626),
.B(n_519),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_719),
.B(n_572),
.Y(n_737)
);

AOI221x1_ASAP7_75t_L g738 ( 
.A1(n_686),
.A2(n_330),
.B1(n_332),
.B2(n_368),
.C(n_365),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_642),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_610),
.A2(n_573),
.B1(n_313),
.B2(n_550),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_611),
.B(n_569),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_685),
.B(n_540),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_699),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_707),
.Y(n_744)
);

NOR3xp33_ASAP7_75t_L g745 ( 
.A(n_701),
.B(n_225),
.C(n_218),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_642),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_661),
.B(n_573),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_649),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_679),
.B(n_591),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_708),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_580),
.B(n_546),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_591),
.B(n_566),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_591),
.B(n_566),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_708),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_664),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_689),
.B(n_542),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_696),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_649),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_664),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_712),
.B(n_550),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_673),
.B(n_542),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_651),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_648),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_682),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_626),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_634),
.B(n_566),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_651),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_585),
.B(n_567),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_653),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_680),
.B(n_540),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_634),
.B(n_538),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_680),
.A2(n_561),
.B1(n_541),
.B2(n_544),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_634),
.B(n_648),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_682),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_594),
.A2(n_538),
.B1(n_561),
.B2(n_559),
.C(n_541),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_608),
.B(n_538),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_653),
.Y(n_777)
);

A2O1A1Ixp33_ASAP7_75t_L g778 ( 
.A1(n_631),
.A2(n_544),
.B(n_555),
.C(n_558),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_645),
.B(n_544),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_644),
.B(n_555),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_583),
.A2(n_555),
.B1(n_558),
.B2(n_559),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_686),
.Y(n_782)
);

INVx4_ASAP7_75t_L g783 ( 
.A(n_633),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_645),
.B(n_559),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_675),
.B(n_528),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_671),
.A2(n_716),
.B1(n_709),
.B2(n_714),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_621),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_711),
.B(n_528),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_694),
.B(n_639),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_578),
.A2(n_567),
.B(n_547),
.C(n_560),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_645),
.B(n_547),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_578),
.A2(n_556),
.B1(n_562),
.B2(n_218),
.C(n_225),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_583),
.B(n_614),
.C(n_595),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_593),
.A2(n_606),
.B1(n_625),
.B2(n_657),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_637),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_581),
.B(n_528),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_693),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_596),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_693),
.Y(n_800)
);

OR2x6_ASAP7_75t_L g801 ( 
.A(n_671),
.B(n_547),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_581),
.B(n_551),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_697),
.Y(n_803)
);

AOI221xp5_ASAP7_75t_L g804 ( 
.A1(n_586),
.A2(n_671),
.B1(n_636),
.B2(n_687),
.C(n_721),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_630),
.B(n_551),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_697),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_630),
.B(n_551),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_576),
.B(n_554),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_663),
.B(n_554),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_716),
.A2(n_567),
.B1(n_560),
.B2(n_554),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_556),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_576),
.B(n_554),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_637),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_600),
.Y(n_814)
);

OAI21xp5_ASAP7_75t_L g815 ( 
.A1(n_709),
.A2(n_714),
.B(n_710),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_666),
.B(n_724),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_698),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_L g818 ( 
.A(n_600),
.B(n_222),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_698),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_704),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_640),
.Y(n_821)
);

INVx4_ASAP7_75t_L g822 ( 
.A(n_633),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_581),
.A2(n_567),
.B1(n_560),
.B2(n_562),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_585),
.B(n_560),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_576),
.B(n_596),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_654),
.B(n_226),
.Y(n_826)
);

OAI21xp33_ASAP7_75t_L g827 ( 
.A1(n_667),
.A2(n_356),
.B(n_236),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_681),
.B(n_238),
.Y(n_828)
);

BUFx8_ASAP7_75t_L g829 ( 
.A(n_706),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_668),
.B(n_431),
.Y(n_830)
);

AO22x2_ASAP7_75t_L g831 ( 
.A1(n_706),
.A2(n_471),
.B1(n_470),
.B2(n_447),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_640),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_585),
.B(n_226),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_704),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_603),
.A2(n_357),
.B1(n_358),
.B2(n_363),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_654),
.B(n_229),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_597),
.B(n_358),
.C(n_357),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_624),
.B(n_240),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_603),
.B(n_229),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_603),
.B(n_234),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_623),
.B(n_234),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_SL g842 ( 
.A(n_668),
.B(n_437),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_633),
.A2(n_235),
.B1(n_376),
.B2(n_293),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_716),
.A2(n_710),
.B1(n_717),
.B2(n_706),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_705),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_623),
.B(n_235),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_641),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_641),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_695),
.B(n_366),
.C(n_363),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_623),
.B(n_635),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_589),
.Y(n_851)
);

AOI221xp5_ASAP7_75t_L g852 ( 
.A1(n_609),
.A2(n_366),
.B1(n_367),
.B2(n_370),
.C(n_371),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_633),
.B(n_242),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_L g854 ( 
.A(n_600),
.B(n_293),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_577),
.A2(n_336),
.B(n_345),
.C(n_520),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_635),
.B(n_364),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_635),
.B(n_364),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_658),
.B(n_246),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_607),
.B(n_375),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_248),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_607),
.B(n_375),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_616),
.B(n_376),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_658),
.B(n_259),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_616),
.B(n_658),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_717),
.B(n_384),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_717),
.B(n_384),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_688),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_717),
.A2(n_522),
.B1(n_390),
.B2(n_379),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_717),
.B(n_575),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_604),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_717),
.B(n_575),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_720),
.B(n_260),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_600),
.B(n_385),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_628),
.A2(n_587),
.B1(n_588),
.B2(n_577),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_579),
.B(n_385),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_600),
.B(n_386),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_618),
.B(n_629),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_604),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_605),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_720),
.B(n_266),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_605),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_618),
.B(n_386),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_587),
.A2(n_378),
.B1(n_379),
.B2(n_380),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_618),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_705),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_579),
.B(n_582),
.Y(n_886)
);

OAI221xp5_ASAP7_75t_L g887 ( 
.A1(n_720),
.A2(n_378),
.B1(n_380),
.B2(n_382),
.C(n_388),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_588),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_722),
.B(n_268),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_618),
.B(n_382),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_SL g891 ( 
.A(n_722),
.B(n_440),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_850),
.A2(n_678),
.B(n_609),
.Y(n_892)
);

OR2x6_ASAP7_75t_L g893 ( 
.A(n_731),
.B(n_722),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_804),
.A2(n_632),
.B1(n_670),
.B2(n_683),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_760),
.B(n_618),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_773),
.B(n_472),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_725),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_789),
.B(n_722),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_756),
.B(n_632),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_L g900 ( 
.A(n_825),
.B(n_284),
.C(n_271),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_743),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_824),
.A2(n_678),
.B(n_620),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_877),
.A2(n_678),
.B(n_620),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_756),
.B(n_632),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_816),
.B(n_629),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_734),
.B(n_688),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_763),
.Y(n_907)
);

BUFx8_ASAP7_75t_L g908 ( 
.A(n_830),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_877),
.A2(n_620),
.B(n_599),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_725),
.B(n_629),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_741),
.B(n_476),
.Y(n_911)
);

O2A1O1Ixp33_ASAP7_75t_SL g912 ( 
.A1(n_768),
.A2(n_643),
.B(n_647),
.C(n_655),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_810),
.A2(n_601),
.B(n_592),
.Y(n_913)
);

CKINVDCx10_ASAP7_75t_R g914 ( 
.A(n_801),
.Y(n_914)
);

BUFx12f_ASAP7_75t_L g915 ( 
.A(n_732),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_734),
.B(n_688),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_811),
.B(n_632),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_795),
.B(n_799),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_755),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_725),
.B(n_629),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_771),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_811),
.A2(n_780),
.B(n_749),
.C(n_764),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_782),
.A2(n_660),
.B1(n_613),
.B2(n_601),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_725),
.B(n_629),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_870),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_851),
.Y(n_926)
);

NOR2x1_ASAP7_75t_L g927 ( 
.A(n_728),
.B(n_592),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_759),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_809),
.A2(n_627),
.B(n_599),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_774),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_735),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_780),
.B(n_632),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_766),
.B(n_486),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_829),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_810),
.A2(n_619),
.B(n_602),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_765),
.B(n_665),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_886),
.A2(n_627),
.B(n_599),
.Y(n_937)
);

HB1xp67_ASAP7_75t_L g938 ( 
.A(n_797),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_768),
.A2(n_638),
.B(n_627),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_815),
.A2(n_646),
.B(n_638),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_797),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_747),
.B(n_670),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_785),
.B(n_761),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_802),
.B(n_683),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_765),
.B(n_665),
.Y(n_945)
);

O2A1O1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_793),
.A2(n_662),
.B(n_582),
.C(n_590),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_788),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_802),
.B(n_662),
.Y(n_948)
);

AOI21xp33_ASAP7_75t_L g949 ( 
.A1(n_740),
.A2(n_598),
.B(n_590),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_730),
.A2(n_598),
.B(n_650),
.C(n_652),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_726),
.A2(n_742),
.B(n_833),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_736),
.B(n_638),
.Y(n_952)
);

AOI21x1_ASAP7_75t_L g953 ( 
.A1(n_869),
.A2(n_615),
.B(n_691),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_736),
.A2(n_794),
.B1(n_880),
.B2(n_872),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_737),
.B(n_646),
.Y(n_955)
);

BUFx6f_ASAP7_75t_L g956 ( 
.A(n_735),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_839),
.A2(n_650),
.B(n_646),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_779),
.A2(n_650),
.B(n_652),
.C(n_674),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_840),
.A2(n_674),
.B(n_652),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_798),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_778),
.A2(n_677),
.B(n_674),
.C(n_615),
.Y(n_961)
);

AO21x1_ASAP7_75t_L g962 ( 
.A1(n_873),
.A2(n_656),
.B(n_617),
.Y(n_962)
);

BUFx2_ASAP7_75t_SL g963 ( 
.A(n_765),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_765),
.B(n_665),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_776),
.B(n_488),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_800),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_803),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_783),
.B(n_665),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_878),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_784),
.A2(n_677),
.B(n_656),
.C(n_715),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_853),
.B(n_713),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_SL g972 ( 
.A(n_842),
.B(n_490),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_891),
.B(n_491),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_841),
.A2(n_677),
.B(n_691),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_828),
.A2(n_389),
.B(n_388),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_806),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_846),
.A2(n_702),
.B(n_700),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_817),
.Y(n_978)
);

INVx2_ASAP7_75t_SL g979 ( 
.A(n_829),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_853),
.B(n_713),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_826),
.B(n_665),
.Y(n_981)
);

BUFx4f_ASAP7_75t_L g982 ( 
.A(n_735),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_856),
.A2(n_857),
.B(n_812),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_831),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_783),
.B(n_672),
.Y(n_985)
);

O2A1O1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_887),
.A2(n_723),
.B(n_718),
.C(n_715),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_752),
.A2(n_718),
.B(n_703),
.C(n_702),
.Y(n_987)
);

O2A1O1Ixp5_ASAP7_75t_L g988 ( 
.A1(n_808),
.A2(n_703),
.B(n_700),
.C(n_723),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_770),
.A2(n_676),
.B(n_672),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_836),
.B(n_672),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_858),
.B(n_713),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_822),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_822),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_739),
.A2(n_676),
.B(n_672),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_858),
.B(n_713),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_753),
.B(n_612),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_873),
.A2(n_617),
.B(n_507),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_739),
.A2(n_672),
.B(n_684),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_819),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_814),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_814),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_860),
.B(n_713),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_860),
.B(n_713),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_820),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_863),
.B(n_729),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_863),
.B(n_676),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_746),
.A2(n_684),
.B(n_676),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_792),
.B(n_676),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_746),
.A2(n_684),
.B(n_511),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_814),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_834),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_748),
.A2(n_684),
.B(n_511),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_748),
.A2(n_684),
.B(n_511),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_879),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_823),
.B(n_389),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_874),
.B(n_390),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_845),
.B(n_285),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_814),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_758),
.A2(n_506),
.B(n_507),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_885),
.B(n_888),
.Y(n_1020)
);

AND2x4_ASAP7_75t_SL g1021 ( 
.A(n_801),
.B(n_612),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_781),
.B(n_291),
.Y(n_1022)
);

NOR3xp33_ASAP7_75t_L g1023 ( 
.A(n_828),
.B(n_292),
.C(n_325),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_758),
.A2(n_506),
.B(n_507),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_838),
.B(n_295),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_872),
.B(n_298),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_880),
.A2(n_317),
.B1(n_301),
.B2(n_304),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_831),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_838),
.B(n_312),
.Y(n_1029)
);

BUFx4f_ASAP7_75t_L g1030 ( 
.A(n_727),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_805),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_762),
.A2(n_506),
.B(n_507),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_791),
.A2(n_520),
.B(n_515),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_744),
.B(n_326),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_827),
.B(n_331),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_889),
.B(n_340),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_750),
.B(n_342),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_762),
.A2(n_769),
.B(n_767),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_889),
.B(n_343),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_754),
.B(n_344),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_871),
.A2(n_511),
.B(n_506),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_884),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_884),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_751),
.B(n_346),
.Y(n_1044)
);

OAI321xp33_ASAP7_75t_L g1045 ( 
.A1(n_868),
.A2(n_801),
.A3(n_775),
.B1(n_852),
.B2(n_733),
.C(n_772),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_807),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_786),
.B(n_351),
.Y(n_1047)
);

OAI22x1_ASAP7_75t_L g1048 ( 
.A1(n_831),
.A2(n_391),
.B1(n_354),
.B2(n_352),
.Y(n_1048)
);

AOI22x1_ASAP7_75t_L g1049 ( 
.A1(n_867),
.A2(n_510),
.B1(n_514),
.B2(n_520),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_844),
.B(n_243),
.Y(n_1050)
);

O2A1O1Ixp5_ASAP7_75t_L g1051 ( 
.A1(n_876),
.A2(n_515),
.B(n_520),
.C(n_510),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_868),
.A2(n_515),
.B(n_520),
.C(n_514),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_786),
.B(n_767),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_835),
.A2(n_883),
.B(n_875),
.C(n_859),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_769),
.A2(n_510),
.B(n_514),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_745),
.B(n_612),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_777),
.B(n_250),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_777),
.A2(n_864),
.B(n_861),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_837),
.B(n_849),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_844),
.B(n_612),
.Y(n_1060)
);

AOI33xp33_ASAP7_75t_L g1061 ( 
.A1(n_843),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.B3(n_14),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_862),
.A2(n_515),
.B(n_514),
.C(n_510),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_867),
.A2(n_289),
.B(n_255),
.Y(n_1063)
);

AO21x2_ASAP7_75t_L g1064 ( 
.A1(n_876),
.A2(n_522),
.B(n_529),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_884),
.B(n_890),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_733),
.B(n_262),
.Y(n_1067)
);

CKINVDCx10_ASAP7_75t_R g1068 ( 
.A(n_738),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_787),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_884),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_865),
.B(n_290),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_787),
.A2(n_525),
.B1(n_529),
.B2(n_522),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_866),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_882),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1025),
.B(n_790),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_SL g1076 ( 
.A1(n_973),
.A2(n_319),
.B1(n_265),
.B2(n_269),
.Y(n_1076)
);

OR2x6_ASAP7_75t_L g1077 ( 
.A(n_934),
.B(n_790),
.Y(n_1077)
);

CKINVDCx14_ASAP7_75t_R g1078 ( 
.A(n_911),
.Y(n_1078)
);

OAI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_922),
.A2(n_821),
.B1(n_796),
.B2(n_848),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_954),
.B(n_796),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1025),
.B(n_813),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_943),
.A2(n_918),
.B1(n_1020),
.B2(n_898),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1029),
.B(n_813),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_1029),
.A2(n_855),
.B(n_818),
.C(n_854),
.Y(n_1084)
);

NOR2xp67_ASAP7_75t_L g1085 ( 
.A(n_979),
.B(n_821),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_SL g1086 ( 
.A1(n_906),
.A2(n_848),
.B(n_847),
.C(n_832),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_918),
.B(n_832),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1006),
.A2(n_847),
.B(n_881),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_983),
.A2(n_310),
.B(n_274),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_896),
.B(n_522),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1039),
.B(n_264),
.Y(n_1091)
);

AOI33xp33_ASAP7_75t_L g1092 ( 
.A1(n_1027),
.A2(n_11),
.A3(n_12),
.B1(n_15),
.B2(n_19),
.B3(n_20),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_907),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_907),
.B(n_277),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_915),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1023),
.A2(n_335),
.B1(n_278),
.B2(n_280),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_913),
.A2(n_339),
.B(n_288),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_916),
.B(n_19),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_921),
.B(n_28),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_921),
.B(n_33),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_919),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_522),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_928),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_930),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_1023),
.A2(n_348),
.B1(n_282),
.B2(n_297),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_925),
.Y(n_1106)
);

BUFx4f_ASAP7_75t_L g1107 ( 
.A(n_893),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_947),
.B(n_35),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_935),
.A2(n_306),
.B(n_333),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_926),
.Y(n_1110)
);

AND2x4_ASAP7_75t_L g1111 ( 
.A(n_938),
.B(n_941),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_SL g1112 ( 
.A(n_982),
.B(n_350),
.Y(n_1112)
);

INVx4_ASAP7_75t_L g1113 ( 
.A(n_956),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_951),
.A2(n_338),
.B(n_497),
.Y(n_1114)
);

AND2x6_ASAP7_75t_L g1115 ( 
.A(n_1060),
.B(n_522),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1054),
.A2(n_529),
.B(n_525),
.C(n_522),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_956),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_975),
.A2(n_529),
.B1(n_522),
.B2(n_42),
.C(n_43),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_960),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_956),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_1005),
.A2(n_252),
.B(n_208),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_953),
.A2(n_252),
.B(n_208),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_942),
.A2(n_497),
.B(n_495),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_R g1124 ( 
.A(n_972),
.B(n_112),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_966),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_892),
.A2(n_497),
.B(n_495),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_932),
.A2(n_497),
.B(n_495),
.Y(n_1127)
);

NOR2xp67_ASAP7_75t_L g1128 ( 
.A(n_901),
.B(n_933),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_917),
.A2(n_497),
.B(n_495),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_967),
.Y(n_1130)
);

A2O1A1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_1045),
.A2(n_529),
.B(n_522),
.C(n_497),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_938),
.B(n_941),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_893),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_SL g1134 ( 
.A(n_1030),
.B(n_529),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_899),
.A2(n_904),
.B(n_957),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_959),
.A2(n_497),
.B(n_495),
.Y(n_1136)
);

OR2x6_ASAP7_75t_SL g1137 ( 
.A(n_1074),
.B(n_1068),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1030),
.B(n_529),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_976),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1031),
.B(n_41),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1046),
.B(n_529),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_965),
.B(n_46),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_956),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_978),
.B(n_208),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1035),
.A2(n_252),
.B1(n_208),
.B2(n_498),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_940),
.A2(n_495),
.B(n_497),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_999),
.B(n_208),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_893),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_1004),
.A2(n_1011),
.B1(n_948),
.B2(n_894),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1035),
.A2(n_495),
.B(n_252),
.C(n_51),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_1059),
.B(n_47),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1069),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1028),
.A2(n_48),
.B1(n_53),
.B2(n_54),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1041),
.A2(n_997),
.B(n_962),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_908),
.Y(n_1155)
);

AND2x4_ASAP7_75t_L g1156 ( 
.A(n_931),
.B(n_55),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_894),
.B(n_58),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_944),
.B(n_61),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_923),
.A2(n_61),
.B1(n_65),
.B2(n_67),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1026),
.A2(n_68),
.B(n_252),
.C(n_495),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1022),
.A2(n_252),
.B1(n_84),
.B2(n_88),
.Y(n_1161)
);

AOI22xp5_ASAP7_75t_L g1162 ( 
.A1(n_1071),
.A2(n_252),
.B1(n_498),
.B2(n_91),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_969),
.Y(n_1163)
);

NOR3xp33_ASAP7_75t_L g1164 ( 
.A(n_1036),
.B(n_900),
.C(n_1016),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_902),
.A2(n_78),
.B(n_89),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1000),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_908),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_L g1168 ( 
.A1(n_1048),
.A2(n_498),
.B1(n_103),
.B2(n_108),
.Y(n_1168)
);

BUFx10_ASAP7_75t_L g1169 ( 
.A(n_1071),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1015),
.A2(n_96),
.B1(n_113),
.B2(n_116),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_984),
.A2(n_914),
.B1(n_1073),
.B2(n_927),
.Y(n_1171)
);

BUFx8_ASAP7_75t_L g1172 ( 
.A(n_1056),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_897),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_974),
.A2(n_117),
.B(n_120),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_931),
.B(n_1021),
.Y(n_1175)
);

O2A1O1Ixp5_ASAP7_75t_L g1176 ( 
.A1(n_905),
.A2(n_498),
.B(n_134),
.C(n_135),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_900),
.A2(n_498),
.B(n_143),
.C(n_144),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1017),
.B(n_498),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1000),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1014),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_897),
.B(n_128),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_1034),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_L g1183 ( 
.A(n_1044),
.B(n_152),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_1000),
.Y(n_1184)
);

BUFx12f_ASAP7_75t_L g1185 ( 
.A(n_1000),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_952),
.A2(n_498),
.B(n_162),
.C(n_163),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_992),
.B(n_498),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_929),
.A2(n_159),
.B(n_170),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1065),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1037),
.A2(n_498),
.B(n_179),
.C(n_182),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_993),
.B(n_175),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_1010),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1040),
.B(n_191),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_993),
.B(n_996),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_SL g1195 ( 
.A1(n_950),
.A2(n_945),
.B(n_924),
.C(n_964),
.Y(n_1195)
);

OR2x2_ASAP7_75t_L g1196 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_912),
.A2(n_977),
.B(n_989),
.Y(n_1197)
);

AOI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_952),
.A2(n_996),
.B1(n_981),
.B2(n_990),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1061),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_937),
.A2(n_903),
.B(n_1058),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1066),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_963),
.B(n_955),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_994),
.A2(n_1007),
.B(n_998),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1066),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_955),
.B(n_1060),
.Y(n_1205)
);

A2O1A1Ixp33_ASAP7_75t_L g1206 ( 
.A1(n_946),
.A2(n_990),
.B(n_981),
.C(n_986),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1010),
.B(n_1042),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_958),
.A2(n_895),
.B(n_970),
.C(n_1033),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_1010),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_L g1210 ( 
.A1(n_971),
.A2(n_991),
.B(n_1003),
.C(n_1002),
.Y(n_1210)
);

BUFx2_ASAP7_75t_L g1211 ( 
.A(n_1001),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1008),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1010),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1018),
.B(n_1042),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_949),
.B(n_1057),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1001),
.B(n_1018),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1064),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1018),
.B(n_1042),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_SL g1219 ( 
.A(n_980),
.B(n_995),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1050),
.B(n_1042),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1018),
.B(n_1043),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_SL g1222 ( 
.A1(n_909),
.A2(n_1063),
.B(n_939),
.C(n_987),
.Y(n_1222)
);

CKINVDCx14_ASAP7_75t_R g1223 ( 
.A(n_1043),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1151),
.A2(n_968),
.B(n_985),
.C(n_936),
.Y(n_1224)
);

BUFx12f_ASAP7_75t_L g1225 ( 
.A(n_1095),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1091),
.A2(n_910),
.B(n_920),
.C(n_1062),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1167),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1200),
.A2(n_1043),
.B(n_1070),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1203),
.A2(n_1135),
.B(n_1082),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_SL g1230 ( 
.A1(n_1098),
.A2(n_1052),
.B(n_1067),
.C(n_1009),
.Y(n_1230)
);

INVx3_ASAP7_75t_SL g1231 ( 
.A(n_1110),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1142),
.A2(n_1051),
.B(n_988),
.C(n_961),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1082),
.A2(n_1070),
.B(n_1043),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1078),
.B(n_1070),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1155),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1075),
.A2(n_1051),
.B(n_988),
.C(n_1038),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1199),
.A2(n_1157),
.B1(n_1159),
.B2(n_1108),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1101),
.Y(n_1239)
);

A2O1A1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1193),
.A2(n_961),
.B(n_1012),
.C(n_1013),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1122),
.A2(n_1049),
.B(n_1024),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1116),
.A2(n_1064),
.B(n_1032),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1182),
.B(n_1019),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1206),
.A2(n_1055),
.B(n_1072),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1197),
.A2(n_1072),
.B(n_1081),
.Y(n_1245)
);

AO32x2_ASAP7_75t_L g1246 ( 
.A1(n_1159),
.A2(n_1149),
.A3(n_1079),
.B1(n_1161),
.B2(n_1170),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1121),
.A2(n_1217),
.A3(n_1079),
.B(n_1088),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1093),
.Y(n_1248)
);

OA21x2_ASAP7_75t_L g1249 ( 
.A1(n_1154),
.A2(n_1126),
.B(n_1146),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1111),
.B(n_1132),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1152),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1083),
.A2(n_1222),
.B(n_1208),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1164),
.A2(n_1084),
.B(n_1183),
.C(n_1160),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1129),
.A2(n_1136),
.B(n_1127),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1076),
.B(n_1094),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1123),
.A2(n_1165),
.B(n_1210),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1174),
.A2(n_1188),
.B(n_1114),
.Y(n_1257)
);

AO22x2_ASAP7_75t_L g1258 ( 
.A1(n_1196),
.A2(n_1149),
.B1(n_1215),
.B2(n_1205),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1195),
.A2(n_1219),
.B(n_1080),
.Y(n_1259)
);

AOI211x1_ASAP7_75t_L g1260 ( 
.A1(n_1099),
.A2(n_1100),
.B(n_1140),
.C(n_1103),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1169),
.B(n_1111),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1219),
.A2(n_1202),
.B(n_1086),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_1185),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1205),
.B(n_1115),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1104),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1132),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1117),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1137),
.Y(n_1268)
);

NAND3xp33_ASAP7_75t_L g1269 ( 
.A(n_1118),
.B(n_1092),
.C(n_1105),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1128),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1096),
.A2(n_1156),
.B1(n_1198),
.B2(n_1125),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1153),
.A2(n_1171),
.B1(n_1201),
.B2(n_1106),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1223),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_1162),
.A2(n_1109),
.B(n_1097),
.C(n_1220),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1107),
.Y(n_1275)
);

OAI22x1_ASAP7_75t_L g1276 ( 
.A1(n_1133),
.A2(n_1148),
.B1(n_1156),
.B2(n_1139),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1119),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1090),
.Y(n_1278)
);

OA21x2_ASAP7_75t_L g1279 ( 
.A1(n_1131),
.A2(n_1147),
.B(n_1144),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1144),
.A2(n_1147),
.B(n_1141),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1115),
.B(n_1212),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1113),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1115),
.B(n_1130),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1158),
.A2(n_1168),
.B(n_1089),
.C(n_1145),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1141),
.A2(n_1221),
.B(n_1214),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1218),
.A2(n_1191),
.B(n_1138),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1134),
.A2(n_1207),
.B(n_1216),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1077),
.B(n_1204),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1177),
.A2(n_1190),
.B(n_1186),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1107),
.A2(n_1077),
.B1(n_1211),
.B2(n_1194),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1221),
.A2(n_1102),
.B(n_1176),
.Y(n_1291)
);

O2A1O1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1077),
.A2(n_1173),
.B(n_1187),
.C(n_1112),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1102),
.A2(n_1179),
.B(n_1112),
.Y(n_1293)
);

AO32x2_ASAP7_75t_L g1294 ( 
.A1(n_1209),
.A2(n_1213),
.A3(n_1113),
.B1(n_1169),
.B2(n_1172),
.Y(n_1294)
);

INVxp67_ASAP7_75t_SL g1295 ( 
.A(n_1166),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1179),
.A2(n_1192),
.B(n_1184),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1166),
.A2(n_1192),
.B(n_1184),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1115),
.A2(n_1085),
.B1(n_1175),
.B2(n_1172),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1163),
.A2(n_1180),
.B(n_1189),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1166),
.A2(n_1192),
.B(n_1184),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1209),
.B(n_1213),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_1117),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1178),
.A2(n_1124),
.B(n_1181),
.C(n_1117),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1120),
.A2(n_922),
.B(n_1200),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1120),
.A2(n_984),
.A3(n_1082),
.B1(n_1159),
.B2(n_1149),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1120),
.Y(n_1306)
);

O2A1O1Ixp33_ASAP7_75t_SL g1307 ( 
.A1(n_1143),
.A2(n_922),
.B(n_1098),
.C(n_1005),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1143),
.A2(n_922),
.B(n_1200),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1143),
.B(n_773),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1091),
.A2(n_831),
.B1(n_1048),
.B2(n_804),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1093),
.Y(n_1311)
);

AO21x1_ASAP7_75t_L g1312 ( 
.A1(n_1161),
.A2(n_1082),
.B(n_1091),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1313)
);

OAI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1314)
);

AO21x2_ASAP7_75t_L g1315 ( 
.A1(n_1154),
.A2(n_1217),
.B(n_1200),
.Y(n_1315)
);

BUFx6f_ASAP7_75t_L g1316 ( 
.A(n_1185),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1101),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1091),
.B(n_757),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1093),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1091),
.A2(n_831),
.B1(n_1048),
.B2(n_804),
.Y(n_1321)
);

AO22x1_ASAP7_75t_L g1322 ( 
.A1(n_1091),
.A2(n_973),
.B1(n_829),
.B2(n_1039),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1324)
);

AO21x1_ASAP7_75t_L g1325 ( 
.A1(n_1161),
.A2(n_1082),
.B(n_1091),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1091),
.B(n_757),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1082),
.B(n_757),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1154),
.A2(n_1135),
.B(n_1197),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1078),
.Y(n_1331)
);

AOI31xp67_ASAP7_75t_L g1332 ( 
.A1(n_1080),
.A2(n_1217),
.A3(n_905),
.B(n_1198),
.Y(n_1332)
);

A2O1A1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1091),
.A2(n_1025),
.B(n_1029),
.C(n_1039),
.Y(n_1333)
);

AOI221x1_ASAP7_75t_L g1334 ( 
.A1(n_1161),
.A2(n_1048),
.B1(n_1150),
.B2(n_1151),
.C(n_1159),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1107),
.B(n_1175),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1151),
.A2(n_922),
.B1(n_954),
.B2(n_918),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1101),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1091),
.B(n_757),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1200),
.A2(n_1197),
.B(n_1122),
.Y(n_1342)
);

AO21x1_ASAP7_75t_L g1343 ( 
.A1(n_1161),
.A2(n_1082),
.B(n_1091),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1121),
.A2(n_1217),
.A3(n_997),
.B(n_962),
.Y(n_1348)
);

OAI21xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1151),
.A2(n_1029),
.B(n_1025),
.Y(n_1349)
);

A2O1A1Ixp33_ASAP7_75t_L g1350 ( 
.A1(n_1091),
.A2(n_1025),
.B(n_1029),
.C(n_1039),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1185),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1154),
.A2(n_1135),
.B(n_1197),
.Y(n_1353)
);

BUFx12f_ASAP7_75t_L g1354 ( 
.A(n_1095),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1356)
);

AO31x2_ASAP7_75t_L g1357 ( 
.A1(n_1121),
.A2(n_1217),
.A3(n_997),
.B(n_962),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1151),
.A2(n_1029),
.B(n_1025),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1359)
);

OAI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_1095),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1091),
.B(n_1029),
.C(n_1025),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1363)
);

INVx4_ASAP7_75t_SL g1364 ( 
.A(n_1115),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1121),
.A2(n_1217),
.A3(n_997),
.B(n_962),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1206),
.A2(n_922),
.B(n_1082),
.Y(n_1366)
);

OA21x2_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_1197),
.B(n_1122),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1101),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1095),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1101),
.Y(n_1370)
);

O2A1O1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1151),
.A2(n_1025),
.B(n_1029),
.C(n_757),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1082),
.B(n_757),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1122),
.A2(n_1197),
.B(n_1203),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1082),
.B(n_1087),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1091),
.B(n_757),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_1095),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1200),
.A2(n_922),
.B(n_1006),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1091),
.B(n_757),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1082),
.B(n_757),
.Y(n_1379)
);

AO31x2_ASAP7_75t_L g1380 ( 
.A1(n_1121),
.A2(n_1217),
.A3(n_997),
.B(n_962),
.Y(n_1380)
);

INVx3_ASAP7_75t_SL g1381 ( 
.A(n_1231),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1310),
.A2(n_1321),
.B1(n_1362),
.B2(n_1337),
.Y(n_1382)
);

BUFx4f_ASAP7_75t_SL g1383 ( 
.A(n_1225),
.Y(n_1383)
);

INVx6_ASAP7_75t_L g1384 ( 
.A(n_1316),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1265),
.Y(n_1385)
);

CKINVDCx11_ASAP7_75t_R g1386 ( 
.A(n_1376),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1277),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1315),
.Y(n_1388)
);

BUFx12f_ASAP7_75t_L g1389 ( 
.A(n_1361),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1333),
.A2(n_1350),
.B(n_1349),
.Y(n_1390)
);

BUFx4_ASAP7_75t_SL g1391 ( 
.A(n_1227),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1238),
.A2(n_1269),
.B1(n_1255),
.B2(n_1343),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1329),
.B(n_1372),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1379),
.B(n_1318),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1317),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1312),
.A2(n_1325),
.B1(n_1347),
.B2(n_1326),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1334),
.B2(n_1360),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1250),
.B(n_1266),
.Y(n_1398)
);

AOI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1358),
.A2(n_1341),
.B1(n_1378),
.B2(n_1328),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1375),
.B(n_1320),
.Y(n_1400)
);

CKINVDCx14_ASAP7_75t_R g1401 ( 
.A(n_1331),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1326),
.A2(n_1360),
.B1(n_1366),
.B2(n_1347),
.Y(n_1402)
);

BUFx4_ASAP7_75t_SL g1403 ( 
.A(n_1263),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1371),
.B(n_1311),
.Y(n_1404)
);

CKINVDCx14_ASAP7_75t_R g1405 ( 
.A(n_1354),
.Y(n_1405)
);

CKINVDCx6p67_ASAP7_75t_R g1406 ( 
.A(n_1369),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1344),
.A2(n_1366),
.B1(n_1355),
.B2(n_1323),
.Y(n_1407)
);

CKINVDCx11_ASAP7_75t_R g1408 ( 
.A(n_1361),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1344),
.A2(n_1355),
.B(n_1253),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1340),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1271),
.A2(n_1323),
.B1(n_1327),
.B2(n_1319),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1267),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1268),
.Y(n_1413)
);

BUFx4f_ASAP7_75t_SL g1414 ( 
.A(n_1316),
.Y(n_1414)
);

BUFx12f_ASAP7_75t_L g1415 ( 
.A(n_1316),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1271),
.A2(n_1319),
.B1(n_1345),
.B2(n_1374),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1327),
.A2(n_1374),
.B1(n_1345),
.B2(n_1260),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1294),
.Y(n_1418)
);

BUFx2_ASAP7_75t_SL g1419 ( 
.A(n_1273),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1258),
.A2(n_1272),
.B1(n_1276),
.B2(n_1370),
.Y(n_1420)
);

BUFx12f_ASAP7_75t_L g1421 ( 
.A(n_1236),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1267),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1267),
.Y(n_1423)
);

INVx6_ASAP7_75t_L g1424 ( 
.A(n_1302),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1258),
.A2(n_1305),
.B1(n_1290),
.B2(n_1246),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1368),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1235),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1351),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1270),
.A2(n_1309),
.B1(n_1278),
.B2(n_1290),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_SL g1430 ( 
.A1(n_1298),
.A2(n_1274),
.B(n_1259),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_SL g1431 ( 
.A1(n_1305),
.A2(n_1246),
.B1(n_1322),
.B2(n_1279),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1251),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1351),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1243),
.A2(n_1288),
.B1(n_1279),
.B2(n_1244),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1299),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1244),
.A2(n_1264),
.B1(n_1261),
.B2(n_1283),
.Y(n_1436)
);

CKINVDCx11_ASAP7_75t_R g1437 ( 
.A(n_1364),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1234),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1264),
.A2(n_1283),
.B1(n_1234),
.B2(n_1305),
.Y(n_1439)
);

OAI22xp5_ASAP7_75t_L g1440 ( 
.A1(n_1284),
.A2(n_1252),
.B1(n_1229),
.B2(n_1224),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1246),
.A2(n_1335),
.B1(n_1275),
.B2(n_1281),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1335),
.A2(n_1245),
.B1(n_1364),
.B2(n_1280),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1294),
.B(n_1306),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1306),
.B(n_1295),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1364),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1304),
.A2(n_1308),
.B1(n_1233),
.B2(n_1282),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1313),
.A2(n_1346),
.B1(n_1352),
.B2(n_1336),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1289),
.A2(n_1226),
.B1(n_1293),
.B2(n_1262),
.Y(n_1448)
);

CKINVDCx11_ASAP7_75t_R g1449 ( 
.A(n_1294),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1292),
.Y(n_1450)
);

BUFx12f_ASAP7_75t_L g1451 ( 
.A(n_1303),
.Y(n_1451)
);

BUFx4f_ASAP7_75t_SL g1452 ( 
.A(n_1307),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1286),
.A2(n_1377),
.B(n_1363),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1285),
.B(n_1301),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1332),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1301),
.A2(n_1287),
.B1(n_1296),
.B2(n_1291),
.Y(n_1456)
);

OAI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1240),
.A2(n_1232),
.B1(n_1237),
.B2(n_1228),
.Y(n_1457)
);

BUFx8_ASAP7_75t_L g1458 ( 
.A(n_1297),
.Y(n_1458)
);

OAI21xp5_ASAP7_75t_SL g1459 ( 
.A1(n_1300),
.A2(n_1242),
.B(n_1330),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1315),
.B(n_1247),
.Y(n_1460)
);

CKINVDCx20_ASAP7_75t_R g1461 ( 
.A(n_1249),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1257),
.A2(n_1256),
.B1(n_1342),
.B2(n_1367),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1342),
.A2(n_1367),
.B1(n_1254),
.B2(n_1241),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1247),
.B(n_1348),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1247),
.B(n_1380),
.Y(n_1465)
);

OAI21xp33_ASAP7_75t_L g1466 ( 
.A1(n_1353),
.A2(n_1339),
.B(n_1314),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1324),
.A2(n_1338),
.B1(n_1373),
.B2(n_1359),
.Y(n_1467)
);

OAI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1230),
.A2(n_1356),
.B1(n_1380),
.B2(n_1357),
.Y(n_1468)
);

INVx6_ASAP7_75t_L g1469 ( 
.A(n_1357),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1357),
.A2(n_1349),
.B1(n_1358),
.B2(n_1362),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1365),
.A2(n_1380),
.B1(n_1048),
.B2(n_1310),
.Y(n_1471)
);

BUFx12f_ASAP7_75t_L g1472 ( 
.A(n_1365),
.Y(n_1472)
);

INVx3_ASAP7_75t_SL g1473 ( 
.A(n_1231),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1329),
.B(n_1372),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1225),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1267),
.Y(n_1476)
);

CKINVDCx11_ASAP7_75t_R g1477 ( 
.A(n_1376),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1239),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1231),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1349),
.A2(n_1358),
.B(n_1362),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1248),
.Y(n_1481)
);

INVx6_ASAP7_75t_L g1482 ( 
.A(n_1316),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1329),
.B(n_1372),
.Y(n_1483)
);

INVx4_ASAP7_75t_L g1484 ( 
.A(n_1316),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1310),
.A2(n_1048),
.B1(n_1321),
.B2(n_804),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1239),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1337),
.A2(n_671),
.B1(n_831),
.B2(n_801),
.Y(n_1487)
);

OAI22xp33_ASAP7_75t_L g1488 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1337),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1337),
.A2(n_801),
.B1(n_891),
.B2(n_1137),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1350),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1337),
.A2(n_671),
.B1(n_831),
.B2(n_801),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1316),
.Y(n_1492)
);

CKINVDCx6p67_ASAP7_75t_R g1493 ( 
.A(n_1225),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1350),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1337),
.A2(n_671),
.B1(n_831),
.B2(n_801),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1329),
.B(n_1372),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1239),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1248),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1350),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_SL g1500 ( 
.A1(n_1337),
.A2(n_671),
.B1(n_831),
.B2(n_801),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1376),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1239),
.Y(n_1502)
);

BUFx2_ASAP7_75t_SL g1503 ( 
.A(n_1376),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1239),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1239),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1310),
.A2(n_1048),
.B1(n_1321),
.B2(n_804),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1310),
.A2(n_1048),
.B1(n_1321),
.B2(n_804),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1225),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1310),
.A2(n_1048),
.B1(n_1321),
.B2(n_804),
.Y(n_1509)
);

OAI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1337),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1239),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1350),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_SL g1513 ( 
.A1(n_1255),
.A2(n_1328),
.B1(n_1341),
.B2(n_1318),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1349),
.A2(n_1358),
.B1(n_1362),
.B2(n_1350),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1310),
.A2(n_1048),
.B1(n_1321),
.B2(n_804),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1425),
.B(n_1402),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1438),
.Y(n_1517)
);

AO21x2_ASAP7_75t_L g1518 ( 
.A1(n_1460),
.A2(n_1465),
.B(n_1464),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1453),
.A2(n_1462),
.B(n_1463),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1389),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1404),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1425),
.B(n_1402),
.Y(n_1522)
);

OAI21x1_ASAP7_75t_L g1523 ( 
.A1(n_1462),
.A2(n_1463),
.B(n_1457),
.Y(n_1523)
);

OAI21x1_ASAP7_75t_L g1524 ( 
.A1(n_1468),
.A2(n_1467),
.B(n_1447),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1393),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1435),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1385),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1467),
.A2(n_1447),
.B(n_1440),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1474),
.B(n_1483),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1443),
.B(n_1387),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1417),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1472),
.B(n_1430),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1454),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1400),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1388),
.Y(n_1535)
);

INVx4_ASAP7_75t_SL g1536 ( 
.A(n_1452),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1395),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1454),
.Y(n_1538)
);

BUFx6f_ASAP7_75t_L g1539 ( 
.A(n_1437),
.Y(n_1539)
);

INVx4_ASAP7_75t_L g1540 ( 
.A(n_1452),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1410),
.Y(n_1541)
);

INVx4_ASAP7_75t_SL g1542 ( 
.A(n_1469),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1496),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1426),
.Y(n_1544)
);

AND2x6_ASAP7_75t_L g1545 ( 
.A(n_1450),
.B(n_1456),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1478),
.B(n_1486),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1497),
.Y(n_1547)
);

BUFx2_ASAP7_75t_R g1548 ( 
.A(n_1503),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1484),
.B(n_1492),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1461),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1504),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1505),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1466),
.A2(n_1459),
.B(n_1390),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1446),
.A2(n_1448),
.B(n_1455),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1394),
.B(n_1409),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1411),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1416),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1439),
.Y(n_1559)
);

BUFx3_ASAP7_75t_L g1560 ( 
.A(n_1422),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1418),
.B(n_1396),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1396),
.B(n_1436),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1407),
.B(n_1399),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1436),
.B(n_1434),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1434),
.B(n_1431),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1424),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1439),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1431),
.B(n_1470),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1445),
.Y(n_1569)
);

BUFx2_ASAP7_75t_SL g1570 ( 
.A(n_1432),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1480),
.B(n_1392),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1487),
.A2(n_1491),
.B1(n_1500),
.B2(n_1495),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_SL g1573 ( 
.A1(n_1489),
.A2(n_1499),
.B1(n_1494),
.B2(n_1514),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1424),
.Y(n_1574)
);

AO21x2_ASAP7_75t_L g1575 ( 
.A1(n_1397),
.A2(n_1510),
.B(n_1488),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1391),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1441),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1441),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1481),
.Y(n_1579)
);

INVx2_ASAP7_75t_SL g1580 ( 
.A(n_1498),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_SL g1581 ( 
.A(n_1479),
.Y(n_1581)
);

BUFx6f_ASAP7_75t_L g1582 ( 
.A(n_1451),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1444),
.Y(n_1583)
);

OAI21x1_ASAP7_75t_L g1584 ( 
.A1(n_1442),
.A2(n_1490),
.B(n_1512),
.Y(n_1584)
);

OAI21x1_ASAP7_75t_L g1585 ( 
.A1(n_1471),
.A2(n_1382),
.B(n_1429),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1423),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1398),
.B(n_1449),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1382),
.B(n_1513),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1485),
.A2(n_1515),
.B(n_1509),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1471),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1420),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1412),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1420),
.B(n_1476),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1423),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1427),
.B(n_1491),
.Y(n_1595)
);

OAI21x1_ASAP7_75t_L g1596 ( 
.A1(n_1485),
.A2(n_1515),
.B(n_1509),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1458),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1487),
.A2(n_1495),
.B1(n_1500),
.B2(n_1506),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1421),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1384),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1482),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1428),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1433),
.Y(n_1603)
);

INVx4_ASAP7_75t_L g1604 ( 
.A(n_1482),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1419),
.B(n_1507),
.Y(n_1605)
);

AO21x2_ASAP7_75t_L g1606 ( 
.A1(n_1506),
.A2(n_1507),
.B(n_1492),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1414),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1414),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1381),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1391),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1401),
.B(n_1473),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1415),
.Y(n_1612)
);

AO21x2_ASAP7_75t_L g1613 ( 
.A1(n_1589),
.A2(n_1403),
.B(n_1413),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1550),
.B(n_1405),
.Y(n_1614)
);

AO32x1_ASAP7_75t_L g1615 ( 
.A1(n_1598),
.A2(n_1403),
.A3(n_1408),
.B1(n_1386),
.B2(n_1477),
.Y(n_1615)
);

AO32x2_ASAP7_75t_L g1616 ( 
.A1(n_1580),
.A2(n_1406),
.A3(n_1493),
.B1(n_1383),
.B2(n_1501),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1550),
.B(n_1475),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1530),
.B(n_1508),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1525),
.B(n_1543),
.Y(n_1619)
);

CKINVDCx14_ASAP7_75t_R g1620 ( 
.A(n_1576),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1530),
.B(n_1587),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1521),
.Y(n_1622)
);

A2O1A1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1596),
.A2(n_1588),
.B(n_1563),
.C(n_1562),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1537),
.Y(n_1624)
);

AO32x2_ASAP7_75t_L g1625 ( 
.A1(n_1580),
.A2(n_1538),
.A3(n_1533),
.B1(n_1566),
.B2(n_1574),
.Y(n_1625)
);

OAI22xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1573),
.A2(n_1571),
.B1(n_1555),
.B2(n_1576),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1546),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1579),
.B(n_1551),
.Y(n_1628)
);

INVx4_ASAP7_75t_L g1629 ( 
.A(n_1536),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1557),
.B(n_1558),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1540),
.B(n_1581),
.Y(n_1631)
);

OAI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1605),
.A2(n_1562),
.B1(n_1568),
.B2(n_1572),
.C(n_1516),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1551),
.B(n_1583),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_SL g1634 ( 
.A(n_1545),
.B(n_1532),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1570),
.B(n_1561),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1575),
.A2(n_1557),
.B(n_1558),
.C(n_1605),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1584),
.A2(n_1523),
.B(n_1554),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1537),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1539),
.A2(n_1569),
.B1(n_1540),
.B2(n_1610),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1529),
.B(n_1531),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1609),
.B(n_1611),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1540),
.B(n_1548),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1611),
.B(n_1564),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_L g1644 ( 
.A1(n_1522),
.A2(n_1565),
.B(n_1585),
.C(n_1559),
.Y(n_1644)
);

AOI211xp5_ASAP7_75t_L g1645 ( 
.A1(n_1565),
.A2(n_1595),
.B(n_1567),
.C(n_1559),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1592),
.Y(n_1646)
);

OAI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1545),
.A2(n_1528),
.B(n_1585),
.Y(n_1647)
);

O2A1O1Ixp5_ASAP7_75t_L g1648 ( 
.A1(n_1602),
.A2(n_1603),
.B(n_1600),
.C(n_1601),
.Y(n_1648)
);

BUFx3_ASAP7_75t_L g1649 ( 
.A(n_1599),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1539),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1545),
.B(n_1575),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1527),
.B(n_1534),
.Y(n_1652)
);

AND2x4_ASAP7_75t_SL g1653 ( 
.A(n_1539),
.B(n_1569),
.Y(n_1653)
);

CKINVDCx8_ASAP7_75t_R g1654 ( 
.A(n_1539),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1542),
.B(n_1597),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1577),
.A2(n_1578),
.B(n_1591),
.C(n_1528),
.Y(n_1656)
);

OAI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1591),
.A2(n_1569),
.B1(n_1541),
.B2(n_1556),
.Y(n_1657)
);

CKINVDCx11_ASAP7_75t_R g1658 ( 
.A(n_1569),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1544),
.B(n_1547),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1590),
.A2(n_1606),
.B1(n_1556),
.B2(n_1544),
.C(n_1547),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1545),
.B(n_1517),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1552),
.A2(n_1607),
.B1(n_1608),
.B2(n_1517),
.Y(n_1662)
);

A2O1A1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1593),
.A2(n_1523),
.B(n_1554),
.C(n_1524),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1545),
.A2(n_1524),
.B(n_1519),
.Y(n_1664)
);

CKINVDCx6p67_ASAP7_75t_R g1665 ( 
.A(n_1599),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1593),
.A2(n_1519),
.B(n_1582),
.C(n_1607),
.Y(n_1666)
);

AO32x2_ASAP7_75t_L g1667 ( 
.A1(n_1533),
.A2(n_1538),
.A3(n_1594),
.B1(n_1586),
.B2(n_1604),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1535),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1664),
.B(n_1553),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1664),
.B(n_1553),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1624),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1637),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1630),
.B(n_1553),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1643),
.B(n_1553),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1628),
.B(n_1627),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1668),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1630),
.B(n_1535),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1636),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1625),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1526),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1625),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1647),
.B(n_1651),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1518),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1659),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1625),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1667),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1667),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1667),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1646),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1661),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1662),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1641),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1613),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1676),
.B(n_1635),
.Y(n_1697)
);

AOI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1680),
.A2(n_1632),
.B1(n_1626),
.B2(n_1623),
.C(n_1645),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1680),
.B(n_1622),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1671),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1671),
.Y(n_1701)
);

INVx3_ASAP7_75t_L g1702 ( 
.A(n_1671),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1669),
.A2(n_1634),
.B(n_1615),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1691),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1676),
.B(n_1621),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1680),
.B(n_1619),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_SL g1707 ( 
.A(n_1693),
.B(n_1639),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1669),
.A2(n_1615),
.B(n_1642),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1693),
.B(n_1679),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1695),
.B(n_1629),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1669),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1670),
.B(n_1633),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1693),
.B(n_1652),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1670),
.B(n_1655),
.Y(n_1714)
);

OAI31xp33_ASAP7_75t_L g1715 ( 
.A1(n_1670),
.A2(n_1632),
.A3(n_1644),
.B(n_1657),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1682),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1673),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1679),
.B(n_1660),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1682),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1672),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1672),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1672),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1694),
.B(n_1666),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1694),
.B(n_1656),
.Y(n_1724)
);

INVx2_ASAP7_75t_SL g1725 ( 
.A(n_1688),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1675),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1682),
.Y(n_1727)
);

HB1xp67_ASAP7_75t_L g1728 ( 
.A(n_1673),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1679),
.B(n_1660),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1718),
.B(n_1678),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1702),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1702),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1720),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1718),
.B(n_1678),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1706),
.B(n_1674),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1720),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1706),
.B(n_1674),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1699),
.B(n_1674),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1699),
.B(n_1520),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1714),
.B(n_1692),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1709),
.B(n_1686),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1692),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1709),
.B(n_1686),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1721),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1695),
.Y(n_1749)
);

OR2x6_ASAP7_75t_L g1750 ( 
.A(n_1703),
.B(n_1696),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1729),
.B(n_1695),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1721),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1686),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1722),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1710),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1713),
.B(n_1724),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1705),
.B(n_1692),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1722),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1723),
.B(n_1696),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1724),
.B(n_1681),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1705),
.B(n_1688),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1726),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1712),
.B(n_1688),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1688),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1726),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1731),
.B(n_1725),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1731),
.B(n_1711),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1734),
.Y(n_1771)
);

INVx2_ASAP7_75t_SL g1772 ( 
.A(n_1756),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1757),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1749),
.B(n_1751),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1739),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1737),
.B(n_1711),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1739),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1712),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1748),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1748),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1752),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1755),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1737),
.B(n_1711),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1732),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1738),
.B(n_1697),
.Y(n_1785)
);

AND2x4_ASAP7_75t_SL g1786 ( 
.A(n_1742),
.B(n_1614),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1743),
.B(n_1697),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1757),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1743),
.B(n_1697),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1751),
.B(n_1707),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1732),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_L g1792 ( 
.A(n_1756),
.B(n_1708),
.Y(n_1792)
);

OR2x2_ASAP7_75t_L g1793 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1730),
.B(n_1695),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1732),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1759),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1735),
.B(n_1695),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1735),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1764),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1767),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1767),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1753),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1741),
.B(n_1704),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1733),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1741),
.B(n_1704),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1745),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1746),
.B(n_1681),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1792),
.B(n_1744),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1785),
.B(n_1744),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1774),
.B(n_1745),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1790),
.B(n_1746),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1785),
.B(n_1763),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1773),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1798),
.B(n_1788),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1770),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1802),
.B(n_1758),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1787),
.B(n_1763),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1806),
.B(n_1758),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1787),
.B(n_1765),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1789),
.B(n_1769),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1770),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1806),
.B(n_1747),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1786),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1771),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1771),
.Y(n_1825)
);

OAI222xp33_ASAP7_75t_L g1826 ( 
.A1(n_1794),
.A2(n_1750),
.B1(n_1762),
.B2(n_1703),
.C1(n_1754),
.C2(n_1761),
.Y(n_1826)
);

OAI21xp5_ASAP7_75t_SL g1827 ( 
.A1(n_1797),
.A2(n_1708),
.B(n_1698),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1778),
.B(n_1681),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1772),
.B(n_1681),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1775),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1775),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1793),
.B(n_1747),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1786),
.B(n_1620),
.Y(n_1833)
);

AND2x2_ASAP7_75t_L g1834 ( 
.A(n_1789),
.B(n_1765),
.Y(n_1834)
);

OR2x2_ASAP7_75t_L g1835 ( 
.A(n_1793),
.B(n_1736),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1807),
.B(n_1736),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1777),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1772),
.B(n_1681),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1769),
.B(n_1766),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1777),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1779),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1803),
.B(n_1683),
.Y(n_1842)
);

NOR2x1_ASAP7_75t_L g1843 ( 
.A(n_1779),
.B(n_1649),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1776),
.B(n_1754),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1776),
.B(n_1766),
.Y(n_1845)
);

OAI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1827),
.A2(n_1823),
.B1(n_1750),
.B2(n_1820),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1813),
.B(n_1683),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1821),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1821),
.Y(n_1849)
);

OAI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1820),
.A2(n_1750),
.B1(n_1698),
.B2(n_1687),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1826),
.A2(n_1750),
.B(n_1615),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1840),
.Y(n_1852)
);

OAI221xp5_ASAP7_75t_L g1853 ( 
.A1(n_1842),
.A2(n_1750),
.B1(n_1762),
.B2(n_1715),
.C(n_1725),
.Y(n_1853)
);

AOI32xp33_ASAP7_75t_L g1854 ( 
.A1(n_1808),
.A2(n_1761),
.A3(n_1754),
.B1(n_1760),
.B2(n_1814),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1820),
.B(n_1783),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1808),
.A2(n_1715),
.B1(n_1760),
.B2(n_1761),
.Y(n_1856)
);

OAI22xp5_ASAP7_75t_L g1857 ( 
.A1(n_1844),
.A2(n_1687),
.B1(n_1683),
.B2(n_1719),
.Y(n_1857)
);

INVxp67_ASAP7_75t_SL g1858 ( 
.A(n_1829),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1840),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1844),
.B(n_1783),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1844),
.A2(n_1683),
.B1(n_1687),
.B2(n_1719),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1811),
.B(n_1683),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1843),
.A2(n_1687),
.B1(n_1727),
.B2(n_1719),
.Y(n_1863)
);

AOI222xp33_ASAP7_75t_L g1864 ( 
.A1(n_1838),
.A2(n_1685),
.B1(n_1828),
.B2(n_1754),
.C1(n_1761),
.C2(n_1760),
.Y(n_1864)
);

AOI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1812),
.A2(n_1760),
.B1(n_1685),
.B2(n_1613),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1815),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1833),
.B(n_1710),
.Y(n_1867)
);

INVxp67_ASAP7_75t_L g1868 ( 
.A(n_1824),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1825),
.Y(n_1869)
);

INVx2_ASAP7_75t_SL g1870 ( 
.A(n_1822),
.Y(n_1870)
);

AOI21xp33_ASAP7_75t_L g1871 ( 
.A1(n_1830),
.A2(n_1728),
.B(n_1717),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1812),
.B(n_1687),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1848),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1870),
.B(n_1855),
.Y(n_1874)
);

XNOR2x1_ASAP7_75t_L g1875 ( 
.A(n_1850),
.B(n_1582),
.Y(n_1875)
);

OAI22xp33_ASAP7_75t_L g1876 ( 
.A1(n_1853),
.A2(n_1696),
.B1(n_1690),
.B2(n_1688),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1846),
.B(n_1810),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1867),
.B(n_1810),
.Y(n_1878)
);

AOI211xp5_ASAP7_75t_L g1879 ( 
.A1(n_1851),
.A2(n_1871),
.B(n_1863),
.C(n_1858),
.Y(n_1879)
);

AOI21xp33_ASAP7_75t_L g1880 ( 
.A1(n_1858),
.A2(n_1837),
.B(n_1831),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1860),
.B(n_1817),
.Y(n_1881)
);

OAI221xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1856),
.A2(n_1835),
.B1(n_1832),
.B2(n_1836),
.C(n_1822),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1849),
.Y(n_1883)
);

AOI21xp33_ASAP7_75t_L g1884 ( 
.A1(n_1868),
.A2(n_1841),
.B(n_1728),
.Y(n_1884)
);

OAI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1865),
.A2(n_1690),
.B1(n_1689),
.B2(n_1835),
.Y(n_1885)
);

NAND3xp33_ASAP7_75t_SL g1886 ( 
.A(n_1856),
.B(n_1816),
.C(n_1832),
.Y(n_1886)
);

OAI322xp33_ASAP7_75t_L g1887 ( 
.A1(n_1868),
.A2(n_1836),
.A3(n_1818),
.B1(n_1805),
.B2(n_1717),
.C1(n_1740),
.C2(n_1689),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1866),
.B(n_1817),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1852),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1869),
.B(n_1819),
.Y(n_1890)
);

AOI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1857),
.A2(n_1690),
.B1(n_1689),
.B2(n_1673),
.C(n_1701),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1859),
.Y(n_1892)
);

AOI221xp5_ASAP7_75t_L g1893 ( 
.A1(n_1861),
.A2(n_1690),
.B1(n_1689),
.B2(n_1700),
.C(n_1701),
.Y(n_1893)
);

OAI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1882),
.A2(n_1847),
.B1(n_1862),
.B2(n_1872),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1881),
.B(n_1819),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1888),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_1874),
.B(n_1665),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1890),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1886),
.B(n_1834),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1892),
.B(n_1834),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1878),
.B(n_1839),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1873),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1883),
.Y(n_1903)
);

AOI322xp5_ASAP7_75t_L g1904 ( 
.A1(n_1885),
.A2(n_1845),
.A3(n_1839),
.B1(n_1690),
.B2(n_1689),
.C1(n_1685),
.C2(n_1684),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1889),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1900),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1899),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1897),
.Y(n_1908)
);

AND2x4_ASAP7_75t_L g1909 ( 
.A(n_1902),
.B(n_1877),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1901),
.B(n_1887),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1900),
.Y(n_1911)
);

INVx1_ASAP7_75t_SL g1912 ( 
.A(n_1895),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1903),
.Y(n_1913)
);

OA211x2_ASAP7_75t_L g1914 ( 
.A1(n_1894),
.A2(n_1891),
.B(n_1893),
.C(n_1631),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1896),
.B(n_1880),
.Y(n_1915)
);

OAI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1904),
.A2(n_1879),
.B1(n_1875),
.B2(n_1854),
.C(n_1884),
.Y(n_1916)
);

OAI211xp5_ASAP7_75t_L g1917 ( 
.A1(n_1907),
.A2(n_1910),
.B(n_1916),
.C(n_1915),
.Y(n_1917)
);

AOI222xp33_ASAP7_75t_L g1918 ( 
.A1(n_1907),
.A2(n_1909),
.B1(n_1911),
.B2(n_1876),
.C1(n_1906),
.C2(n_1913),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1909),
.A2(n_1884),
.B1(n_1905),
.B2(n_1898),
.C(n_1700),
.Y(n_1919)
);

NOR2x1_ASAP7_75t_L g1920 ( 
.A(n_1912),
.B(n_1612),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1908),
.A2(n_1864),
.B(n_1781),
.Y(n_1921)
);

XOR2x2_ASAP7_75t_L g1922 ( 
.A(n_1914),
.B(n_1617),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1909),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1919),
.A2(n_1845),
.B1(n_1784),
.B2(n_1804),
.C(n_1791),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_SL g1925 ( 
.A(n_1923),
.B(n_1917),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1918),
.A2(n_1781),
.B(n_1780),
.Y(n_1926)
);

AOI221xp5_ASAP7_75t_L g1927 ( 
.A1(n_1921),
.A2(n_1701),
.B1(n_1700),
.B2(n_1795),
.C(n_1784),
.Y(n_1927)
);

O2A1O1Ixp33_ASAP7_75t_L g1928 ( 
.A1(n_1920),
.A2(n_1791),
.B(n_1804),
.C(n_1795),
.Y(n_1928)
);

NOR2xp67_ASAP7_75t_L g1929 ( 
.A(n_1922),
.B(n_1780),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1917),
.A2(n_1796),
.B1(n_1782),
.B2(n_1801),
.C(n_1800),
.Y(n_1930)
);

NOR3xp33_ASAP7_75t_L g1931 ( 
.A(n_1917),
.B(n_1612),
.C(n_1658),
.Y(n_1931)
);

AND2x2_ASAP7_75t_SL g1932 ( 
.A(n_1931),
.B(n_1925),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1929),
.B(n_1926),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1924),
.B(n_1809),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1930),
.B(n_1809),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1927),
.B(n_1768),
.Y(n_1936)
);

XOR2xp5_ASAP7_75t_L g1937 ( 
.A(n_1928),
.B(n_1612),
.Y(n_1937)
);

NOR4xp75_ASAP7_75t_L g1938 ( 
.A(n_1934),
.B(n_1616),
.C(n_1650),
.D(n_1618),
.Y(n_1938)
);

OAI211xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1933),
.A2(n_1616),
.B(n_1608),
.C(n_1654),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1935),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1932),
.Y(n_1941)
);

NOR4xp25_ASAP7_75t_L g1942 ( 
.A(n_1941),
.B(n_1932),
.C(n_1936),
.D(n_1937),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1942),
.Y(n_1943)
);

XOR2x2_ASAP7_75t_L g1944 ( 
.A(n_1943),
.B(n_1940),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1943),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1945),
.B(n_1935),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1944),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1946),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1947),
.Y(n_1949)
);

AOI21xp5_ASAP7_75t_L g1950 ( 
.A1(n_1949),
.A2(n_1939),
.B(n_1938),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1950),
.A2(n_1948),
.B(n_1653),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1951),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1952),
.A2(n_1782),
.B1(n_1801),
.B2(n_1800),
.C(n_1799),
.Y(n_1953)
);

AOI211xp5_ASAP7_75t_L g1954 ( 
.A1(n_1953),
.A2(n_1560),
.B(n_1616),
.C(n_1549),
.Y(n_1954)
);


endmodule