module fake_jpeg_8761_n_115 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_115);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_115;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_17),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_9),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_10),
.B1(n_18),
.B2(n_11),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_28),
.B1(n_31),
.B2(n_25),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_22),
.B1(n_20),
.B2(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_18),
.B1(n_16),
.B2(n_9),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_19),
.B(n_21),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_32),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_37),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_45),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_22),
.B(n_20),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_16),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_12),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_54),
.B1(n_58),
.B2(n_56),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_20),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g63 ( 
.A1(n_51),
.A2(n_41),
.B(n_22),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_51),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_62),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_60),
.A2(n_28),
.B1(n_33),
.B2(n_50),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_65),
.B(n_66),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_36),
.C(n_19),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_52),
.C(n_51),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_28),
.B(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_75),
.C(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_77),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_67),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_28),
.Y(n_78)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_26),
.C(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_67),
.Y(n_81)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_64),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_63),
.C(n_61),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_84),
.B(n_85),
.C(n_88),
.Y(n_92)
);

AOI221xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_13),
.B1(n_80),
.B2(n_3),
.C(n_4),
.Y(n_91)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_26),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_83),
.A2(n_73),
.B1(n_78),
.B2(n_79),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_95),
.B1(n_33),
.B2(n_26),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_91),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_84),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_100),
.C(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_33),
.B(n_1),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_99),
.A2(n_13),
.B(n_91),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_7),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_103),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_104),
.B(n_105),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_15),
.C(n_6),
.Y(n_105)
);

MAJx2_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_8),
.C(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_8),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_109),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_107),
.B(n_0),
.Y(n_110)
);

AOI211xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_108),
.B(n_3),
.C(n_4),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_112),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_3),
.Y(n_115)
);


endmodule