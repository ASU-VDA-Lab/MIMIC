module fake_jpeg_1703_n_389 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_389);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_389;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_73),
.Y(n_82)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_45),
.Y(n_131)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g108 ( 
.A(n_47),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_15),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_59),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_56),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_63),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_67),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_69),
.Y(n_104)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

AO22x1_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_74),
.B1(n_80),
.B2(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_78),
.Y(n_86)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_39),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_32),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_34),
.B1(n_32),
.B2(n_21),
.Y(n_84)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_84),
.A2(n_85),
.B(n_114),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_59),
.A2(n_34),
.B1(n_32),
.B2(n_21),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_34),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_50),
.B(n_35),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_94),
.Y(n_169)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_80),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_97),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_81),
.B(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_98),
.B(n_100),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_20),
.B(n_22),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_99),
.A2(n_108),
.B(n_104),
.C(n_83),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_17),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_45),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_110),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_102),
.B(n_103),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_20),
.B1(n_36),
.B2(n_23),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_105),
.A2(n_92),
.B1(n_133),
.B2(n_89),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_48),
.B(n_38),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_38),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_113),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_36),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_23),
.B1(n_17),
.B2(n_16),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_43),
.B(n_16),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_43),
.B(n_0),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_49),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_9),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_49),
.A2(n_22),
.B1(n_29),
.B2(n_2),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_130),
.B1(n_3),
.B2(n_4),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_49),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_136),
.B(n_138),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_137),
.A2(n_141),
.B1(n_153),
.B2(n_159),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_13),
.C(n_12),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_103),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_144),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_5),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_147),
.B(n_154),
.Y(n_204)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_152),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_6),
.Y(n_154)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_6),
.Y(n_155)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_155),
.B(n_175),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_156),
.Y(n_216)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_120),
.Y(n_157)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_9),
.B1(n_11),
.B2(n_6),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_93),
.A2(n_8),
.B1(n_82),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_162),
.A2(n_145),
.B1(n_154),
.B2(n_169),
.Y(n_214)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_119),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_87),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_170),
.Y(n_194)
);

O2A1O1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_112),
.B(n_124),
.C(n_116),
.Y(n_209)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_172),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_108),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_86),
.B(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_173),
.B(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_174),
.B(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_125),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_104),
.A2(n_126),
.B1(n_122),
.B2(n_87),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_122),
.B(n_121),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_108),
.A2(n_104),
.B1(n_92),
.B2(n_127),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_128),
.B1(n_116),
.B2(n_131),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_112),
.B1(n_96),
.B2(n_109),
.Y(n_219)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_89),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_127),
.C(n_133),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_187),
.B(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_134),
.B(n_128),
.C(n_121),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_142),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_214),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_SL g230 ( 
.A(n_209),
.B(n_163),
.C(n_181),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_135),
.A2(n_131),
.B1(n_124),
.B2(n_109),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_175),
.B1(n_178),
.B2(n_156),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_96),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_215),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_155),
.B(n_96),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_112),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_217),
.B(n_221),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_165),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_182),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_219),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_151),
.B(n_169),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_135),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_148),
.B(n_146),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_164),
.B(n_179),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_152),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_224),
.B(n_234),
.Y(n_282)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_205),
.A2(n_166),
.B1(n_163),
.B2(n_168),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_245),
.B1(n_248),
.B2(n_253),
.Y(n_258)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_163),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_231),
.B(n_232),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_177),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_176),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_235),
.B(n_252),
.Y(n_261)
);

BUFx24_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

INVx13_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_194),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_188),
.Y(n_240)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_241),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_191),
.A2(n_144),
.B1(n_143),
.B2(n_150),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_250),
.B1(n_251),
.B2(n_256),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_209),
.A2(n_181),
.B(n_176),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_197),
.B(n_198),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_205),
.A2(n_181),
.B1(n_140),
.B2(n_157),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_212),
.A2(n_149),
.B(n_158),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_249),
.A2(n_193),
.B(n_192),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_210),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_208),
.B(n_213),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_195),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_187),
.B(n_185),
.C(n_220),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_189),
.B(n_193),
.C(n_190),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_226),
.A2(n_219),
.B(n_185),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_257),
.A2(n_263),
.B(n_272),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_224),
.B(n_207),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_260),
.B(n_279),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_195),
.B1(n_217),
.B2(n_191),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_228),
.B1(n_223),
.B2(n_252),
.Y(n_289)
);

XNOR2x2_ASAP7_75t_SL g296 ( 
.A(n_267),
.B(n_244),
.Y(n_296)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_184),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_270),
.Y(n_285)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_203),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_203),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_267),
.C(n_234),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_233),
.A2(n_200),
.B(n_218),
.Y(n_272)
);

AND2x6_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_206),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_236),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_278),
.A2(n_246),
.B(n_236),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_198),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_197),
.B(n_196),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_280),
.Y(n_298)
);

AO22x1_ASAP7_75t_SL g281 ( 
.A1(n_248),
.A2(n_196),
.B1(n_183),
.B2(n_216),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_247),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_286),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_235),
.B1(n_228),
.B2(n_231),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_294),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_303),
.C(n_307),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_289),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_290),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_258),
.A2(n_239),
.B1(n_223),
.B2(n_232),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_291),
.A2(n_293),
.B1(n_304),
.B2(n_259),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_292),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_278),
.A2(n_239),
.B1(n_240),
.B2(n_225),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_238),
.Y(n_294)
);

XOR2x1_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_227),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_299),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_276),
.A2(n_237),
.B1(n_243),
.B2(n_241),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_306),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_268),
.B(n_281),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_229),
.C(n_251),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_241),
.B1(n_216),
.B2(n_183),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_236),
.C(n_282),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_273),
.B(n_257),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_276),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_312),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_313),
.B(n_321),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_261),
.C(n_263),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_318),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_316),
.B(n_330),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_280),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_300),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_303),
.B(n_269),
.C(n_283),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_296),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_324),
.A2(n_302),
.B(n_293),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_294),
.B(n_265),
.Y(n_328)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_328),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_297),
.B(n_274),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_307),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_334),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_291),
.Y(n_334)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_320),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_335),
.A2(n_341),
.B1(n_345),
.B2(n_323),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_328),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_339),
.B(n_330),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_346),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_326),
.A2(n_319),
.B1(n_313),
.B2(n_317),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_343),
.A2(n_295),
.B(n_324),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_285),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_344),
.Y(n_359)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_311),
.B(n_296),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

NAND2x1p5_ASAP7_75t_L g349 ( 
.A(n_332),
.B(n_341),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_349),
.B(n_357),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_351),
.B(n_354),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_337),
.A2(n_317),
.B1(n_298),
.B2(n_312),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_352),
.A2(n_353),
.B(n_355),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_337),
.A2(n_315),
.B1(n_317),
.B2(n_298),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_342),
.A2(n_315),
.B1(n_323),
.B2(n_310),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_318),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_331),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_360),
.A2(n_310),
.B(n_347),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_356),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_359),
.B(n_340),
.C(n_331),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_363),
.B(n_364),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_333),
.C(n_346),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_365),
.B(n_350),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_325),
.C(n_336),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_366),
.B(n_367),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_358),
.B(n_325),
.C(n_336),
.Y(n_367)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_371),
.B(n_372),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_368),
.A2(n_356),
.B(n_349),
.Y(n_372)
);

NAND2x1_ASAP7_75t_SL g374 ( 
.A(n_369),
.B(n_299),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_374),
.B(n_375),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_353),
.B(n_343),
.Y(n_375)
);

AOI322xp5_ASAP7_75t_L g377 ( 
.A1(n_370),
.A2(n_369),
.A3(n_275),
.B1(n_270),
.B2(n_361),
.C1(n_327),
.C2(n_321),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_374),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_379),
.B(n_376),
.C(n_373),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_SL g384 ( 
.A(n_381),
.B(n_382),
.C(n_383),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_329),
.Y(n_383)
);

NOR3xp33_ASAP7_75t_SL g385 ( 
.A(n_382),
.B(n_380),
.C(n_318),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_385),
.A2(n_295),
.B(n_352),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_386),
.A2(n_384),
.B1(n_286),
.B2(n_306),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_304),
.B(n_301),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_388),
.B(n_281),
.Y(n_389)
);


endmodule