module fake_netlist_5_1012_n_1975 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1975);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1975;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_108),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_97),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_139),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_10),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_17),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_80),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_84),
.Y(n_214)
);

BUFx4f_ASAP7_75t_SL g215 ( 
.A(n_39),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_99),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_202),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_177),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_172),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_125),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_129),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_86),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_103),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_137),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_63),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_29),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_194),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_74),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_61),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_44),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_133),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_169),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_63),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_144),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_55),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_163),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_126),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_39),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_29),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_65),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_110),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_7),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_79),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_130),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_167),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_58),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_191),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_178),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_145),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_118),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_138),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_112),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_190),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_155),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_111),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_136),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_64),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_3),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_87),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_131),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_160),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_181),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_17),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_42),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_16),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_81),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_113),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_52),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_93),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_117),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_127),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_43),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_106),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_68),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_16),
.Y(n_289)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_171),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_30),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_193),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_71),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_28),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_3),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_56),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_59),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_4),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_122),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_170),
.Y(n_301)
);

BUFx10_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_151),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_77),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_92),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_15),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_105),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_96),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_20),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_124),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_73),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_195),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_134),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_24),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_11),
.Y(n_317)
);

BUFx5_ASAP7_75t_L g318 ( 
.A(n_32),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_76),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_95),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_186),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_128),
.Y(n_322)
);

BUFx8_ASAP7_75t_SL g323 ( 
.A(n_147),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_123),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_24),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_156),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_164),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_197),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_22),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_101),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_201),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_31),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_46),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_158),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_25),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_5),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_12),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_0),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_62),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_33),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_104),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_120),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_18),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_98),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_88),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_27),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_62),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_59),
.Y(n_349)
);

BUFx5_ASAP7_75t_L g350 ( 
.A(n_149),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_13),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_162),
.Y(n_352)
);

INVx4_ASAP7_75t_R g353 ( 
.A(n_56),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_146),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_19),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g356 ( 
.A(n_12),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_19),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_153),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_85),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_140),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_11),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_148),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_35),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_27),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_75),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_142),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g367 ( 
.A(n_28),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_26),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_30),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_42),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_173),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_44),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_33),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_22),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_54),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_9),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_188),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_82),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_15),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_143),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_51),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_165),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_166),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_55),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_184),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_8),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_200),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_20),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_141),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_83),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_38),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_180),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_176),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_107),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_40),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_67),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_91),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_53),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_192),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_60),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_13),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_183),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_45),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_89),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_318),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_318),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_318),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_318),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_318),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_318),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_401),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_205),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_308),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_205),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_367),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_311),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_223),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_209),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_228),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_237),
.Y(n_425)
);

INVxp33_ASAP7_75t_SL g426 ( 
.A(n_401),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_245),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_239),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_238),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_325),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_352),
.B(n_1),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_223),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_244),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_225),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_232),
.B(n_2),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_400),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_225),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_248),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_236),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_311),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_379),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_302),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_214),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_252),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_377),
.Y(n_449)
);

NOR2xp67_ASAP7_75t_L g450 ( 
.A(n_232),
.B(n_2),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_379),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_253),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_207),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_222),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_254),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_227),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_213),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_236),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_403),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_233),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_274),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_389),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_234),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_241),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_260),
.Y(n_466)
);

NOR2xp67_ASAP7_75t_L g467 ( 
.A(n_338),
.B(n_7),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_276),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_280),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_286),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_240),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_269),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_277),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_352),
.B(n_8),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_240),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_289),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_297),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_271),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_298),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_213),
.B(n_199),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_291),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_268),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_295),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_216),
.B(n_10),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_303),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_284),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_284),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_304),
.B(n_14),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_271),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_302),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_340),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_340),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_307),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_296),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_214),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_317),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_326),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_330),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_363),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_333),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_334),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_337),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_268),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_373),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_285),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_381),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_285),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_482),
.B(n_235),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_430),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_413),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_434),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_427),
.A2(n_275),
.B1(n_243),
.B2(n_335),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_458),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_503),
.B(n_338),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_409),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_423),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_431),
.A2(n_273),
.B(n_216),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_415),
.B(n_224),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_410),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_449),
.B(n_217),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_437),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_415),
.B(n_218),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_437),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_412),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_405),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_419),
.B(n_243),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_R g533 ( 
.A(n_423),
.B(n_219),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_480),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_424),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_458),
.B(n_283),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_424),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_416),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_484),
.A2(n_281),
.B(n_273),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_421),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_432),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_405),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_443),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_406),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_480),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g548 ( 
.A(n_419),
.B(n_411),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_425),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_425),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_480),
.B(n_283),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_435),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_428),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_439),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_420),
.B(n_442),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_428),
.B(n_433),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_441),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_426),
.B(n_251),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_407),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_459),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_433),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_480),
.B(n_394),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_440),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_440),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_471),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_407),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_447),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_475),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_504),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_R g573 ( 
.A(n_447),
.B(n_452),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_452),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_445),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_495),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_414),
.B(n_394),
.Y(n_577)
);

CKINVDCx11_ASAP7_75t_R g578 ( 
.A(n_478),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_495),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_504),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_456),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_R g583 ( 
.A(n_456),
.B(n_468),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_506),
.Y(n_584)
);

XNOR2x2_ASAP7_75t_R g585 ( 
.A(n_489),
.B(n_14),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_474),
.B(n_282),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_417),
.B(n_224),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_486),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_586),
.B(n_468),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_517),
.B(n_436),
.Y(n_591)
);

INVx2_ASAP7_75t_SL g592 ( 
.A(n_536),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_561),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_561),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_462),
.Y(n_595)
);

BUFx6f_ASAP7_75t_L g596 ( 
.A(n_534),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_555),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_536),
.B(n_470),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_534),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_534),
.A2(n_438),
.B1(n_488),
.B2(n_467),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_526),
.B(n_560),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_513),
.Y(n_603)
);

BUFx10_ASAP7_75t_L g604 ( 
.A(n_548),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_534),
.B(n_418),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_534),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_534),
.A2(n_438),
.B1(n_450),
.B2(n_454),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_510),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_469),
.Y(n_612)
);

BUFx2_ASAP7_75t_L g613 ( 
.A(n_573),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_519),
.B(n_493),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_510),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_530),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_547),
.B(n_469),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_579),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_517),
.B(n_476),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_547),
.B(n_476),
.Y(n_620)
);

AND2x6_ASAP7_75t_L g621 ( 
.A(n_547),
.B(n_281),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_551),
.B(n_288),
.Y(n_622)
);

AND2x6_ASAP7_75t_L g623 ( 
.A(n_564),
.B(n_288),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_517),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_531),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_519),
.B(n_477),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_579),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_513),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_579),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_531),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_531),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_516),
.B(n_454),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_531),
.B(n_477),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_545),
.B(n_479),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_577),
.B(n_429),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_535),
.B(n_479),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_513),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_539),
.A2(n_388),
.B1(n_301),
.B2(n_359),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_545),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_528),
.B(n_485),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_575),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_545),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_513),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_583),
.Y(n_644)
);

BUFx10_ASAP7_75t_L g645 ( 
.A(n_537),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_524),
.B(n_485),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_518),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_569),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_545),
.Y(n_649)
);

INVx5_ASAP7_75t_L g650 ( 
.A(n_518),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

BUFx10_ASAP7_75t_L g652 ( 
.A(n_549),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_588),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_525),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_463),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_518),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_518),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_533),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_569),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_532),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_525),
.B(n_496),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_542),
.B(n_496),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_542),
.B(n_500),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_518),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_542),
.B(n_500),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_522),
.B(n_490),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_569),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_550),
.B(n_501),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g669 ( 
.A(n_518),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_521),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_521),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_523),
.B(n_453),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_521),
.Y(n_673)
);

AOI22xp33_ASAP7_75t_L g674 ( 
.A1(n_539),
.A2(n_301),
.B1(n_359),
.B2(n_460),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_521),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_553),
.B(n_501),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_575),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_521),
.B(n_293),
.Y(n_678)
);

BUFx4f_ASAP7_75t_L g679 ( 
.A(n_521),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_556),
.B(n_502),
.Y(n_680)
);

BUFx8_ASAP7_75t_SL g681 ( 
.A(n_538),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_539),
.A2(n_556),
.B1(n_568),
.B2(n_523),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_515),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_557),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_578),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_563),
.B(n_502),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_556),
.B(n_390),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_565),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_568),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_566),
.B(n_293),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_570),
.Y(n_691)
);

OAI22xp33_ASAP7_75t_L g692 ( 
.A1(n_574),
.A2(n_294),
.B1(n_369),
.B2(n_336),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_539),
.Y(n_694)
);

BUFx6f_ASAP7_75t_SL g695 ( 
.A(n_572),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_580),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_580),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_569),
.B(n_399),
.Y(n_698)
);

AND2x2_ASAP7_75t_SL g699 ( 
.A(n_582),
.B(n_293),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_582),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_581),
.B(n_293),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_584),
.B(n_208),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_584),
.B(n_455),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_508),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_508),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_515),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_576),
.B(n_226),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_543),
.B(n_457),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_511),
.Y(n_709)
);

BUFx10_ASAP7_75t_L g710 ( 
.A(n_543),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_511),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_540),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_576),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_512),
.B(n_214),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_544),
.B(n_309),
.Y(n_715)
);

BUFx4f_ASAP7_75t_L g716 ( 
.A(n_512),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_514),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_514),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_520),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_544),
.B(n_461),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_576),
.B(n_247),
.Y(n_721)
);

INVxp33_ASAP7_75t_L g722 ( 
.A(n_587),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_587),
.B(n_444),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_520),
.B(n_464),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_576),
.B(n_203),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_546),
.B(n_465),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_527),
.B(n_204),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_527),
.B(n_466),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_529),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_529),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_546),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_558),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_558),
.B(n_206),
.Y(n_733)
);

AO22x2_ASAP7_75t_L g734 ( 
.A1(n_585),
.A2(n_354),
.B1(n_346),
.B2(n_345),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_589),
.Y(n_735)
);

AND2x2_ASAP7_75t_SL g736 ( 
.A(n_589),
.B(n_249),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_541),
.B(n_210),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_SL g738 ( 
.A(n_552),
.B(n_275),
.C(n_505),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_571),
.B(n_472),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_567),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_559),
.A2(n_473),
.B1(n_499),
.B2(n_498),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_736),
.A2(n_263),
.B1(n_358),
.B2(n_362),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_602),
.B(n_309),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_590),
.B(n_640),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_606),
.B(n_255),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_590),
.B(n_324),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_653),
.B(n_612),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_653),
.B(n_324),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_614),
.B(n_666),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_507),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_612),
.B(n_335),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_713),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_736),
.B(n_266),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_715),
.B(n_279),
.C(n_272),
.Y(n_755)
);

NAND2x1_ASAP7_75t_L g756 ( 
.A(n_596),
.B(n_287),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_646),
.A2(n_392),
.B1(n_319),
.B2(n_331),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_596),
.B(n_305),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_596),
.B(n_312),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_658),
.B(n_302),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_626),
.B(n_392),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_713),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_739),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_640),
.B(n_662),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_596),
.B(n_320),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_648),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_648),
.Y(n_767)
);

BUFx8_ASAP7_75t_L g768 ( 
.A(n_691),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_663),
.B(n_215),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_600),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_665),
.B(n_219),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_680),
.B(n_220),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_600),
.B(n_321),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_607),
.B(n_601),
.C(n_619),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_723),
.B(n_316),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_600),
.B(n_322),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_600),
.B(n_329),
.Y(n_777)
);

INVx4_ASAP7_75t_L g778 ( 
.A(n_624),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_592),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_632),
.B(n_595),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_696),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_619),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_696),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_696),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_621),
.B(n_674),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_593),
.B(n_332),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_594),
.B(n_342),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_648),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_592),
.B(n_365),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_655),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_661),
.B(n_220),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_633),
.B(n_221),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_699),
.B(n_371),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_697),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_724),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_624),
.B(n_481),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_634),
.B(n_221),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_700),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_638),
.A2(n_385),
.B1(n_387),
.B2(n_397),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_646),
.B(n_402),
.Y(n_800)
);

NAND2xp33_ASAP7_75t_L g801 ( 
.A(n_621),
.B(n_214),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_630),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_659),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_681),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_684),
.B(n_402),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_699),
.B(n_211),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_722),
.B(n_339),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_647),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_605),
.A2(n_261),
.B(n_300),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_659),
.Y(n_810)
);

BUFx8_ASAP7_75t_L g811 ( 
.A(n_613),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_719),
.B(n_212),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_617),
.B(n_229),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_719),
.B(n_230),
.Y(n_814)
);

O2A1O1Ixp5_ASAP7_75t_L g815 ( 
.A1(n_702),
.A2(n_483),
.B(n_497),
.C(n_494),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_731),
.Y(n_816)
);

NAND2x1p5_ASAP7_75t_L g817 ( 
.A(n_630),
.B(n_487),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_722),
.B(n_341),
.Y(n_818)
);

INVx8_ASAP7_75t_L g819 ( 
.A(n_591),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_735),
.B(n_231),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_687),
.B(n_242),
.Y(n_821)
);

BUFx6f_ASAP7_75t_L g822 ( 
.A(n_639),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_621),
.B(n_214),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_639),
.B(n_246),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_704),
.B(n_250),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_620),
.B(n_710),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_635),
.B(n_347),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_737),
.B(n_690),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_705),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_688),
.B(n_256),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_690),
.B(n_348),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_701),
.B(n_351),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_709),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_711),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_717),
.B(n_257),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_667),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_667),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_644),
.B(n_316),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_667),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_710),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_718),
.B(n_258),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_608),
.Y(n_844)
);

NOR3xp33_ASAP7_75t_L g845 ( 
.A(n_715),
.B(n_361),
.C(n_355),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_729),
.B(n_259),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_701),
.B(n_357),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_708),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_724),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_608),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_610),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_616),
.B(n_364),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_708),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_708),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_610),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_710),
.B(n_262),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_597),
.B(n_264),
.Y(n_857)
);

BUFx12f_ASAP7_75t_L g858 ( 
.A(n_712),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_625),
.B(n_265),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_720),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_742),
.B(n_368),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_599),
.B(n_727),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_615),
.Y(n_863)
);

NOR3xp33_ASAP7_75t_L g864 ( 
.A(n_738),
.B(n_391),
.C(n_370),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_631),
.B(n_267),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_732),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_642),
.B(n_278),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_591),
.A2(n_360),
.B1(n_292),
.B2(n_299),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_649),
.B(n_306),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_733),
.B(n_372),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_591),
.B(n_374),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_615),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_618),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_622),
.A2(n_214),
.B1(n_350),
.B2(n_290),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_728),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_591),
.B(n_375),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_622),
.A2(n_214),
.B1(n_270),
.B2(n_290),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_310),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_668),
.B(n_313),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_720),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_732),
.B(n_314),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_720),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_621),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_732),
.B(n_315),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_732),
.B(n_327),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_676),
.B(n_316),
.Y(n_886)
);

BUFx5_ASAP7_75t_L g887 ( 
.A(n_621),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_686),
.B(n_562),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_694),
.B(n_328),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_726),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_728),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_618),
.Y(n_892)
);

OR2x2_ASAP7_75t_L g893 ( 
.A(n_740),
.B(n_386),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_622),
.A2(n_350),
.B1(n_270),
.B2(n_290),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_694),
.B(n_343),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_726),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_627),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_726),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_627),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_695),
.A2(n_380),
.B1(n_382),
.B2(n_383),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_730),
.B(n_366),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_716),
.B(n_378),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_730),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_695),
.A2(n_404),
.B1(n_393),
.B2(n_396),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_725),
.B(n_350),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_621),
.Y(n_906)
);

AND2x2_ASAP7_75t_SL g907 ( 
.A(n_714),
.B(n_492),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_716),
.B(n_350),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_703),
.B(n_398),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_629),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_695),
.A2(n_270),
.B1(n_290),
.B2(n_350),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_716),
.B(n_350),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_660),
.A2(n_270),
.B1(n_290),
.B2(n_350),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_785),
.A2(n_682),
.B(n_669),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_907),
.A2(n_679),
.B(n_672),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_745),
.B(n_688),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_763),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_907),
.A2(n_679),
.B(n_672),
.Y(n_918)
);

CKINVDCx8_ASAP7_75t_R g919 ( 
.A(n_804),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_889),
.A2(n_679),
.B(n_672),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_862),
.A2(n_672),
.B(n_689),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_764),
.B(n_862),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_895),
.A2(n_609),
.B(n_611),
.Y(n_923)
);

OAI21xp33_ASAP7_75t_L g924 ( 
.A1(n_747),
.A2(n_692),
.B(n_703),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_793),
.A2(n_678),
.B(n_702),
.C(n_721),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_781),
.B(n_703),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_764),
.B(n_703),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_795),
.B(n_693),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_908),
.A2(n_609),
.B(n_611),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_795),
.B(n_603),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_912),
.A2(n_609),
.B(n_611),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_905),
.A2(n_714),
.B(n_656),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_748),
.A2(n_678),
.B(n_721),
.C(n_707),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_849),
.B(n_603),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_746),
.A2(n_656),
.B(n_671),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_783),
.B(n_636),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_808),
.A2(n_656),
.B(n_637),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_802),
.Y(n_938)
);

BUFx3_ASAP7_75t_L g939 ( 
.A(n_858),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_761),
.B(n_741),
.C(n_712),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_645),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_754),
.A2(n_670),
.B(n_673),
.Y(n_942)
);

BUFx6f_ASAP7_75t_L g943 ( 
.A(n_802),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_774),
.A2(n_603),
.B1(n_657),
.B2(n_675),
.Y(n_944)
);

NAND3xp33_ASAP7_75t_L g945 ( 
.A(n_761),
.B(n_395),
.C(n_707),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_849),
.B(n_641),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_875),
.A2(n_651),
.B(n_654),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_875),
.B(n_641),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_886),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_802),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_891),
.A2(n_629),
.B(n_677),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_752),
.B(n_685),
.C(n_604),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_784),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_SL g954 ( 
.A(n_768),
.B(n_645),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_808),
.A2(n_637),
.B(n_628),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_830),
.A2(n_677),
.B(n_706),
.C(n_683),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_816),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_790),
.Y(n_958)
);

OAI21xp33_ASAP7_75t_L g959 ( 
.A1(n_807),
.A2(n_734),
.B(n_491),
.Y(n_959)
);

INVx1_ASAP7_75t_SL g960 ( 
.A(n_751),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_743),
.A2(n_782),
.B1(n_830),
.B2(n_891),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_881),
.A2(n_637),
.B(n_628),
.Y(n_962)
);

HB1xp67_ASAP7_75t_L g963 ( 
.A(n_790),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_782),
.B(n_622),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_884),
.A2(n_637),
.B(n_628),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_744),
.B(n_604),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_825),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_799),
.A2(n_683),
.B(n_706),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_885),
.A2(n_628),
.B(n_657),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_743),
.A2(n_734),
.B1(n_647),
.B2(n_664),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_806),
.A2(n_623),
.B(n_622),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_802),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_792),
.B(n_622),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_760),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_770),
.A2(n_664),
.B(n_647),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_770),
.A2(n_664),
.B(n_647),
.Y(n_976)
);

AO32x2_ASAP7_75t_L g977 ( 
.A1(n_778),
.A2(n_623),
.A3(n_734),
.B1(n_604),
.B2(n_353),
.Y(n_977)
);

NOR2x1p5_ASAP7_75t_SL g978 ( 
.A(n_887),
.B(n_270),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_779),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_792),
.B(n_623),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_797),
.B(n_623),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_800),
.A2(n_779),
.B(n_789),
.C(n_828),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_842),
.B(n_652),
.Y(n_983)
);

AOI21x1_ASAP7_75t_L g984 ( 
.A1(n_758),
.A2(n_487),
.B(n_491),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_794),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_770),
.A2(n_664),
.B(n_643),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_870),
.B(n_652),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_807),
.B(n_652),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_797),
.B(n_623),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_771),
.B(n_772),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_757),
.B(n_685),
.C(n_492),
.Y(n_991)
);

OAI21xp33_ASAP7_75t_L g992 ( 
.A1(n_818),
.A2(n_344),
.B(n_356),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_770),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_848),
.A2(n_854),
.B1(n_860),
.B2(n_898),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_826),
.A2(n_643),
.B(n_650),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_859),
.A2(n_643),
.B(n_650),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_749),
.B(n_323),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_844),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_818),
.B(n_344),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_829),
.B(n_344),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_865),
.A2(n_643),
.B(n_650),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_771),
.B(n_623),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_833),
.A2(n_643),
.B(n_650),
.C(n_270),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_833),
.A2(n_650),
.B(n_270),
.C(n_290),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_822),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_772),
.B(n_290),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_822),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_801),
.A2(n_224),
.B(n_132),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_L g1009 ( 
.A(n_888),
.B(n_323),
.C(n_376),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_768),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_811),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_791),
.B(n_21),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_811),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_867),
.A2(n_66),
.B(n_198),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_869),
.A2(n_121),
.B(n_72),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_791),
.B(n_21),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_805),
.A2(n_384),
.B(n_376),
.C(n_356),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_822),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_861),
.A2(n_384),
.B(n_376),
.Y(n_1019)
);

OA21x2_ASAP7_75t_L g1020 ( 
.A1(n_759),
.A2(n_196),
.B(n_187),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_798),
.Y(n_1021)
);

AO22x1_ASAP7_75t_L g1022 ( 
.A1(n_755),
.A2(n_384),
.B1(n_356),
.B2(n_26),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_831),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_829),
.B(n_23),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_780),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_870),
.A2(n_182),
.B(n_179),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_850),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_835),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_836),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_821),
.B(n_23),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_851),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_878),
.B(n_853),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_824),
.A2(n_175),
.B(n_168),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_887),
.B(n_161),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_857),
.A2(n_25),
.B(n_31),
.C(n_32),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_866),
.A2(n_152),
.B(n_119),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_755),
.A2(n_786),
.B(n_787),
.C(n_847),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_796),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_866),
.A2(n_116),
.B(n_114),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_822),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_880),
.A2(n_109),
.B1(n_100),
.B2(n_94),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_796),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_834),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_882),
.B(n_34),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_890),
.B(n_36),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_896),
.B(n_37),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_812),
.A2(n_90),
.B(n_78),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_765),
.A2(n_70),
.B(n_38),
.Y(n_1048)
);

OAI22x1_ASAP7_75t_L g1049 ( 
.A1(n_840),
.A2(n_834),
.B1(n_847),
.B2(n_909),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_769),
.B(n_37),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_L g1051 ( 
.A(n_864),
.B(n_41),
.C(n_45),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_773),
.A2(n_777),
.B(n_776),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_852),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_769),
.B(n_41),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_901),
.A2(n_46),
.B(n_47),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_815),
.A2(n_48),
.B(n_49),
.C(n_50),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_814),
.B(n_48),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_815),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_753),
.A2(n_53),
.B(n_54),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_778),
.B(n_832),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_855),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_766),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_902),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_863),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_893),
.Y(n_1065)
);

O2A1O1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_813),
.A2(n_57),
.B(n_845),
.C(n_879),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_762),
.A2(n_841),
.B(n_767),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_788),
.A2(n_839),
.B(n_803),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_810),
.A2(n_838),
.B(n_823),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_900),
.Y(n_1070)
);

AO21x1_ASAP7_75t_L g1071 ( 
.A1(n_845),
.A2(n_913),
.B(n_817),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_817),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_820),
.A2(n_843),
.B(n_846),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_827),
.B(n_837),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_871),
.B(n_876),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_909),
.B(n_876),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_872),
.B(n_897),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_873),
.B(n_910),
.Y(n_1078)
);

NOR2xp67_ASAP7_75t_L g1079 ( 
.A(n_904),
.B(n_868),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_892),
.A2(n_899),
.B(n_883),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_756),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_883),
.A2(n_906),
.B(n_809),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_883),
.A2(n_906),
.B(n_856),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_874),
.A2(n_894),
.B(n_877),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_871),
.B(n_819),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_874),
.A2(n_877),
.B(n_894),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_911),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_819),
.B(n_887),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_887),
.A2(n_883),
.B(n_906),
.Y(n_1089)
);

NOR2xp67_ASAP7_75t_SL g1090 ( 
.A(n_906),
.B(n_887),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_819),
.A2(n_887),
.B(n_864),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_745),
.A2(n_793),
.B(n_748),
.C(n_754),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_745),
.B(n_764),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_750),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_903),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_785),
.A2(n_606),
.B(n_600),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_745),
.A2(n_764),
.B(n_862),
.C(n_590),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_745),
.A2(n_795),
.B(n_875),
.C(n_849),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_802),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_785),
.A2(n_606),
.B(n_600),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_785),
.A2(n_606),
.B(n_600),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_785),
.A2(n_606),
.B(n_600),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_745),
.B(n_764),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_785),
.A2(n_600),
.B(n_596),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_914),
.A2(n_932),
.B(n_1052),
.Y(n_1105)
);

OAI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1097),
.A2(n_1103),
.B(n_1093),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_922),
.A2(n_1086),
.B1(n_990),
.B2(n_961),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1096),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_916),
.A2(n_1076),
.B1(n_927),
.B2(n_1012),
.Y(n_1109)
);

O2A1O1Ixp5_ASAP7_75t_L g1110 ( 
.A1(n_1016),
.A2(n_1006),
.B(n_920),
.C(n_980),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1098),
.B(n_928),
.Y(n_1111)
);

NAND3xp33_ASAP7_75t_SL g1112 ( 
.A(n_960),
.B(n_966),
.C(n_997),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1024),
.A2(n_1079),
.B1(n_921),
.B2(n_1050),
.Y(n_1113)
);

OAI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1082),
.A2(n_1100),
.B(n_1096),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_926),
.B(n_936),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1101),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1101),
.A2(n_1102),
.B(n_1089),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1094),
.B(n_941),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_962),
.A2(n_965),
.B(n_1068),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1000),
.B(n_999),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_946),
.B(n_948),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_932),
.A2(n_1052),
.B(n_920),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_985),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1068),
.A2(n_1069),
.B(n_923),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1069),
.A2(n_923),
.B(n_969),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1074),
.B(n_988),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_917),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_943),
.Y(n_1128)
);

NAND3x1_ASAP7_75t_L g1129 ( 
.A(n_952),
.B(n_1009),
.C(n_1051),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1065),
.B(n_974),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_929),
.A2(n_931),
.B(n_1067),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1092),
.A2(n_924),
.B(n_1037),
.C(n_982),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1032),
.B(n_1021),
.Y(n_1133)
);

AOI21x1_ASAP7_75t_L g1134 ( 
.A1(n_915),
.A2(n_918),
.B(n_973),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1080),
.A2(n_935),
.B(n_976),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1023),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1028),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1025),
.B(n_1075),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1066),
.A2(n_1084),
.B(n_1073),
.C(n_1026),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1029),
.B(n_1049),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_930),
.B(n_934),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1073),
.A2(n_915),
.B(n_918),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_958),
.Y(n_1143)
);

O2A1O1Ixp5_ASAP7_75t_L g1144 ( 
.A1(n_981),
.A2(n_989),
.B(n_1002),
.C(n_971),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_956),
.A2(n_925),
.B(n_964),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1054),
.B(n_1030),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_919),
.Y(n_1147)
);

OAI21x1_ASAP7_75t_SL g1148 ( 
.A1(n_1091),
.A2(n_1083),
.B(n_1088),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_943),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_944),
.A2(n_942),
.B(n_933),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_1003),
.A2(n_968),
.B(n_1004),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1005),
.B(n_1007),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_957),
.Y(n_1153)
);

NAND2x1_ASAP7_75t_L g1154 ( 
.A(n_1090),
.B(n_1005),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1087),
.A2(n_1080),
.B(n_951),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_935),
.A2(n_975),
.B(n_995),
.Y(n_1156)
);

AOI21xp33_ASAP7_75t_L g1157 ( 
.A1(n_945),
.A2(n_1057),
.B(n_1063),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_949),
.B(n_967),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_959),
.A2(n_992),
.B(n_1019),
.C(n_1091),
.Y(n_1159)
);

AOI221xp5_ASAP7_75t_L g1160 ( 
.A1(n_1022),
.A2(n_1070),
.B1(n_940),
.B2(n_963),
.C(n_1043),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1034),
.A2(n_1083),
.B(n_937),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_955),
.A2(n_1001),
.B(n_996),
.Y(n_1162)
);

AOI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_987),
.A2(n_1085),
.B1(n_926),
.B2(n_1053),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_979),
.B(n_1038),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_936),
.B(n_1042),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_947),
.A2(n_1078),
.B(n_1077),
.Y(n_1166)
);

AOI21xp33_ASAP7_75t_L g1167 ( 
.A1(n_1035),
.A2(n_1046),
.B(n_1045),
.Y(n_1167)
);

BUFx6f_ASAP7_75t_L g1168 ( 
.A(n_943),
.Y(n_1168)
);

BUFx8_ASAP7_75t_L g1169 ( 
.A(n_1010),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_986),
.A2(n_994),
.B(n_1072),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1044),
.A2(n_1017),
.B(n_1058),
.C(n_1056),
.Y(n_1171)
);

OAI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_970),
.A2(n_1008),
.B(n_1095),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1008),
.A2(n_1062),
.B(n_1027),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_993),
.A2(n_1060),
.B(n_938),
.Y(n_1174)
);

AND2x4_ASAP7_75t_L g1175 ( 
.A(n_1007),
.B(n_1072),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_939),
.B(n_1011),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1041),
.A2(n_950),
.B1(n_1018),
.B2(n_972),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_950),
.A2(n_1018),
.B1(n_972),
.B2(n_991),
.Y(n_1178)
);

O2A1O1Ixp5_ASAP7_75t_L g1179 ( 
.A1(n_1071),
.A2(n_984),
.B(n_1048),
.C(n_1081),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1013),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_998),
.B(n_1031),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_938),
.A2(n_1099),
.B(n_1040),
.Y(n_1182)
);

O2A1O1Ixp5_ASAP7_75t_L g1183 ( 
.A1(n_1048),
.A2(n_1015),
.B(n_1014),
.C(n_1047),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1040),
.A2(n_1099),
.B(n_1033),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1061),
.B(n_1064),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_983),
.B(n_950),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_972),
.Y(n_1187)
);

OR2x6_ASAP7_75t_L g1188 ( 
.A(n_1018),
.B(n_1059),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_977),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_1036),
.A2(n_1039),
.B(n_1020),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1055),
.A2(n_1020),
.B(n_978),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_954),
.B(n_977),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_977),
.B(n_750),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_919),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1025),
.Y(n_1197)
);

NAND2x1_ASAP7_75t_L g1198 ( 
.A(n_1090),
.B(n_770),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1199)
);

OAI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_988),
.B(n_745),
.Y(n_1203)
);

OR2x6_ASAP7_75t_L g1204 ( 
.A(n_939),
.B(n_819),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_919),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_921),
.A2(n_942),
.B(n_920),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_953),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_926),
.B(n_936),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_919),
.Y(n_1209)
);

AOI221xp5_ASAP7_75t_L g1210 ( 
.A1(n_1093),
.A2(n_745),
.B1(n_747),
.B2(n_1103),
.C(n_692),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1093),
.B(n_1103),
.Y(n_1211)
);

AND2x6_ASAP7_75t_L g1212 ( 
.A(n_1088),
.B(n_883),
.Y(n_1212)
);

OAI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1097),
.A2(n_745),
.B(n_990),
.C(n_922),
.Y(n_1214)
);

OAI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_990),
.A2(n_745),
.B1(n_1103),
.B2(n_1093),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1025),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1093),
.B(n_745),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_926),
.B(n_936),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_988),
.B(n_745),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1097),
.A2(n_745),
.B(n_990),
.C(n_922),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1093),
.B(n_1103),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_943),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1093),
.A2(n_1103),
.B1(n_922),
.B2(n_1097),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1093),
.A2(n_1103),
.B1(n_922),
.B2(n_1097),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_SL g1232 ( 
.A(n_1097),
.B(n_1076),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1233)
);

BUFx3_ASAP7_75t_L g1234 ( 
.A(n_939),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_990),
.A2(n_745),
.B(n_1093),
.Y(n_1235)
);

INVxp67_ASAP7_75t_L g1236 ( 
.A(n_1025),
.Y(n_1236)
);

AOI221xp5_ASAP7_75t_L g1237 ( 
.A1(n_1093),
.A2(n_745),
.B1(n_747),
.B2(n_1103),
.C(n_692),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1093),
.B(n_1103),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_926),
.B(n_936),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1025),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_921),
.A2(n_942),
.B(n_920),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_985),
.Y(n_1244)
);

AOI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1076),
.A2(n_745),
.B1(n_1103),
.B2(n_1093),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1097),
.A2(n_914),
.B(n_1093),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_914),
.A2(n_600),
.B(n_596),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_921),
.A2(n_920),
.B(n_942),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_920),
.A2(n_918),
.B(n_915),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_921),
.A2(n_942),
.B(n_920),
.Y(n_1252)
);

AO21x1_ASAP7_75t_L g1253 ( 
.A1(n_990),
.A2(n_745),
.B(n_922),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1093),
.B(n_1103),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1104),
.A2(n_1082),
.B(n_1100),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1118),
.B(n_1120),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1218),
.A2(n_1210),
.B1(n_1237),
.B2(n_1232),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1105),
.A2(n_1161),
.B(n_1139),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1175),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1197),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1147),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1217),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1240),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1175),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1228),
.B(n_1149),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1122),
.A2(n_1150),
.B(n_1142),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1150),
.A2(n_1225),
.B(n_1214),
.Y(n_1267)
);

NAND2x1p5_ASAP7_75t_L g1268 ( 
.A(n_1228),
.B(n_1149),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_SL g1269 ( 
.A(n_1232),
.B(n_1205),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1245),
.B(n_1211),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1216),
.A2(n_1194),
.B1(n_1138),
.B2(n_1254),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1227),
.A2(n_1238),
.B1(n_1107),
.B2(n_1229),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1229),
.B(n_1231),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1117),
.A2(n_1195),
.B(n_1108),
.Y(n_1274)
);

OR2x6_ASAP7_75t_L g1275 ( 
.A(n_1204),
.B(n_1176),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1127),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1126),
.B(n_1130),
.Y(n_1277)
);

INVxp67_ASAP7_75t_L g1278 ( 
.A(n_1143),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1207),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1136),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1137),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1164),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_1236),
.Y(n_1283)
);

NOR2xp67_ASAP7_75t_L g1284 ( 
.A(n_1112),
.B(n_1209),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1199),
.A2(n_1223),
.B(n_1233),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1115),
.B(n_1208),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1199),
.A2(n_1223),
.B(n_1233),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1115),
.B(n_1208),
.Y(n_1288)
);

AND2x4_ASAP7_75t_L g1289 ( 
.A(n_1221),
.B(n_1239),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1107),
.A2(n_1231),
.B1(n_1106),
.B2(n_1235),
.Y(n_1290)
);

CKINVDCx8_ASAP7_75t_R g1291 ( 
.A(n_1180),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1200),
.A2(n_1213),
.B(n_1247),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1200),
.A2(n_1213),
.B(n_1247),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1106),
.A2(n_1235),
.B1(n_1248),
.B2(n_1215),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1169),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1169),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1203),
.B(n_1224),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1215),
.A2(n_1248),
.B(n_1201),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1221),
.B(n_1239),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1165),
.B(n_1133),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1121),
.B(n_1109),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1165),
.B(n_1204),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1196),
.A2(n_1222),
.B(n_1220),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1168),
.Y(n_1304)
);

HB1xp67_ASAP7_75t_L g1305 ( 
.A(n_1187),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1109),
.A2(n_1111),
.B1(n_1159),
.B2(n_1113),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1204),
.B(n_1244),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1202),
.A2(n_1219),
.B(n_1249),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1146),
.B(n_1141),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1234),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1253),
.B(n_1193),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1113),
.B(n_1132),
.Y(n_1312)
);

NAND2xp33_ASAP7_75t_L g1313 ( 
.A(n_1129),
.B(n_1212),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1160),
.B(n_1163),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1158),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1191),
.A2(n_1145),
.B(n_1148),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1140),
.B(n_1153),
.Y(n_1317)
);

INVx3_ASAP7_75t_SL g1318 ( 
.A(n_1176),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1181),
.B(n_1185),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1152),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1181),
.B(n_1185),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1176),
.Y(n_1322)
);

INVx3_ASAP7_75t_L g1323 ( 
.A(n_1152),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1168),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1128),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1128),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1166),
.B(n_1172),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1178),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1154),
.B(n_1198),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1186),
.B(n_1166),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1188),
.B(n_1157),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1155),
.A2(n_1250),
.B(n_1172),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1192),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1155),
.B(n_1167),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1188),
.Y(n_1335)
);

BUFx12f_ASAP7_75t_L g1336 ( 
.A(n_1188),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1178),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1157),
.A2(n_1167),
.B1(n_1189),
.B2(n_1250),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1189),
.B(n_1173),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1189),
.Y(n_1340)
);

NAND2x1p5_ASAP7_75t_L g1341 ( 
.A(n_1182),
.B(n_1170),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1177),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1173),
.B(n_1171),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1183),
.A2(n_1179),
.B(n_1110),
.C(n_1116),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1191),
.B(n_1145),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1177),
.B(n_1174),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1212),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_L g1348 ( 
.A(n_1251),
.B(n_1134),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1184),
.B(n_1114),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1206),
.A2(n_1252),
.B(n_1242),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1124),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1226),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1230),
.Y(n_1353)
);

AOI222xp33_ASAP7_75t_L g1354 ( 
.A1(n_1212),
.A2(n_1255),
.B1(n_1241),
.B2(n_1243),
.C1(n_1246),
.C2(n_1190),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1212),
.B(n_1252),
.Y(n_1355)
);

AOI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1206),
.A2(n_1242),
.B(n_1144),
.Y(n_1356)
);

BUFx12f_ASAP7_75t_L g1357 ( 
.A(n_1151),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1135),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1119),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1131),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1125),
.B(n_1156),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1162),
.A2(n_1105),
.B(n_1161),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1218),
.B(n_1093),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1194),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_SL g1365 ( 
.A(n_1234),
.Y(n_1365)
);

AOI222xp33_ASAP7_75t_L g1366 ( 
.A1(n_1210),
.A2(n_745),
.B1(n_1237),
.B2(n_1218),
.C1(n_747),
.C2(n_1103),
.Y(n_1366)
);

NOR2xp33_ASAP7_75t_L g1367 ( 
.A(n_1218),
.B(n_745),
.Y(n_1367)
);

OAI321xp33_ASAP7_75t_L g1368 ( 
.A1(n_1245),
.A2(n_745),
.A3(n_1103),
.B1(n_1093),
.B2(n_922),
.C(n_1097),
.Y(n_1368)
);

AOI211xp5_ASAP7_75t_L g1369 ( 
.A1(n_1218),
.A2(n_745),
.B(n_916),
.C(n_602),
.Y(n_1369)
);

A2O1A1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1218),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1218),
.B(n_1093),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1118),
.B(n_750),
.Y(n_1372)
);

INVx3_ASAP7_75t_SL g1373 ( 
.A(n_1147),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1118),
.B(n_750),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1123),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1218),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1376)
);

BUFx12f_ASAP7_75t_L g1377 ( 
.A(n_1169),
.Y(n_1377)
);

INVx5_ASAP7_75t_L g1378 ( 
.A(n_1149),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1218),
.B(n_745),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1149),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1218),
.B(n_745),
.Y(n_1381)
);

INVx1_ASAP7_75t_SL g1382 ( 
.A(n_1197),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1218),
.B(n_1093),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1149),
.Y(n_1384)
);

O2A1O1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1235),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1385)
);

O2A1O1Ixp33_ASAP7_75t_L g1386 ( 
.A1(n_1235),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1150),
.A2(n_1142),
.B(n_1122),
.Y(n_1387)
);

BUFx3_ASAP7_75t_L g1388 ( 
.A(n_1197),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1123),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1115),
.B(n_1208),
.Y(n_1390)
);

O2A1O1Ixp33_ASAP7_75t_L g1391 ( 
.A1(n_1235),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1126),
.B(n_780),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1218),
.A2(n_745),
.B1(n_1076),
.B2(n_990),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1197),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1218),
.A2(n_745),
.B1(n_1076),
.B2(n_990),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1126),
.B(n_780),
.Y(n_1396)
);

AO21x1_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_1107),
.B(n_1109),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1147),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1175),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1218),
.A2(n_745),
.B(n_1097),
.C(n_1093),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1118),
.B(n_750),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1340),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1367),
.A2(n_1379),
.B1(n_1381),
.B2(n_1269),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1282),
.Y(n_1404)
);

CKINVDCx10_ASAP7_75t_R g1405 ( 
.A(n_1365),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1256),
.B(n_1372),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1281),
.Y(n_1407)
);

INVx6_ASAP7_75t_L g1408 ( 
.A(n_1304),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1374),
.B(n_1401),
.Y(n_1409)
);

INVx5_ASAP7_75t_L g1410 ( 
.A(n_1304),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1393),
.B(n_1395),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1346),
.A2(n_1334),
.B(n_1306),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1304),
.Y(n_1413)
);

HB1xp67_ASAP7_75t_L g1414 ( 
.A(n_1337),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1269),
.A2(n_1314),
.B1(n_1271),
.B2(n_1290),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1335),
.B(n_1259),
.Y(n_1416)
);

AO21x1_ASAP7_75t_L g1417 ( 
.A1(n_1369),
.A2(n_1386),
.B(n_1385),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1363),
.B(n_1371),
.Y(n_1418)
);

NAND2x1_ASAP7_75t_L g1419 ( 
.A(n_1320),
.B(n_1323),
.Y(n_1419)
);

AO21x1_ASAP7_75t_SL g1420 ( 
.A1(n_1257),
.A2(n_1312),
.B(n_1311),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1363),
.B(n_1371),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1344),
.A2(n_1266),
.B(n_1258),
.Y(n_1422)
);

INVx6_ASAP7_75t_L g1423 ( 
.A(n_1378),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1378),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1369),
.A2(n_1383),
.B1(n_1370),
.B2(n_1400),
.Y(n_1425)
);

NAND2x1p5_ASAP7_75t_L g1426 ( 
.A(n_1378),
.B(n_1320),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1383),
.B(n_1270),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_1282),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1277),
.B(n_1300),
.Y(n_1429)
);

BUFx2_ASAP7_75t_SL g1430 ( 
.A(n_1365),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1366),
.A2(n_1376),
.B(n_1368),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1366),
.A2(n_1397),
.B1(n_1290),
.B2(n_1294),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1328),
.Y(n_1433)
);

AOI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1306),
.A2(n_1298),
.B(n_1356),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1294),
.A2(n_1273),
.B1(n_1272),
.B2(n_1270),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1296),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1375),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1388),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1389),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1291),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1362),
.A2(n_1303),
.B(n_1308),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1392),
.B(n_1396),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1336),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1394),
.Y(n_1444)
);

AO21x1_ASAP7_75t_L g1445 ( 
.A1(n_1391),
.A2(n_1272),
.B(n_1301),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1342),
.Y(n_1446)
);

BUFx12f_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

AOI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1285),
.A2(n_1292),
.B(n_1293),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1279),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1273),
.A2(n_1343),
.B1(n_1287),
.B2(n_1312),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1267),
.A2(n_1309),
.B1(n_1342),
.B2(n_1327),
.Y(n_1451)
);

AO21x1_ASAP7_75t_L g1452 ( 
.A1(n_1309),
.A2(n_1330),
.B(n_1327),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1341),
.A2(n_1350),
.B(n_1351),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1319),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1317),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1315),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1286),
.Y(n_1457)
);

CKINVDCx11_ASAP7_75t_R g1458 ( 
.A(n_1295),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1380),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1332),
.A2(n_1338),
.B(n_1348),
.Y(n_1460)
);

CKINVDCx6p67_ASAP7_75t_R g1461 ( 
.A(n_1373),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1360),
.A2(n_1353),
.B(n_1352),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1321),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1326),
.Y(n_1464)
);

AO21x2_ASAP7_75t_L g1465 ( 
.A1(n_1358),
.A2(n_1387),
.B(n_1355),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1297),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1311),
.Y(n_1467)
);

BUFx10_ASAP7_75t_L g1468 ( 
.A(n_1261),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1307),
.Y(n_1469)
);

BUFx8_ASAP7_75t_SL g1470 ( 
.A(n_1364),
.Y(n_1470)
);

INVx8_ASAP7_75t_L g1471 ( 
.A(n_1380),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1399),
.B(n_1264),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1345),
.A2(n_1331),
.B1(n_1313),
.B2(n_1284),
.Y(n_1473)
);

NAND2x1p5_ASAP7_75t_L g1474 ( 
.A(n_1399),
.B(n_1347),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1286),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1384),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1361),
.A2(n_1359),
.B(n_1349),
.Y(n_1477)
);

INVx8_ASAP7_75t_L g1478 ( 
.A(n_1384),
.Y(n_1478)
);

BUFx8_ASAP7_75t_SL g1479 ( 
.A(n_1398),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1302),
.B(n_1260),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1288),
.B(n_1390),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1324),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1339),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1384),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1316),
.Y(n_1485)
);

OAI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1368),
.A2(n_1275),
.B1(n_1322),
.B2(n_1318),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1263),
.Y(n_1487)
);

INVx4_ASAP7_75t_L g1488 ( 
.A(n_1275),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1357),
.A2(n_1333),
.B1(n_1316),
.B2(n_1275),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1263),
.A2(n_1382),
.B1(n_1283),
.B2(n_1262),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1302),
.A2(n_1382),
.B1(n_1390),
.B2(n_1299),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1349),
.Y(n_1492)
);

INVx6_ASAP7_75t_L g1493 ( 
.A(n_1288),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1289),
.B(n_1299),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1278),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1289),
.A2(n_1276),
.B1(n_1305),
.B2(n_1361),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1325),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_L g1498 ( 
.A1(n_1329),
.A2(n_1310),
.B1(n_1268),
.B2(n_1265),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1354),
.A2(n_1366),
.B1(n_1379),
.B2(n_1367),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1354),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1274),
.A2(n_1114),
.B(n_1108),
.Y(n_1501)
);

AND2x4_ASAP7_75t_L g1502 ( 
.A(n_1335),
.B(n_1259),
.Y(n_1502)
);

AOI222xp33_ASAP7_75t_L g1503 ( 
.A1(n_1367),
.A2(n_1381),
.B1(n_1379),
.B2(n_745),
.C1(n_747),
.C2(n_752),
.Y(n_1503)
);

OAI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1367),
.A2(n_1093),
.B1(n_1103),
.B2(n_922),
.Y(n_1504)
);

CKINVDCx8_ASAP7_75t_R g1505 ( 
.A(n_1261),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1336),
.Y(n_1506)
);

BUFx6f_ASAP7_75t_L g1507 ( 
.A(n_1304),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1392),
.B(n_1396),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1344),
.A2(n_1110),
.B(n_1122),
.Y(n_1509)
);

BUFx2_ASAP7_75t_SL g1510 ( 
.A(n_1365),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1304),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1257),
.A2(n_745),
.B(n_1097),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1280),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1393),
.A2(n_745),
.B1(n_1103),
.B2(n_1093),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1367),
.A2(n_745),
.B1(n_916),
.B2(n_1379),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1280),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1256),
.B(n_1372),
.Y(n_1517)
);

NAND2x1p5_ASAP7_75t_L g1518 ( 
.A(n_1304),
.B(n_1378),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_SL g1519 ( 
.A1(n_1367),
.A2(n_745),
.B1(n_1076),
.B2(n_1379),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1393),
.A2(n_745),
.B1(n_1103),
.B2(n_1093),
.Y(n_1520)
);

BUFx6f_ASAP7_75t_L g1521 ( 
.A(n_1304),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1366),
.A2(n_1379),
.B1(n_1381),
.B2(n_1367),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1367),
.B(n_1218),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1280),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1304),
.Y(n_1525)
);

BUFx12f_ASAP7_75t_L g1526 ( 
.A(n_1296),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1388),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1280),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1462),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1462),
.Y(n_1530)
);

OA21x2_ASAP7_75t_L g1531 ( 
.A1(n_1448),
.A2(n_1431),
.B(n_1432),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1433),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1442),
.B(n_1427),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1433),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1402),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1477),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1483),
.B(n_1467),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1480),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1485),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1479),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1522),
.B(n_1508),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1450),
.B(n_1429),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1522),
.B(n_1418),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1402),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1480),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1492),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1443),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1492),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1454),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1452),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1460),
.B(n_1454),
.Y(n_1552)
);

OR2x6_ASAP7_75t_L g1553 ( 
.A(n_1488),
.B(n_1412),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1446),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1446),
.Y(n_1555)
);

OR2x6_ASAP7_75t_L g1556 ( 
.A(n_1488),
.B(n_1445),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1465),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1434),
.A2(n_1417),
.B(n_1441),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1414),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1414),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1435),
.B(n_1432),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1404),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1435),
.B(n_1420),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1453),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1456),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1501),
.A2(n_1451),
.B(n_1512),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1509),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1463),
.B(n_1451),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1425),
.A2(n_1499),
.B(n_1489),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1509),
.A2(n_1422),
.B(n_1500),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1509),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1466),
.Y(n_1572)
);

HB1xp67_ASAP7_75t_L g1573 ( 
.A(n_1455),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1428),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1524),
.B(n_1500),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1437),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1524),
.B(n_1460),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1439),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1479),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1416),
.B(n_1502),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1422),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1487),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1407),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1528),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1513),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1516),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1443),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1415),
.B(n_1406),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1464),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1416),
.B(n_1502),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1489),
.B(n_1473),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1517),
.B(n_1409),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1499),
.A2(n_1473),
.B(n_1411),
.Y(n_1593)
);

INVx5_ASAP7_75t_L g1594 ( 
.A(n_1410),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1449),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1490),
.B(n_1496),
.Y(n_1596)
);

OR2x6_ASAP7_75t_L g1597 ( 
.A(n_1443),
.B(n_1430),
.Y(n_1597)
);

HB1xp67_ASAP7_75t_L g1598 ( 
.A(n_1482),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1421),
.B(n_1469),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1486),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1496),
.A2(n_1419),
.B(n_1474),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1444),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1519),
.B(n_1515),
.Y(n_1603)
);

BUFx3_ASAP7_75t_L g1604 ( 
.A(n_1506),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1486),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1490),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_1470),
.Y(n_1607)
);

OR2x6_ASAP7_75t_L g1608 ( 
.A(n_1510),
.B(n_1472),
.Y(n_1608)
);

AO21x2_ASAP7_75t_L g1609 ( 
.A1(n_1504),
.A2(n_1520),
.B(n_1514),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1426),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1523),
.B(n_1403),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1426),
.A2(n_1518),
.B(n_1498),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1491),
.B(n_1481),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1552),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.B(n_1497),
.Y(n_1615)
);

NOR3xp33_ASAP7_75t_L g1616 ( 
.A(n_1603),
.B(n_1403),
.C(n_1504),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1552),
.B(n_1506),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1570),
.B(n_1506),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1476),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1567),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1553),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1566),
.B(n_1484),
.Y(n_1622)
);

BUFx2_ASAP7_75t_L g1623 ( 
.A(n_1553),
.Y(n_1623)
);

BUFx3_ASAP7_75t_L g1624 ( 
.A(n_1608),
.Y(n_1624)
);

HB1xp67_ASAP7_75t_L g1625 ( 
.A(n_1532),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1566),
.B(n_1539),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1530),
.A2(n_1503),
.B(n_1494),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1571),
.B(n_1459),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1555),
.B(n_1495),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1581),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1561),
.A2(n_1611),
.B1(n_1569),
.B2(n_1609),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1529),
.B(n_1438),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1568),
.B(n_1459),
.Y(n_1633)
);

AND2x4_ASAP7_75t_L g1634 ( 
.A(n_1553),
.B(n_1475),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1569),
.A2(n_1440),
.B1(n_1505),
.B2(n_1447),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1529),
.B(n_1527),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1558),
.B(n_1459),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1532),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1558),
.B(n_1457),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1608),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1609),
.A2(n_1493),
.B1(n_1461),
.B2(n_1447),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1549),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1554),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1568),
.B(n_1511),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1561),
.A2(n_1518),
.B(n_1525),
.Y(n_1645)
);

NOR2xp33_ASAP7_75t_L g1646 ( 
.A(n_1544),
.B(n_1493),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1647)
);

OAI221xp5_ASAP7_75t_L g1648 ( 
.A1(n_1569),
.A2(n_1493),
.B1(n_1505),
.B2(n_1440),
.C(n_1423),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1547),
.B(n_1461),
.Y(n_1649)
);

AOI221xp5_ASAP7_75t_L g1650 ( 
.A1(n_1609),
.A2(n_1424),
.B1(n_1525),
.B2(n_1413),
.C(n_1521),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1608),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1531),
.B(n_1521),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1554),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1531),
.B(n_1521),
.Y(n_1654)
);

OAI21xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1650),
.A2(n_1612),
.B(n_1556),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1614),
.B(n_1549),
.Y(n_1656)
);

OAI21xp33_ASAP7_75t_L g1657 ( 
.A1(n_1616),
.A2(n_1606),
.B(n_1542),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1614),
.B(n_1543),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_R g1660 ( 
.A(n_1646),
.B(n_1607),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1648),
.A2(n_1591),
.B1(n_1569),
.B2(n_1596),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1620),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1615),
.B(n_1565),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1615),
.B(n_1572),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1629),
.B(n_1550),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1648),
.A2(n_1591),
.B1(n_1596),
.B2(n_1593),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1629),
.B(n_1535),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_L g1668 ( 
.A(n_1616),
.B(n_1533),
.C(n_1588),
.D(n_1562),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1643),
.B(n_1545),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1635),
.B(n_1600),
.C(n_1605),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1647),
.Y(n_1671)
);

NAND3xp33_ASAP7_75t_L g1672 ( 
.A(n_1631),
.B(n_1593),
.C(n_1531),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_L g1673 ( 
.A(n_1641),
.B(n_1531),
.C(n_1600),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1631),
.A2(n_1635),
.B1(n_1588),
.B2(n_1646),
.C(n_1641),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1643),
.B(n_1598),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1628),
.B(n_1536),
.Y(n_1676)
);

NOR3xp33_ASAP7_75t_L g1677 ( 
.A(n_1650),
.B(n_1605),
.C(n_1548),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1649),
.B(n_1593),
.C(n_1582),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1618),
.A2(n_1601),
.B(n_1612),
.Y(n_1679)
);

AND2x2_ASAP7_75t_L g1680 ( 
.A(n_1617),
.B(n_1536),
.Y(n_1680)
);

AOI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1627),
.A2(n_1593),
.B1(n_1563),
.B2(n_1613),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1617),
.B(n_1537),
.Y(n_1682)
);

OAI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1645),
.A2(n_1597),
.B1(n_1556),
.B2(n_1541),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1537),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1633),
.B(n_1559),
.Y(n_1685)
);

OAI221xp5_ASAP7_75t_SL g1686 ( 
.A1(n_1645),
.A2(n_1563),
.B1(n_1556),
.B2(n_1597),
.C(n_1608),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1627),
.A2(n_1574),
.B1(n_1573),
.B2(n_1602),
.C(n_1592),
.Y(n_1687)
);

AOI221xp5_ASAP7_75t_L g1688 ( 
.A1(n_1627),
.A2(n_1592),
.B1(n_1560),
.B2(n_1599),
.C(n_1575),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1627),
.A2(n_1613),
.B1(n_1580),
.B2(n_1590),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1649),
.A2(n_1597),
.B1(n_1587),
.B2(n_1548),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1618),
.B(n_1538),
.C(n_1610),
.Y(n_1691)
);

OAI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1649),
.A2(n_1597),
.B1(n_1604),
.B2(n_1587),
.C(n_1608),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1652),
.B(n_1541),
.Y(n_1693)
);

OAI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1618),
.A2(n_1597),
.B1(n_1604),
.B2(n_1587),
.C(n_1546),
.Y(n_1694)
);

NOR3xp33_ASAP7_75t_SL g1695 ( 
.A(n_1644),
.B(n_1579),
.C(n_1540),
.Y(n_1695)
);

OAI221xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1621),
.A2(n_1599),
.B1(n_1604),
.B2(n_1575),
.C(n_1546),
.Y(n_1696)
);

NOR2xp67_ASAP7_75t_L g1697 ( 
.A(n_1630),
.B(n_1594),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1652),
.B(n_1576),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1632),
.B(n_1578),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1620),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1654),
.B(n_1564),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1627),
.B(n_1589),
.Y(n_1702)
);

AOI221xp5_ASAP7_75t_L g1703 ( 
.A1(n_1644),
.A2(n_1583),
.B1(n_1585),
.B2(n_1586),
.C(n_1584),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1624),
.A2(n_1546),
.B1(n_1610),
.B2(n_1580),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1634),
.B(n_1580),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1653),
.B(n_1595),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1658),
.B(n_1621),
.Y(n_1707)
);

OR2x6_ASAP7_75t_L g1708 ( 
.A(n_1679),
.B(n_1621),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1671),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1671),
.B(n_1653),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1662),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1658),
.B(n_1623),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1702),
.B(n_1625),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1662),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1663),
.B(n_1642),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1687),
.B(n_1625),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1673),
.A2(n_1601),
.B(n_1619),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1700),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1698),
.B(n_1638),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1700),
.Y(n_1720)
);

NAND2x1_ASAP7_75t_L g1721 ( 
.A(n_1697),
.B(n_1642),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1680),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1664),
.B(n_1642),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1701),
.B(n_1622),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1697),
.B(n_1624),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1680),
.Y(n_1726)
);

AND2x4_ASAP7_75t_L g1727 ( 
.A(n_1705),
.B(n_1624),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1667),
.B(n_1636),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1655),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1691),
.B(n_1624),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1706),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1684),
.B(n_1619),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1688),
.B(n_1626),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1684),
.B(n_1619),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1676),
.B(n_1626),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1659),
.B(n_1637),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1732),
.B(n_1693),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1718),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1709),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1732),
.B(n_1734),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1656),
.Y(n_1743)
);

INVxp67_ASAP7_75t_L g1744 ( 
.A(n_1716),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1709),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1713),
.B(n_1681),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1710),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1725),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1729),
.B(n_1655),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1718),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1707),
.B(n_1656),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1729),
.B(n_1681),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1710),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1711),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1721),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1713),
.B(n_1703),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1711),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1714),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1714),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1731),
.B(n_1682),
.Y(n_1761)
);

OAI21xp33_ASAP7_75t_L g1762 ( 
.A1(n_1733),
.A2(n_1657),
.B(n_1668),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1720),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1718),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1722),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1722),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1724),
.B(n_1689),
.Y(n_1767)
);

NAND3xp33_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1678),
.C(n_1657),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1728),
.B(n_1470),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1707),
.B(n_1640),
.Y(n_1770)
);

NAND2x1_ASAP7_75t_L g1771 ( 
.A(n_1725),
.B(n_1678),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1726),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1731),
.B(n_1685),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1735),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1736),
.B(n_1640),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1736),
.B(n_1651),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1736),
.B(n_1651),
.Y(n_1777)
);

NOR2x1_ASAP7_75t_L g1778 ( 
.A(n_1721),
.B(n_1672),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1738),
.B(n_1651),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1726),
.Y(n_1780)
);

AND2x4_ASAP7_75t_L g1781 ( 
.A(n_1748),
.B(n_1725),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1741),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1741),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1745),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.B(n_1728),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1745),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1754),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1754),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_L g1790 ( 
.A(n_1762),
.B(n_1737),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1757),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1762),
.B(n_1737),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1768),
.A2(n_1672),
.B1(n_1683),
.B2(n_1674),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1757),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1758),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1758),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1759),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1759),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1799)
);

INVxp67_ASAP7_75t_SL g1800 ( 
.A(n_1778),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1744),
.B(n_1712),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1760),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1749),
.B(n_1708),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1760),
.Y(n_1804)
);

INVxp67_ASAP7_75t_L g1805 ( 
.A(n_1756),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1763),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1763),
.Y(n_1807)
);

OR2x2_ASAP7_75t_L g1808 ( 
.A(n_1746),
.B(n_1733),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1752),
.B(n_1708),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1747),
.B(n_1716),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1752),
.B(n_1708),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1744),
.B(n_1712),
.Y(n_1813)
);

AO21x1_ASAP7_75t_SL g1814 ( 
.A1(n_1756),
.A2(n_1717),
.B(n_1719),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1765),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1755),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1752),
.B(n_1773),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1766),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1766),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1772),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1774),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1772),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1761),
.B(n_1715),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1780),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1761),
.B(n_1715),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1780),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1797),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1797),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1793),
.B(n_1768),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1782),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1781),
.B(n_1748),
.Y(n_1831)
);

INVxp67_ASAP7_75t_SL g1832 ( 
.A(n_1800),
.Y(n_1832)
);

OA21x2_ASAP7_75t_L g1833 ( 
.A1(n_1800),
.A2(n_1750),
.B(n_1740),
.Y(n_1833)
);

OAI221xp5_ASAP7_75t_L g1834 ( 
.A1(n_1805),
.A2(n_1771),
.B1(n_1778),
.B2(n_1708),
.C(n_1769),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1781),
.Y(n_1835)
);

AND3x2_ASAP7_75t_L g1836 ( 
.A(n_1805),
.B(n_1677),
.C(n_1725),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1817),
.B(n_1747),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1792),
.B(n_1458),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1783),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1781),
.B(n_1755),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1785),
.Y(n_1842)
);

CKINVDCx16_ASAP7_75t_R g1843 ( 
.A(n_1784),
.Y(n_1843)
);

NOR2xp33_ASAP7_75t_L g1844 ( 
.A(n_1790),
.B(n_1458),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1787),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1790),
.A2(n_1755),
.B(n_1730),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1784),
.B(n_1767),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1809),
.Y(n_1848)
);

INVx1_ASAP7_75t_SL g1849 ( 
.A(n_1809),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1801),
.B(n_1753),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1816),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1808),
.B(n_1767),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1799),
.B(n_1767),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1788),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1813),
.B(n_1739),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1799),
.B(n_1742),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1789),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1823),
.B(n_1774),
.Y(n_1858)
);

INVxp67_ASAP7_75t_L g1859 ( 
.A(n_1814),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1825),
.B(n_1810),
.Y(n_1860)
);

INVx1_ASAP7_75t_SL g1861 ( 
.A(n_1812),
.Y(n_1861)
);

INVxp67_ASAP7_75t_SL g1862 ( 
.A(n_1816),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1810),
.B(n_1774),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1812),
.Y(n_1864)
);

AOI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1829),
.A2(n_1771),
.B(n_1803),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1827),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1829),
.B(n_1803),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1835),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1828),
.Y(n_1869)
);

INVx1_ASAP7_75t_SL g1870 ( 
.A(n_1848),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1830),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1832),
.A2(n_1666),
.B(n_1661),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1843),
.B(n_1742),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1840),
.Y(n_1874)
);

AOI22xp5_ASAP7_75t_L g1875 ( 
.A1(n_1834),
.A2(n_1730),
.B1(n_1670),
.B2(n_1694),
.Y(n_1875)
);

AOI32xp33_ASAP7_75t_L g1876 ( 
.A1(n_1852),
.A2(n_1730),
.A3(n_1770),
.B1(n_1727),
.B2(n_1821),
.Y(n_1876)
);

AOI31xp33_ASAP7_75t_L g1877 ( 
.A1(n_1859),
.A2(n_1405),
.A3(n_1690),
.B(n_1730),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1842),
.Y(n_1878)
);

OAI21xp33_ASAP7_75t_L g1879 ( 
.A1(n_1852),
.A2(n_1686),
.B(n_1791),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1845),
.Y(n_1880)
);

AOI22xp5_ASAP7_75t_L g1881 ( 
.A1(n_1849),
.A2(n_1692),
.B1(n_1727),
.B2(n_1811),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1862),
.Y(n_1882)
);

CKINVDCx20_ASAP7_75t_R g1883 ( 
.A(n_1844),
.Y(n_1883)
);

OAI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1846),
.A2(n_1795),
.B(n_1794),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1833),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1854),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1847),
.B(n_1775),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1857),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1861),
.A2(n_1727),
.B1(n_1818),
.B2(n_1815),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1851),
.Y(n_1890)
);

NAND3xp33_ASAP7_75t_L g1891 ( 
.A(n_1836),
.B(n_1798),
.C(n_1796),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1864),
.B(n_1739),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1882),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1883),
.B(n_1844),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1890),
.Y(n_1895)
);

INVx1_ASAP7_75t_SL g1896 ( 
.A(n_1868),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1885),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1873),
.B(n_1847),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1870),
.B(n_1853),
.Y(n_1899)
);

NAND2xp33_ASAP7_75t_SL g1900 ( 
.A(n_1883),
.B(n_1660),
.Y(n_1900)
);

AOI22xp33_ASAP7_75t_L g1901 ( 
.A1(n_1879),
.A2(n_1853),
.B1(n_1831),
.B2(n_1860),
.Y(n_1901)
);

NOR2x1_ASAP7_75t_L g1902 ( 
.A(n_1891),
.B(n_1846),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1866),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1865),
.A2(n_1856),
.B1(n_1839),
.B2(n_1850),
.Y(n_1904)
);

INVxp67_ASAP7_75t_L g1905 ( 
.A(n_1867),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1887),
.B(n_1856),
.Y(n_1906)
);

INVxp67_ASAP7_75t_L g1907 ( 
.A(n_1884),
.Y(n_1907)
);

AOI22xp33_ASAP7_75t_SL g1908 ( 
.A1(n_1865),
.A2(n_1839),
.B1(n_1841),
.B2(n_1851),
.Y(n_1908)
);

NOR2x1p5_ASAP7_75t_SL g1909 ( 
.A(n_1885),
.B(n_1863),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1869),
.B(n_1841),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1841),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1889),
.B(n_1855),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1892),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1902),
.A2(n_1872),
.B(n_1875),
.Y(n_1914)
);

AOI221xp5_ASAP7_75t_L g1915 ( 
.A1(n_1907),
.A2(n_1872),
.B1(n_1886),
.B2(n_1888),
.C(n_1880),
.Y(n_1915)
);

AOI22xp5_ASAP7_75t_L g1916 ( 
.A1(n_1894),
.A2(n_1881),
.B1(n_1874),
.B2(n_1878),
.Y(n_1916)
);

NAND3xp33_ASAP7_75t_L g1917 ( 
.A(n_1908),
.B(n_1876),
.C(n_1877),
.Y(n_1917)
);

OAI21xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1904),
.A2(n_1838),
.B(n_1837),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1896),
.B(n_1819),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1893),
.B(n_1436),
.Y(n_1920)
);

AOI221xp5_ASAP7_75t_L g1921 ( 
.A1(n_1905),
.A2(n_1802),
.B1(n_1804),
.B2(n_1806),
.C(n_1807),
.Y(n_1921)
);

OAI221xp5_ASAP7_75t_L g1922 ( 
.A1(n_1901),
.A2(n_1858),
.B1(n_1695),
.B2(n_1821),
.C(n_1833),
.Y(n_1922)
);

AOI22xp5_ASAP7_75t_L g1923 ( 
.A1(n_1898),
.A2(n_1820),
.B1(n_1824),
.B2(n_1822),
.Y(n_1923)
);

AOI221x1_ASAP7_75t_L g1924 ( 
.A1(n_1900),
.A2(n_1826),
.B1(n_1764),
.B2(n_1740),
.C(n_1750),
.Y(n_1924)
);

NOR2xp33_ASAP7_75t_L g1925 ( 
.A(n_1900),
.B(n_1436),
.Y(n_1925)
);

OAI221xp5_ASAP7_75t_SL g1926 ( 
.A1(n_1899),
.A2(n_1675),
.B1(n_1669),
.B2(n_1723),
.C(n_1770),
.Y(n_1926)
);

OAI21xp33_ASAP7_75t_SL g1927 ( 
.A1(n_1898),
.A2(n_1743),
.B(n_1751),
.Y(n_1927)
);

NAND4xp75_ASAP7_75t_L g1928 ( 
.A(n_1920),
.B(n_1909),
.C(n_1897),
.D(n_1895),
.Y(n_1928)
);

NOR4xp25_ASAP7_75t_L g1929 ( 
.A(n_1914),
.B(n_1903),
.C(n_1897),
.D(n_1913),
.Y(n_1929)
);

INVxp33_ASAP7_75t_SL g1930 ( 
.A(n_1925),
.Y(n_1930)
);

NOR2x1_ASAP7_75t_L g1931 ( 
.A(n_1917),
.B(n_1910),
.Y(n_1931)
);

NOR2x1_ASAP7_75t_SL g1932 ( 
.A(n_1919),
.B(n_1903),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1916),
.Y(n_1933)
);

AND5x1_ASAP7_75t_L g1934 ( 
.A(n_1915),
.B(n_1909),
.C(n_1912),
.D(n_1913),
.E(n_1910),
.Y(n_1934)
);

NOR2x1_ASAP7_75t_L g1935 ( 
.A(n_1922),
.B(n_1910),
.Y(n_1935)
);

NOR2x1p5_ASAP7_75t_L g1936 ( 
.A(n_1918),
.B(n_1911),
.Y(n_1936)
);

NOR2x1_ASAP7_75t_L g1937 ( 
.A(n_1924),
.B(n_1911),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1923),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1926),
.B(n_1912),
.Y(n_1939)
);

AND4x1_ASAP7_75t_L g1940 ( 
.A(n_1931),
.B(n_1921),
.C(n_1906),
.D(n_1526),
.Y(n_1940)
);

NAND4xp75_ASAP7_75t_L g1941 ( 
.A(n_1937),
.B(n_1927),
.C(n_1906),
.D(n_1833),
.Y(n_1941)
);

NOR2xp33_ASAP7_75t_L g1942 ( 
.A(n_1930),
.B(n_1911),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1929),
.B(n_1773),
.Y(n_1943)
);

NAND4xp25_ASAP7_75t_L g1944 ( 
.A(n_1935),
.B(n_1696),
.C(n_1727),
.D(n_1526),
.Y(n_1944)
);

NOR3xp33_ASAP7_75t_L g1945 ( 
.A(n_1928),
.B(n_1468),
.C(n_1665),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1939),
.A2(n_1704),
.B(n_1779),
.C(n_1777),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1942),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1943),
.A2(n_1933),
.B1(n_1939),
.B2(n_1936),
.Y(n_1948)
);

AOI22xp5_ASAP7_75t_L g1949 ( 
.A1(n_1945),
.A2(n_1938),
.B1(n_1934),
.B2(n_1932),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1941),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1940),
.B(n_1775),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1946),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1944),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1951),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1947),
.B(n_1776),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1948),
.B(n_1750),
.C(n_1740),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1950),
.B(n_1468),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1952),
.Y(n_1958)
);

NOR2xp33_ASAP7_75t_L g1959 ( 
.A(n_1949),
.B(n_1468),
.Y(n_1959)
);

AOI211xp5_ASAP7_75t_L g1960 ( 
.A1(n_1959),
.A2(n_1954),
.B(n_1953),
.C(n_1958),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1955),
.B(n_1951),
.Y(n_1961)
);

AND2x4_ASAP7_75t_SL g1962 ( 
.A(n_1957),
.B(n_1413),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1956),
.B(n_1776),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1961),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1960),
.Y(n_1965)
);

NOR3xp33_ASAP7_75t_L g1966 ( 
.A(n_1964),
.B(n_1963),
.C(n_1962),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1966),
.B(n_1965),
.Y(n_1967)
);

OAI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1966),
.A2(n_1764),
.B1(n_1413),
.B2(n_1525),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_L g1969 ( 
.A(n_1967),
.B(n_1777),
.Y(n_1969)
);

INVxp67_ASAP7_75t_L g1970 ( 
.A(n_1968),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1969),
.B(n_1413),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1971),
.Y(n_1972)
);

AOI22xp33_ASAP7_75t_L g1973 ( 
.A1(n_1972),
.A2(n_1970),
.B1(n_1471),
.B2(n_1478),
.Y(n_1973)
);

OAI221xp5_ASAP7_75t_R g1974 ( 
.A1(n_1973),
.A2(n_1478),
.B1(n_1471),
.B2(n_1408),
.C(n_1423),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1424),
.B(n_1521),
.C(n_1507),
.Y(n_1975)
);


endmodule