module fake_jpeg_2714_n_431 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_431);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_431;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_3),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_41),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_42),
.B(n_45),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_46),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_57),
.B(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_68),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_0),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_16),
.B(n_8),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_16),
.B(n_8),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_78),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_76),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_31),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_0),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_17),
.B(n_15),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_80),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_77),
.A2(n_35),
.B1(n_28),
.B2(n_36),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_81),
.A2(n_86),
.B1(n_117),
.B2(n_61),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_36),
.B1(n_28),
.B2(n_35),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_83),
.A2(n_115),
.B1(n_119),
.B2(n_54),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_40),
.B1(n_24),
.B2(n_32),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_94),
.B1(n_117),
.B2(n_88),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_39),
.B1(n_17),
.B2(n_37),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_91),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_66),
.A2(n_29),
.B1(n_37),
.B2(n_32),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_30),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_40),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_1),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_49),
.B(n_24),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_123),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_44),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_30),
.B1(n_25),
.B2(n_9),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_44),
.A2(n_30),
.B1(n_14),
.B2(n_13),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_50),
.B(n_14),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_80),
.B1(n_70),
.B2(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_126),
.A2(n_144),
.B1(n_164),
.B2(n_124),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_81),
.A2(n_59),
.B1(n_55),
.B2(n_58),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_127),
.A2(n_146),
.B1(n_153),
.B2(n_118),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_107),
.B(n_72),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_131),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_129),
.Y(n_173)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_134),
.B(n_145),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_44),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_136),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_87),
.A2(n_61),
.B(n_63),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_137),
.A2(n_167),
.B(n_96),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_138),
.B(n_98),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_92),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_84),
.B(n_41),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_143),
.Y(n_183)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_53),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_61),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_112),
.A2(n_43),
.B1(n_75),
.B2(n_64),
.Y(n_146)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_148),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_87),
.A2(n_69),
.B1(n_52),
.B2(n_60),
.Y(n_149)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_150),
.B(n_156),
.Y(n_176)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_86),
.A2(n_76),
.B1(n_51),
.B2(n_74),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

OR2x2_ASAP7_75t_SL g155 ( 
.A(n_107),
.B(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_155),
.B(n_168),
.Y(n_174)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_158),
.Y(n_187)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_94),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_160),
.Y(n_201)
);

NAND3xp33_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_121),
.C(n_102),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_92),
.B(n_1),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_166),
.Y(n_200)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_100),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_163),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_85),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_135),
.B1(n_145),
.B2(n_155),
.Y(n_197)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_96),
.B(n_101),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_185),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_177),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_179),
.A2(n_189),
.B1(n_190),
.B2(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_111),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_98),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_186),
.B(n_161),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_143),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_188),
.B(n_192),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_124),
.B1(n_97),
.B2(n_101),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_143),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_93),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_138),
.A2(n_93),
.B1(n_100),
.B2(n_116),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_126),
.B1(n_153),
.B2(n_164),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_195),
.A2(n_203),
.B1(n_148),
.B2(n_133),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_156),
.B1(n_129),
.B2(n_157),
.Y(n_225)
);

OAI22x1_ASAP7_75t_L g199 ( 
.A1(n_137),
.A2(n_111),
.B1(n_125),
.B2(n_105),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_199),
.A2(n_152),
.B1(n_62),
.B2(n_132),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_161),
.A2(n_122),
.B1(n_110),
.B2(n_116),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_130),
.B(n_110),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_162),
.C(n_158),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_151),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_209),
.B(n_223),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_174),
.A2(n_150),
.B(n_167),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_211),
.A2(n_229),
.B(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_168),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_172),
.C(n_181),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_193),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_163),
.B1(n_122),
.B2(n_154),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_221),
.B1(n_228),
.B2(n_230),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_236),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_190),
.Y(n_259)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_171),
.B(n_176),
.Y(n_223)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_224),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_226),
.Y(n_266)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_122),
.B1(n_142),
.B2(n_111),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_174),
.A2(n_147),
.B(n_136),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_179),
.A2(n_166),
.B1(n_125),
.B2(n_105),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_238),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_196),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_178),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_235),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_1),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_240),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_13),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_241),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_177),
.A2(n_30),
.B(n_13),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_242),
.A2(n_200),
.B(n_201),
.Y(n_265)
);

CKINVDCx11_ASAP7_75t_R g243 ( 
.A(n_191),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_243),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_189),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_244),
.A2(n_203),
.B1(n_205),
.B2(n_198),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_182),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_194),
.B1(n_205),
.B2(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_183),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_250),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_264),
.B1(n_267),
.B2(n_268),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_206),
.B1(n_192),
.B2(n_188),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_258),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_215),
.B(n_172),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_262),
.C(n_277),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_231),
.A2(n_216),
.B1(n_232),
.B2(n_226),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_216),
.A2(n_227),
.B1(n_220),
.B2(n_213),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_213),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_207),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_199),
.B(n_184),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_224),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_221),
.A2(n_238),
.B1(n_220),
.B2(n_234),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_223),
.A2(n_170),
.B1(n_185),
.B2(n_200),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_217),
.A2(n_199),
.B1(n_190),
.B2(n_200),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_263),
.B1(n_251),
.B2(n_273),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_241),
.A2(n_178),
.B1(n_198),
.B2(n_202),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_237),
.B1(n_235),
.B2(n_212),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_175),
.C(n_208),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_246),
.B(n_208),
.C(n_173),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_235),
.C(n_191),
.Y(n_307)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_255),
.A2(n_273),
.B1(n_261),
.B2(n_257),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_291),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_211),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_262),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_294),
.A2(n_302),
.B1(n_303),
.B2(n_268),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_296),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_249),
.B(n_209),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_240),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_298),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_266),
.B(n_210),
.Y(n_298)
);

A2O1A1Ixp33_ASAP7_75t_R g299 ( 
.A1(n_260),
.A2(n_210),
.B(n_222),
.C(n_225),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_299),
.B(n_300),
.Y(n_333)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_276),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_301),
.A2(n_309),
.B(n_271),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_251),
.A2(n_244),
.B1(n_242),
.B2(n_230),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_273),
.A2(n_228),
.B1(n_235),
.B2(n_243),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_307),
.C(n_259),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_278),
.B(n_245),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_306),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_275),
.B(n_173),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_278),
.B(n_233),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_274),
.B(n_298),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_313),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_279),
.B(n_258),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_286),
.A2(n_257),
.B1(n_261),
.B2(n_279),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_314),
.A2(n_322),
.B1(n_325),
.B2(n_328),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_323),
.C(n_334),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_320),
.B1(n_284),
.B2(n_283),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_318),
.B(n_307),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_267),
.B1(n_253),
.B2(n_252),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_287),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_326),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_286),
.A2(n_252),
.B1(n_264),
.B2(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_277),
.C(n_248),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_295),
.A2(n_301),
.B1(n_310),
.B2(n_309),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_287),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_294),
.A2(n_299),
.B1(n_305),
.B2(n_300),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_292),
.B(n_250),
.C(n_281),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_302),
.A2(n_274),
.B1(n_280),
.B2(n_270),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_313),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_338),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g338 ( 
.A(n_318),
.B(n_303),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_308),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_332),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_326),
.B(n_291),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_342),
.B(n_358),
.Y(n_364)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_343),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_327),
.A2(n_288),
.B1(n_290),
.B2(n_289),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_345),
.A2(n_349),
.B1(n_350),
.B2(n_357),
.Y(n_368)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_348),
.B(n_354),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_324),
.B(n_224),
.Y(n_351)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_353),
.C(n_330),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_316),
.B(n_270),
.C(n_202),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_355),
.C(n_339),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_333),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_336),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_323),
.B(n_196),
.C(n_233),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_335),
.A2(n_290),
.B1(n_272),
.B2(n_10),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_272),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_346),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_359),
.B(n_366),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_354),
.A2(n_336),
.B1(n_328),
.B2(n_317),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_371),
.Y(n_385)
);

AOI321xp33_ASAP7_75t_L g361 ( 
.A1(n_338),
.A2(n_331),
.A3(n_312),
.B1(n_337),
.B2(n_344),
.C(n_342),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_361),
.A2(n_372),
.B(n_12),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_SL g363 ( 
.A(n_346),
.B(n_325),
.C(n_314),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_363),
.B(n_367),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_365),
.B(n_352),
.C(n_355),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_350),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g371 ( 
.A1(n_344),
.A2(n_333),
.B(n_322),
.Y(n_371)
);

A2O1A1O1Ixp25_ASAP7_75t_L g372 ( 
.A1(n_356),
.A2(n_324),
.B(n_320),
.C(n_332),
.D(n_329),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_330),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_373),
.B(n_340),
.Y(n_382)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_375),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_356),
.A2(n_319),
.B1(n_329),
.B2(n_12),
.Y(n_376)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_376),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_377),
.B(n_380),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_365),
.B(n_358),
.C(n_339),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_347),
.C(n_319),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_383),
.B(n_388),
.C(n_390),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_11),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_369),
.B(n_11),
.Y(n_386)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_364),
.B(n_2),
.C(n_4),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_389),
.A2(n_370),
.B(n_372),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_2),
.C(n_5),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_385),
.B(n_362),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_391),
.B(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_381),
.A2(n_360),
.B1(n_371),
.B2(n_374),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_395),
.Y(n_404)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_394),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_363),
.C(n_368),
.Y(n_395)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_378),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_396),
.B(n_403),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_385),
.A2(n_376),
.B1(n_362),
.B2(n_361),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_387),
.A2(n_379),
.B1(n_377),
.B2(n_388),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_399),
.B(n_6),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_12),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_2),
.B(n_5),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_2),
.C(n_5),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_402),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_401),
.A2(n_7),
.B(n_5),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_406),
.A2(n_407),
.B1(n_411),
.B2(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_395),
.B(n_6),
.C(n_7),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_408),
.B(n_409),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_398),
.B(n_6),
.C(n_7),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_393),
.B(n_400),
.Y(n_411)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_415),
.Y(n_424)
);

BUFx24_ASAP7_75t_SL g416 ( 
.A(n_404),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_416),
.B(n_420),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_413),
.B(n_392),
.C(n_391),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_417),
.B(n_418),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_392),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_412),
.C(n_411),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_403),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_419),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_421),
.B(n_425),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_423),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_424),
.B(n_422),
.Y(n_428)
);

A2O1A1Ixp33_ASAP7_75t_L g429 ( 
.A1(n_428),
.A2(n_426),
.B(n_405),
.C(n_414),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_429),
.B(n_6),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_430),
.B(n_7),
.Y(n_431)
);


endmodule