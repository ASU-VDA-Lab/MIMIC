module fake_aes_2959_n_22 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_22);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_22;
wire n_20;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_4), .Y(n_9) );
CKINVDCx20_ASAP7_75t_R g10 ( .A(n_5), .Y(n_10) );
INVx2_ASAP7_75t_SL g11 ( .A(n_4), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
BUFx2_ASAP7_75t_L g14 ( .A(n_11), .Y(n_14) );
A2O1A1Ixp33_ASAP7_75t_SL g15 ( .A1(n_13), .A2(n_11), .B(n_9), .C(n_10), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_14), .B(n_13), .Y(n_16) );
OR2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_14), .Y(n_17) );
OAI21xp5_ASAP7_75t_SL g18 ( .A1(n_17), .A2(n_16), .B(n_12), .Y(n_18) );
AOI22xp33_ASAP7_75t_SL g19 ( .A1(n_18), .A2(n_15), .B1(n_1), .B2(n_3), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_19), .Y(n_20) );
OAI322xp33_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_0), .A3(n_1), .B1(n_3), .B2(n_5), .C1(n_6), .C2(n_7), .Y(n_21) );
AOI22xp33_ASAP7_75t_R g22 ( .A1(n_21), .A2(n_0), .B1(n_6), .B2(n_8), .Y(n_22) );
endmodule