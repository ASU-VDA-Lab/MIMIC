module fake_jpeg_11240_n_329 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_49),
.Y(n_64)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_18),
.Y(n_56)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_56),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_36),
.B1(n_25),
.B2(n_27),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_58),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_0),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_38),
.B(n_41),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_60),
.Y(n_70)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_67),
.B(n_68),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_36),
.B1(n_30),
.B2(n_19),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_71),
.B(n_74),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_37),
.B1(n_35),
.B2(n_38),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_73),
.A2(n_99),
.B1(n_28),
.B2(n_35),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_83),
.Y(n_126)
);

BUFx2_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_89),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_56),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_46),
.B(n_31),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_33),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_51),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_41),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_27),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_97),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_35),
.B1(n_38),
.B2(n_32),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_22),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_104),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_42),
.Y(n_132)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_101),
.B1(n_83),
.B2(n_89),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_120),
.B1(n_131),
.B2(n_146),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_115),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_117),
.A2(n_134),
.B1(n_144),
.B2(n_65),
.Y(n_171)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_58),
.B1(n_42),
.B2(n_29),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_145),
.B(n_93),
.Y(n_157)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_80),
.B(n_30),
.CI(n_2),
.CON(n_124),
.SN(n_124)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_124),
.B(n_4),
.Y(n_172)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_92),
.A2(n_58),
.B1(n_42),
.B2(n_29),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_75),
.B1(n_66),
.B2(n_105),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_107),
.A2(n_34),
.B1(n_19),
.B2(n_24),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_132),
.B(n_9),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_77),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_107),
.A2(n_29),
.B1(n_21),
.B2(n_24),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_19),
.B1(n_26),
.B2(n_18),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g161 ( 
.A1(n_137),
.A2(n_75),
.B1(n_66),
.B2(n_85),
.Y(n_161)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_77),
.A2(n_21),
.B1(n_81),
.B2(n_79),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_64),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_166),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_161),
.B1(n_171),
.B2(n_120),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_157),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_126),
.A2(n_70),
.B(n_81),
.C(n_79),
.Y(n_158)
);

O2A1O1Ixp33_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_118),
.B(n_122),
.C(n_12),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_72),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_178),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_78),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_174),
.Y(n_185)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_165),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_112),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_126),
.B(n_93),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_167),
.A2(n_129),
.B(n_128),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_85),
.C(n_72),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_168),
.B(n_137),
.C(n_119),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_169),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_70),
.B1(n_105),
.B2(n_65),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_138),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_172),
.A2(n_124),
.B(n_141),
.C(n_115),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_135),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_176),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_141),
.B(n_16),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_126),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_122),
.B1(n_11),
.B2(n_13),
.Y(n_211)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_121),
.Y(n_180)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_180),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_188),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g186 ( 
.A1(n_159),
.A2(n_132),
.A3(n_124),
.B1(n_143),
.B2(n_117),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_186),
.B(n_206),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_141),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_197),
.B(n_157),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_162),
.B1(n_161),
.B2(n_153),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_202),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_139),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_204),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_167),
.A2(n_111),
.B(n_137),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_137),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_210),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_212),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_15),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_10),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_214),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_217),
.A2(n_237),
.B(n_204),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_196),
.B(n_153),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_207),
.C(n_191),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_224),
.B1(n_211),
.B2(n_208),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_192),
.A2(n_162),
.B1(n_172),
.B2(n_161),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_189),
.A2(n_158),
.B(n_176),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_239),
.B(n_190),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_161),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_181),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_232),
.Y(n_253)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_230),
.Y(n_251)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_201),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_166),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_231),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_195),
.B(n_179),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_235),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_147),
.B(n_154),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_185),
.B(n_154),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_238),
.B(n_205),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_147),
.B(n_156),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_182),
.B1(n_206),
.B2(n_187),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_254),
.B1(n_223),
.B2(n_227),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_245),
.B(n_226),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_232),
.A2(n_208),
.B1(n_183),
.B2(n_200),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_257),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_203),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_250),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_219),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_227),
.B(n_203),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_255),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_205),
.B1(n_194),
.B2(n_213),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_194),
.B1(n_213),
.B2(n_207),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_258),
.A2(n_217),
.B(n_237),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_268),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_272),
.B(n_245),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_251),
.Y(n_266)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_270),
.Y(n_283)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_243),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_216),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_241),
.B(n_228),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g288 ( 
.A(n_273),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_254),
.A2(n_223),
.B1(n_239),
.B2(n_220),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_244),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_250),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_261),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_253),
.B1(n_215),
.B2(n_247),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_285),
.B1(n_273),
.B2(n_265),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_249),
.C(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_291),
.C(n_246),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_269),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_253),
.B1(n_242),
.B2(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_264),
.B(n_274),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_248),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_287),
.A2(n_262),
.B(n_215),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_235),
.C(n_218),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g292 ( 
.A(n_290),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_299),
.B1(n_288),
.B2(n_229),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_300),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_263),
.B1(n_221),
.B2(n_266),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_296),
.A2(n_298),
.B1(n_287),
.B2(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_289),
.A2(n_276),
.B1(n_275),
.B2(n_270),
.Y(n_299)
);

OAI21x1_ASAP7_75t_SL g300 ( 
.A1(n_283),
.A2(n_218),
.B(n_268),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_284),
.B(n_246),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_302),
.C(n_282),
.Y(n_307)
);

OA21x2_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_285),
.B(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_304),
.B1(n_295),
.B2(n_233),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_297),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_310),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_214),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_279),
.C(n_301),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_315),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_286),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_313),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_303),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_310),
.Y(n_320)
);

OAI21x1_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_236),
.B(n_191),
.Y(n_317)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_236),
.A3(n_313),
.B1(n_198),
.B2(n_155),
.C1(n_314),
.C2(n_307),
.Y(n_319)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_155),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_324),
.C(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_323),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_11),
.B(n_14),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_11),
.Y(n_329)
);


endmodule