module fake_jpeg_8435_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_41),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_38),
.B(n_44),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_19),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_48),
.Y(n_85)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_31),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_19),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_52),
.B(n_60),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_30),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_64),
.B(n_66),
.Y(n_94)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_69),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_58),
.B1(n_59),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_22),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_45),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_48),
.B(n_25),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_1),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_47),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_41),
.B1(n_25),
.B2(n_16),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_20),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_81),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_90),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_62),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_17),
.Y(n_103)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_95),
.A2(n_108),
.B1(n_90),
.B2(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_98),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_24),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_68),
.A2(n_32),
.B(n_24),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_102),
.B(n_114),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_2),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_106),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_39),
.C(n_40),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_39),
.C(n_81),
.Y(n_132)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_65),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_82),
.A2(n_40),
.B1(n_36),
.B2(n_21),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_33),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_99),
.B1(n_107),
.B2(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_129),
.B1(n_131),
.B2(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_109),
.Y(n_120)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_69),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_123),
.Y(n_149)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_115),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_71),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_92),
.B1(n_64),
.B2(n_75),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_101),
.C(n_100),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_112),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_17),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_113),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_97),
.A2(n_88),
.B1(n_32),
.B2(n_87),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_96),
.B1(n_32),
.B2(n_114),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_138),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_139),
.A2(n_140),
.B(n_144),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_103),
.B(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_117),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_102),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_150),
.C(n_152),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_132),
.B(n_117),
.C(n_122),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_126),
.A2(n_114),
.B(n_101),
.Y(n_154)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_154),
.A2(n_135),
.B1(n_120),
.B2(n_125),
.C(n_32),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_33),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_118),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

AO221x1_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_136),
.B1(n_83),
.B2(n_96),
.C(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_162),
.Y(n_172)
);

AO221x1_ASAP7_75t_L g162 ( 
.A1(n_141),
.A2(n_131),
.B1(n_119),
.B2(n_121),
.C(n_127),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_142),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_165),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_139),
.Y(n_176)
);

OAI321xp33_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_28),
.A3(n_23),
.B1(n_10),
.B2(n_6),
.C(n_7),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_151),
.A3(n_149),
.B1(n_153),
.B2(n_155),
.C1(n_147),
.C2(n_12),
.Y(n_177)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_168),
.B(n_169),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_146),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_152),
.C(n_154),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_174),
.C(n_179),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_144),
.C(n_140),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_167),
.B1(n_159),
.B2(n_169),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_175),
.A2(n_178),
.B1(n_23),
.B2(n_17),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_176),
.A2(n_160),
.B(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_156),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_143),
.B1(n_147),
.B2(n_28),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_28),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_182),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_180),
.B(n_159),
.Y(n_183)
);

BUFx24_ASAP7_75t_SL g189 ( 
.A(n_183),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_185),
.A2(n_176),
.B1(n_179),
.B2(n_174),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_186),
.A2(n_172),
.B1(n_170),
.B2(n_4),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_7),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_188),
.C(n_171),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_173),
.B(n_8),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_192),
.B(n_194),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_193),
.B(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_186),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_184),
.C(n_8),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_196),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_184),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_190),
.C(n_13),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_202),
.C(n_3),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_2),
.C(n_3),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_197),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_3),
.Y(n_206)
);


endmodule