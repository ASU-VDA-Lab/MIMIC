module fake_jpeg_29448_n_117 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_117);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_117;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_34),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_29),
.B(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_23),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_38),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_18),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_13),
.Y(n_48)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_29),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_54),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_67),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_30),
.C(n_33),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_60),
.C(n_64),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_31),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_22),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_25),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_47),
.A2(n_15),
.B1(n_17),
.B2(n_23),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_47),
.B(n_39),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_17),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_50),
.C(n_49),
.Y(n_84)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_76),
.B1(n_81),
.B2(n_68),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_64),
.A2(n_47),
.B1(n_40),
.B2(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_64),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_38),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_47),
.B(n_54),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_59),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_43),
.B1(n_52),
.B2(n_40),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_49),
.Y(n_93)
);

FAx1_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_86),
.CI(n_88),
.CON(n_97),
.SN(n_97)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_69),
.C(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_91),
.B1(n_38),
.B2(n_71),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_67),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_74),
.A2(n_52),
.B1(n_66),
.B2(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_84),
.B(n_81),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_97),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_88),
.A2(n_80),
.B1(n_73),
.B2(n_75),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_96),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_104)
);

OAI321xp33_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_38),
.A3(n_71),
.B1(n_24),
.B2(n_39),
.C(n_7),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_7),
.B1(n_8),
.B2(n_93),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_94),
.C(n_8),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_105),
.Y(n_111)
);

BUFx24_ASAP7_75t_SL g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_94),
.C(n_95),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_99),
.B(n_98),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_110),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_104),
.B(n_98),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_101),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_113),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_109),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_113),
.C(n_114),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_116),
.Y(n_117)
);


endmodule