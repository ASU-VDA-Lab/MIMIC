module fake_netlist_6_1565_n_1172 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1172);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1172;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_760;
wire n_741;
wire n_209;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_208;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_168;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_1164;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_180;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1160;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1074;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_955;
wire n_337;
wire n_865;
wire n_1138;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_181;
wire n_1127;
wire n_182;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_963;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_1120;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_1139;
wire n_198;
wire n_300;
wire n_718;
wire n_179;
wire n_248;
wire n_222;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_923;
wire n_504;
wire n_1078;
wire n_314;
wire n_1140;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_948;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_977;
wire n_945;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_761;
wire n_428;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_167;
wire n_631;
wire n_174;
wire n_720;
wire n_758;
wire n_516;
wire n_842;
wire n_525;
wire n_1163;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_886;
wire n_448;
wire n_953;
wire n_1017;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_220;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_196;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1041;
wire n_279;
wire n_686;
wire n_796;
wire n_1000;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_719;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_936;
wire n_184;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_216;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_683;
wire n_811;
wire n_630;
wire n_312;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_175;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_1155;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_1053;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_199;
wire n_1167;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_420;
wire n_1153;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_1165;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_1157;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_515;
wire n_434;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1154;
wire n_177;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_170;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_664;
wire n_194;
wire n_171;
wire n_949;
wire n_678;
wire n_192;
wire n_169;
wire n_1007;
wire n_649;
wire n_855;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_139),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_96),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_49),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_149),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_81),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_43),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_17),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_84),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_27),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_109),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_4),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_10),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_39),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_76),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_37),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_10),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_163),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_24),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_0),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_164),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_83),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_85),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_33),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_19),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_146),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_56),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_5),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_115),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_99),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_154),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_117),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_67),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_143),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_102),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_93),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_134),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_17),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_80),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_42),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_46),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_78),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_166),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_168),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_173),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_178),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_186),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_187),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_192),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_198),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_199),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_200),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_203),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_201),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_172),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_171),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_217),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_204),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_246),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_247),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_225),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_249),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_251),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_229),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_230),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_232),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_233),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_234),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_228),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_235),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_239),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_245),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_241),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_242),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_253),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_248),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_238),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_238),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_243),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_243),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_224),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_224),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_247),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_247),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_224),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_224),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_244),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_224),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_290),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_272),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_277),
.Y(n_309)
);

INVxp67_ASAP7_75t_SL g310 ( 
.A(n_255),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_278),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_259),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_260),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_288),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_300),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_257),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_280),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_282),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_299),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_265),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_183),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_258),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

INVxp67_ASAP7_75t_SL g337 ( 
.A(n_270),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_279),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_256),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_291),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_292),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_256),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_268),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_271),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_267),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_296),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_269),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_314),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_316),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_321),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_333),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_314),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_328),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_335),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_328),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_327),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_313),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_322),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_335),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_319),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_315),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_320),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_344),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_320),
.Y(n_376)
);

INVxp33_ASAP7_75t_SL g377 ( 
.A(n_319),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_346),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_R g380 ( 
.A(n_350),
.B(n_274),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_308),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_317),
.Y(n_383)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_348),
.B(n_296),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_350),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_309),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_345),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_311),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_345),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_297),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_323),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_351),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_306),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_359),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_390),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_370),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_371),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_347),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

INVxp33_ASAP7_75t_SL g410 ( 
.A(n_380),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_376),
.B(n_338),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_341),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_388),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_342),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_354),
.Y(n_416)
);

CKINVDCx6p67_ASAP7_75t_R g417 ( 
.A(n_363),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_391),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_397),
.A2(n_305),
.B(n_334),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

OAI22x1_ASAP7_75t_R g423 ( 
.A1(n_372),
.A2(n_297),
.B1(n_301),
.B2(n_302),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_398),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

NAND2x1p5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_351),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_383),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_361),
.B(n_310),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_361),
.B(n_325),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_369),
.B(n_331),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_377),
.B(n_343),
.Y(n_438)
);

AND2x2_ASAP7_75t_SL g439 ( 
.A(n_377),
.B(n_221),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_355),
.B(n_332),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_356),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

AND2x2_ASAP7_75t_SL g444 ( 
.A(n_362),
.B(n_210),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_364),
.B(n_352),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_385),
.Y(n_447)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_385),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_372),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_374),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_276),
.Y(n_452)
);

CKINVDCx6p67_ASAP7_75t_R g453 ( 
.A(n_375),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_358),
.B(n_281),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_358),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_372),
.A2(n_218),
.B1(n_214),
.B2(n_195),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_365),
.B(n_340),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_358),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_358),
.B(n_284),
.Y(n_461)
);

OA21x2_ASAP7_75t_L g462 ( 
.A1(n_357),
.A2(n_169),
.B(n_167),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_358),
.Y(n_463)
);

AND2x6_ASAP7_75t_L g464 ( 
.A(n_358),
.B(n_349),
.Y(n_464)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_390),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_358),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_357),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_365),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_358),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_365),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_358),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_358),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_358),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_358),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_358),
.B(n_285),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_358),
.Y(n_478)
);

INVx6_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_358),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_358),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_358),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_358),
.B(n_286),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_358),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_406),
.B(n_349),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_471),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_400),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_484),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_439),
.A2(n_339),
.B1(n_337),
.B2(n_304),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_405),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_418),
.B(n_287),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_406),
.B(n_301),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_438),
.B(n_302),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_407),
.B(n_304),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_407),
.B(n_195),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_414),
.B(n_214),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_401),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_414),
.B(n_218),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_472),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_176),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_403),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_429),
.B(n_180),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_457),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_460),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_467),
.Y(n_510)
);

BUFx8_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_189),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_409),
.B(n_210),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_409),
.B(n_182),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_416),
.B(n_184),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_422),
.B(n_172),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_478),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_480),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_433),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_456),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_422),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_425),
.B(n_223),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_504),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_495),
.A2(n_439),
.B1(n_479),
.B2(n_465),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_505),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_511),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_507),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_511),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_511),
.Y(n_534)
);

AOI21x1_ASAP7_75t_L g535 ( 
.A1(n_485),
.A2(n_421),
.B(n_462),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_523),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_523),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_493),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_489),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_506),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_493),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_486),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_502),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_512),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_488),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_492),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_509),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_492),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_490),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_492),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_R g552 ( 
.A(n_506),
.B(n_424),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_514),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_494),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_494),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_488),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_499),
.B(n_425),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_496),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_518),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_510),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_526),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_497),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_501),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_515),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_424),
.Y(n_565)
);

NAND3xp33_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_458),
.C(n_402),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_563),
.B(n_444),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_556),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_536),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_527),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_550),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_528),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g573 ( 
.A(n_562),
.B(n_402),
.C(n_424),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_558),
.B(n_452),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_454),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_537),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_555),
.B(n_408),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_540),
.B(n_451),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_530),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_532),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_546),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_548),
.Y(n_582)
);

AO21x2_ASAP7_75t_L g583 ( 
.A1(n_535),
.A2(n_513),
.B(n_503),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_538),
.B(n_454),
.Y(n_584)
);

NAND2xp33_ASAP7_75t_L g585 ( 
.A(n_539),
.B(n_429),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_560),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_541),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_564),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_542),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_557),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_543),
.Y(n_592)
);

AOI21x1_ASAP7_75t_L g593 ( 
.A1(n_553),
.A2(n_421),
.B(n_462),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_556),
.Y(n_594)
);

BUFx4f_ASAP7_75t_L g595 ( 
.A(n_556),
.Y(n_595)
);

NOR2x1p5_ASAP7_75t_L g596 ( 
.A(n_531),
.B(n_453),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_545),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_545),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_544),
.B(n_410),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_553),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_553),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_540),
.A2(n_444),
.B1(n_513),
.B2(n_503),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_547),
.B(n_415),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_551),
.B(n_450),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_549),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_534),
.B(n_455),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_561),
.B(n_461),
.Y(n_609)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_559),
.A2(n_445),
.B1(n_479),
.B2(n_465),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_561),
.B(n_477),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_538),
.Y(n_612)
);

INVx2_ASAP7_75t_SL g613 ( 
.A(n_541),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_550),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_559),
.B(n_441),
.C(n_483),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_561),
.B(n_427),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_538),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_556),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_554),
.B(n_434),
.Y(n_619)
);

INVx5_ASAP7_75t_L g620 ( 
.A(n_556),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_554),
.B(n_434),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_527),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_536),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_561),
.B(n_427),
.Y(n_624)
);

INVx4_ASAP7_75t_L g625 ( 
.A(n_536),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_550),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_531),
.Y(n_627)
);

INVxp67_ASAP7_75t_SL g628 ( 
.A(n_550),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_536),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_550),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_550),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_L g634 ( 
.A(n_552),
.B(n_429),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_561),
.B(n_456),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_561),
.B(n_426),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_527),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_527),
.Y(n_638)
);

INVxp33_ASAP7_75t_SL g639 ( 
.A(n_559),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_561),
.B(n_466),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_527),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_556),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_559),
.B(n_446),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_561),
.B(n_466),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_628),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_636),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_612),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_574),
.B(n_446),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_574),
.B(n_443),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_586),
.A2(n_451),
.B1(n_448),
.B2(n_443),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_612),
.Y(n_651)
);

OAI21xp33_ASAP7_75t_SL g652 ( 
.A1(n_603),
.A2(n_525),
.B(n_491),
.Y(n_652)
);

INVx5_ASAP7_75t_L g653 ( 
.A(n_568),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_603),
.A2(n_449),
.B1(n_447),
.B2(n_426),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_615),
.A2(n_445),
.B1(n_442),
.B2(n_465),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_448),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_595),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_580),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_617),
.Y(n_659)
);

NOR2x1p5_ASAP7_75t_L g660 ( 
.A(n_566),
.B(n_573),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_604),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_570),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_587),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_617),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_591),
.B(n_503),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_448),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_584),
.B(n_609),
.Y(n_668)
);

AND2x2_ASAP7_75t_SL g669 ( 
.A(n_634),
.B(n_440),
.Y(n_669)
);

INVx4_ASAP7_75t_L g670 ( 
.A(n_569),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_584),
.Y(n_671)
);

OAI21xp33_ASAP7_75t_L g672 ( 
.A1(n_586),
.A2(n_567),
.B(n_611),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_568),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_601),
.B(n_488),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_579),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_595),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_607),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_581),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_568),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_582),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_568),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_577),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_611),
.B(n_608),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_575),
.B(n_448),
.Y(n_684)
);

INVxp67_ASAP7_75t_SL g685 ( 
.A(n_628),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_597),
.Y(n_686)
);

BUFx6f_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_589),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_613),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_607),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_608),
.B(n_429),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_622),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_625),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_632),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_575),
.B(n_520),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_576),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_637),
.Y(n_697)
);

AND2x6_ASAP7_75t_L g698 ( 
.A(n_602),
.B(n_488),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_520),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_635),
.B(n_640),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_643),
.B(n_440),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_620),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_598),
.B(n_487),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_635),
.B(n_517),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_R g705 ( 
.A(n_565),
.B(n_440),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_638),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_641),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_623),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_625),
.B(n_430),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_590),
.Y(n_710)
);

OAI21xp33_ASAP7_75t_L g711 ( 
.A1(n_616),
.A2(n_413),
.B(n_411),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_600),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_614),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_629),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_614),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_571),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_592),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_631),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_619),
.B(n_519),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_626),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_651),
.B(n_616),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_719),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_662),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_684),
.B(n_621),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_659),
.B(n_624),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_701),
.B(n_624),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_658),
.B(n_605),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_675),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_687),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_678),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_645),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_663),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_711),
.B(n_640),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_677),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_648),
.B(n_643),
.Y(n_738)
);

INVx1_ASAP7_75t_SL g739 ( 
.A(n_646),
.Y(n_739)
);

NAND3x1_ASAP7_75t_L g740 ( 
.A(n_668),
.B(n_600),
.C(n_610),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_680),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_692),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_685),
.B(n_644),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_666),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_683),
.A2(n_644),
.B1(n_599),
.B2(n_606),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_645),
.B(n_583),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_691),
.A2(n_700),
.B1(n_706),
.B2(n_697),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_688),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_694),
.Y(n_749)
);

NAND2x1p5_ASAP7_75t_L g750 ( 
.A(n_702),
.B(n_669),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_707),
.B(n_605),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_647),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_721),
.B(n_578),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_714),
.B(n_583),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

BUFx2_ASAP7_75t_L g756 ( 
.A(n_647),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_716),
.B(n_630),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_686),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_695),
.B(n_631),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_647),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_690),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_672),
.B(n_633),
.Y(n_762)
);

NAND3x1_ASAP7_75t_L g763 ( 
.A(n_649),
.B(n_435),
.C(n_423),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_661),
.B(n_417),
.Y(n_764)
);

AND2x4_ASAP7_75t_L g765 ( 
.A(n_664),
.B(n_605),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_664),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_664),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_673),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_687),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_710),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_718),
.B(n_421),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_687),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_693),
.B(n_605),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_712),
.Y(n_774)
);

AND2x4_ASAP7_75t_L g775 ( 
.A(n_715),
.B(n_594),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_689),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_722),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_699),
.B(n_430),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_667),
.B(n_594),
.Y(n_779)
);

AO22x2_ASAP7_75t_L g780 ( 
.A1(n_654),
.A2(n_642),
.B1(n_618),
.B2(n_521),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_715),
.B(n_618),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_715),
.B(n_642),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_682),
.B(n_430),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_689),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_681),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_704),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_665),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_689),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_735),
.A2(n_585),
.B(n_652),
.C(n_660),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_747),
.Y(n_790)
);

NOR2x1p5_ASAP7_75t_L g791 ( 
.A(n_737),
.B(n_670),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_728),
.B(n_720),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_736),
.B(n_720),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_725),
.Y(n_794)
);

O2A1O1Ixp5_ASAP7_75t_L g795 ( 
.A1(n_738),
.A2(n_593),
.B(n_717),
.C(n_703),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_740),
.A2(n_655),
.B1(n_650),
.B2(n_656),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_731),
.B(n_670),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_739),
.B(n_720),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_730),
.Y(n_799)
);

NOR2xp67_ASAP7_75t_L g800 ( 
.A(n_769),
.B(n_696),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_739),
.B(n_713),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_761),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_787),
.A2(n_211),
.B1(n_196),
.B2(n_207),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_756),
.B(n_713),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_773),
.B(n_788),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_763),
.A2(n_709),
.B1(n_676),
.B2(n_657),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_786),
.B(n_211),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_776),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_773),
.B(n_705),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_747),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_723),
.B(n_727),
.Y(n_811)
);

INVx2_ASAP7_75t_SL g812 ( 
.A(n_776),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_723),
.B(n_709),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_744),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_727),
.B(n_673),
.Y(n_815)
);

OAI22xp33_ASAP7_75t_L g816 ( 
.A1(n_750),
.A2(n_762),
.B1(n_743),
.B2(n_779),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_748),
.B(n_211),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_749),
.B(n_211),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_758),
.B(n_708),
.Y(n_819)
);

NAND2x1p5_ASAP7_75t_L g820 ( 
.A(n_774),
.B(n_702),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_732),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_SL g822 ( 
.A1(n_770),
.A2(n_702),
.B1(n_431),
.B2(n_430),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_777),
.B(n_211),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_741),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_733),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_742),
.B(n_703),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_733),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_743),
.B(n_679),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_755),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_734),
.B(n_679),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_778),
.A2(n_464),
.B1(n_698),
.B2(n_674),
.Y(n_831)
);

INVx8_ASAP7_75t_L g832 ( 
.A(n_788),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_788),
.B(n_431),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_779),
.B(n_674),
.Y(n_834)
);

OAI22xp33_ASAP7_75t_L g835 ( 
.A1(n_750),
.A2(n_717),
.B1(n_653),
.B2(n_431),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_746),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_772),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_785),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_757),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_759),
.B(n_627),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_751),
.B(n_674),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_757),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_746),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_751),
.B(n_431),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_765),
.B(n_653),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_754),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_729),
.B(n_698),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_754),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_762),
.B(n_653),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_765),
.B(n_657),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_784),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_745),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_745),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_771),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_783),
.B(n_676),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_726),
.B(n_698),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_724),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_811),
.B(n_767),
.Y(n_858)
);

OR2x2_ASAP7_75t_L g859 ( 
.A(n_836),
.B(n_771),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_827),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_846),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_827),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_857),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_802),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_825),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_825),
.Y(n_866)
);

AND2x4_ASAP7_75t_SL g867 ( 
.A(n_804),
.B(n_752),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_836),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_816),
.B(n_752),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_848),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_816),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_832),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_790),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_852),
.B(n_766),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_843),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_801),
.B(n_819),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_839),
.B(n_780),
.Y(n_878)
);

AND2x2_ASAP7_75t_SL g879 ( 
.A(n_853),
.B(n_752),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_829),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_790),
.B(n_766),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_821),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_842),
.B(n_780),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_811),
.B(n_753),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_794),
.Y(n_885)
);

AND2x2_ASAP7_75t_SL g886 ( 
.A(n_792),
.B(n_760),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_801),
.B(n_764),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_828),
.B(n_760),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_798),
.B(n_760),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_810),
.B(n_768),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_799),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_824),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_814),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_854),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_792),
.B(n_775),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_815),
.B(n_775),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_791),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_789),
.A2(n_782),
.B(n_781),
.Y(n_898)
);

AND2x2_ASAP7_75t_SL g899 ( 
.A(n_841),
.B(n_781),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_820),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_815),
.B(n_838),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_793),
.B(n_782),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_826),
.B(n_698),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_823),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_817),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_871),
.A2(n_789),
.B(n_835),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_L g907 ( 
.A(n_869),
.B(n_807),
.C(n_796),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_863),
.B(n_840),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_905),
.B(n_904),
.C(n_873),
.Y(n_909)
);

CKINVDCx10_ASAP7_75t_R g910 ( 
.A(n_863),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_878),
.A2(n_835),
.B(n_849),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_874),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_874),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_L g914 ( 
.A1(n_904),
.A2(n_834),
.B(n_849),
.Y(n_914)
);

OAI22xp5_ASAP7_75t_L g915 ( 
.A1(n_895),
.A2(n_831),
.B1(n_822),
.B2(n_809),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_873),
.A2(n_795),
.B(n_806),
.C(n_818),
.Y(n_916)
);

AOI21xp33_ASAP7_75t_L g917 ( 
.A1(n_905),
.A2(n_795),
.B(n_813),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_883),
.B(n_830),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_898),
.A2(n_844),
.B(n_845),
.Y(n_919)
);

NOR2x1_ASAP7_75t_R g920 ( 
.A(n_864),
.B(n_808),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_895),
.A2(n_850),
.B(n_805),
.Y(n_921)
);

AO21x1_ASAP7_75t_L g922 ( 
.A1(n_881),
.A2(n_820),
.B(n_855),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_864),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_875),
.Y(n_924)
);

O2A1O1Ixp5_ASAP7_75t_L g925 ( 
.A1(n_900),
.A2(n_833),
.B(n_855),
.C(n_856),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_890),
.B(n_813),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_886),
.B(n_797),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_887),
.A2(n_800),
.B(n_803),
.C(n_812),
.Y(n_928)
);

CKINVDCx10_ASAP7_75t_R g929 ( 
.A(n_875),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_886),
.A2(n_803),
.B(n_847),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_877),
.A2(n_851),
.B(n_209),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_899),
.A2(n_832),
.B(n_437),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_899),
.A2(n_832),
.B(n_437),
.Y(n_933)
);

INVx2_ASAP7_75t_SL g934 ( 
.A(n_867),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_901),
.B(n_885),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_880),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_897),
.B(n_627),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_858),
.B(n_596),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_897),
.B(n_436),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_881),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_903),
.A2(n_620),
.B1(n_479),
.B2(n_436),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_891),
.B(n_194),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_874),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_879),
.A2(n_220),
.B(n_216),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_881),
.Y(n_945)
);

A2O1A1Ixp33_ASAP7_75t_L g946 ( 
.A1(n_900),
.A2(n_177),
.B(n_190),
.C(n_175),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_872),
.B(n_620),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_879),
.A2(n_191),
.B1(n_197),
.B2(n_219),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_884),
.B(n_416),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_891),
.B(n_459),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_884),
.B(n_0),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_894),
.B(n_1),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_900),
.A2(n_210),
.B(n_208),
.C(n_212),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_894),
.B(n_1),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_867),
.A2(n_210),
.B(n_213),
.C(n_215),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_902),
.B(n_2),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_2),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_858),
.B(n_3),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_872),
.B(n_432),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_868),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_872),
.B(n_469),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_896),
.B(n_3),
.Y(n_962)
);

BUFx12f_ASAP7_75t_L g963 ( 
.A(n_924),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_910),
.B(n_896),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_906),
.A2(n_888),
.B(n_866),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_937),
.B(n_889),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_929),
.B(n_872),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_916),
.A2(n_882),
.B(n_880),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_907),
.B(n_865),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_949),
.B(n_872),
.Y(n_970)
);

CKINVDCx10_ASAP7_75t_R g971 ( 
.A(n_923),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_940),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_936),
.Y(n_973)
);

BUFx8_ASAP7_75t_L g974 ( 
.A(n_938),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_928),
.A2(n_882),
.B(n_865),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_944),
.A2(n_859),
.B(n_892),
.Y(n_976)
);

AOI21x1_ASAP7_75t_L g977 ( 
.A1(n_958),
.A2(n_860),
.B(n_862),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_907),
.B(n_861),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_931),
.A2(n_859),
.B(n_892),
.Y(n_979)
);

NAND3xp33_ASAP7_75t_SL g980 ( 
.A(n_922),
.B(n_862),
.C(n_893),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_953),
.A2(n_893),
.B(n_876),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_927),
.A2(n_876),
.B(n_870),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_969),
.B(n_909),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_968),
.A2(n_946),
.B(n_954),
.C(n_952),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_975),
.B(n_921),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_978),
.A2(n_948),
.B1(n_915),
.B2(n_919),
.Y(n_986)
);

AO31x2_ASAP7_75t_L g987 ( 
.A1(n_972),
.A2(n_962),
.A3(n_951),
.B(n_957),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_970),
.A2(n_965),
.B1(n_934),
.B2(n_966),
.Y(n_988)
);

HB1xp67_ASAP7_75t_L g989 ( 
.A(n_977),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_980),
.A2(n_920),
.B(n_911),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_976),
.A2(n_930),
.B1(n_918),
.B2(n_926),
.Y(n_991)
);

AND2x6_ASAP7_75t_L g992 ( 
.A(n_967),
.B(n_962),
.Y(n_992)
);

AO32x1_ASAP7_75t_L g993 ( 
.A1(n_973),
.A2(n_945),
.A3(n_941),
.B1(n_912),
.B2(n_913),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_963),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_979),
.B(n_909),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_964),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_974),
.B(n_925),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_971),
.B(n_950),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_981),
.A2(n_961),
.B(n_939),
.Y(n_999)
);

OR2x2_ASAP7_75t_L g1000 ( 
.A(n_982),
.B(n_935),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_974),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_974),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_972),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_967),
.B(n_908),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_980),
.B(n_956),
.C(n_933),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_968),
.A2(n_925),
.B(n_955),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_R g1007 ( 
.A(n_971),
.B(n_4),
.Y(n_1007)
);

INVx4_ASAP7_75t_L g1008 ( 
.A(n_1001),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_992),
.B(n_914),
.Y(n_1009)
);

AND3x1_ASAP7_75t_SL g1010 ( 
.A(n_997),
.B(n_917),
.C(n_940),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_992),
.B(n_960),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_1007),
.Y(n_1012)
);

BUFx8_ASAP7_75t_L g1013 ( 
.A(n_1002),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_994),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_1003),
.Y(n_1015)
);

NAND2x1_ASAP7_75t_L g1016 ( 
.A(n_1008),
.B(n_992),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_1009),
.A2(n_990),
.B(n_1006),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_1011),
.A2(n_985),
.B(n_989),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_1017),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_SL g1020 ( 
.A(n_1016),
.B(n_996),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_1020),
.A2(n_1018),
.B(n_983),
.Y(n_1021)
);

NAND2x1p5_ASAP7_75t_L g1022 ( 
.A(n_1020),
.B(n_996),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_1022),
.B(n_1014),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1022),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_1023),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1023),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1025),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_1028),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_1027),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1029),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1033),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1031),
.B(n_1025),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1032),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_1034),
.B(n_1013),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_1035),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_1037),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1038),
.B(n_1019),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1040),
.Y(n_1041)
);

AND2x4_ASAP7_75t_SL g1042 ( 
.A(n_1039),
.B(n_1036),
.Y(n_1042)
);

INVx2_ASAP7_75t_SL g1043 ( 
.A(n_1042),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_1041),
.Y(n_1044)
);

AND2x2_ASAP7_75t_L g1045 ( 
.A(n_1043),
.B(n_1012),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1044),
.B(n_1021),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1045),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1046),
.B(n_1015),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_1048),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1047),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_1004),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1051),
.Y(n_1052)
);

XOR2x2_ASAP7_75t_L g1053 ( 
.A(n_1050),
.B(n_1013),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_1049),
.B(n_986),
.Y(n_1054)
);

INVxp67_ASAP7_75t_L g1055 ( 
.A(n_1053),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_1052),
.A2(n_998),
.B(n_995),
.C(n_984),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_1055),
.B(n_1054),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1056),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1058),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1059),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1060),
.B(n_987),
.Y(n_1062)
);

INVx1_ASAP7_75t_SL g1063 ( 
.A(n_1061),
.Y(n_1063)
);

INVxp67_ASAP7_75t_SL g1064 ( 
.A(n_1062),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1063),
.Y(n_1065)
);

OAI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1010),
.B1(n_988),
.B2(n_1000),
.Y(n_1066)
);

OAI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1065),
.A2(n_942),
.B1(n_991),
.B2(n_222),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1066),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_1065),
.B(n_1005),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_1068),
.A2(n_993),
.B(n_999),
.Y(n_1070)
);

AOI221xp5_ASAP7_75t_L g1071 ( 
.A1(n_1069),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1067),
.B(n_6),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_1072),
.B(n_987),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_SL g1074 ( 
.A(n_1071),
.B(n_7),
.C(n_8),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_1073),
.B(n_1070),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1074),
.Y(n_1076)
);

NAND4xp75_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_9),
.C(n_11),
.D(n_12),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_1076),
.B(n_399),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1078),
.Y(n_1079)
);

OAI211xp5_ASAP7_75t_SL g1080 ( 
.A1(n_1077),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_1080)
);

AO22x1_ASAP7_75t_L g1081 ( 
.A1(n_1079),
.A2(n_399),
.B1(n_412),
.B2(n_419),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1080),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_1082),
.B(n_13),
.Y(n_1083)
);

NAND3xp33_ASAP7_75t_SL g1084 ( 
.A(n_1081),
.B(n_13),
.C(n_14),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_1085)
);

AOI222xp33_ASAP7_75t_L g1086 ( 
.A1(n_1083),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.C1(n_19),
.C2(n_20),
.Y(n_1086)
);

OAI211xp5_ASAP7_75t_SL g1087 ( 
.A1(n_1084),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1085),
.B(n_21),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_1087),
.A2(n_1086),
.B1(n_23),
.B2(n_24),
.Y(n_1089)
);

NOR2x1_ASAP7_75t_L g1090 ( 
.A(n_1087),
.B(n_22),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1090),
.Y(n_1091)
);

NAND2xp33_ASAP7_75t_SL g1092 ( 
.A(n_1089),
.B(n_23),
.Y(n_1092)
);

OAI211xp5_ASAP7_75t_L g1093 ( 
.A1(n_1091),
.A2(n_1088),
.B(n_26),
.C(n_27),
.Y(n_1093)
);

AOI211x1_ASAP7_75t_SL g1094 ( 
.A1(n_1092),
.A2(n_25),
.B(n_26),
.C(n_28),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_1094),
.B(n_25),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_1093),
.B(n_28),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_1095),
.B(n_29),
.C(n_30),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1096),
.B(n_29),
.Y(n_1098)
);

AO21x1_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_30),
.B(n_428),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_1098),
.B(n_31),
.C(n_32),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1100),
.B(n_34),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1099),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1102),
.B(n_420),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1101),
.Y(n_1104)
);

OR2x2_ASAP7_75t_L g1105 ( 
.A(n_1102),
.B(n_35),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_1104),
.A2(n_36),
.B(n_38),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1103),
.B(n_420),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_1105),
.Y(n_1108)
);

NOR4xp25_ASAP7_75t_L g1109 ( 
.A(n_1108),
.B(n_40),
.C(n_41),
.D(n_44),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1107),
.A2(n_516),
.B1(n_420),
.B2(n_50),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1109),
.A2(n_1106),
.B(n_932),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1110),
.A2(n_420),
.B1(n_522),
.B2(n_51),
.Y(n_1112)
);

AOI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1112),
.A2(n_45),
.B1(n_47),
.B2(n_52),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1111),
.A2(n_947),
.B(n_959),
.Y(n_1114)
);

OR5x1_ASAP7_75t_L g1115 ( 
.A(n_1113),
.B(n_53),
.C(n_54),
.D(n_55),
.E(n_57),
.Y(n_1115)
);

NAND3xp33_ASAP7_75t_SL g1116 ( 
.A(n_1114),
.B(n_58),
.C(n_59),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_1116),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1115),
.A2(n_63),
.B(n_64),
.Y(n_1118)
);

OAI22x1_ASAP7_75t_L g1119 ( 
.A1(n_1118),
.A2(n_1117),
.B1(n_66),
.B2(n_68),
.Y(n_1119)
);

XNOR2xp5_ASAP7_75t_L g1120 ( 
.A(n_1118),
.B(n_65),
.Y(n_1120)
);

OAI22x1_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_72),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1119),
.Y(n_1123)
);

OAI22x1_ASAP7_75t_L g1124 ( 
.A1(n_1123),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_82),
.Y(n_1125)
);

AO21x2_ASAP7_75t_L g1126 ( 
.A1(n_1123),
.A2(n_77),
.B(n_86),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1123),
.A2(n_87),
.B(n_88),
.Y(n_1127)
);

XNOR2x1_ASAP7_75t_L g1128 ( 
.A(n_1125),
.B(n_89),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_514),
.B1(n_484),
.B2(n_482),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1124),
.Y(n_1130)
);

XNOR2x1_ASAP7_75t_L g1131 ( 
.A(n_1130),
.B(n_1127),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1128),
.A2(n_90),
.B(n_92),
.Y(n_1132)
);

XNOR2x1_ASAP7_75t_L g1133 ( 
.A(n_1129),
.B(n_94),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1131),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1133),
.B(n_95),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1132),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1131),
.B(n_97),
.Y(n_1137)
);

OA21x2_ASAP7_75t_L g1138 ( 
.A1(n_1131),
.A2(n_98),
.B(n_100),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1131),
.B(n_101),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1131),
.A2(n_470),
.B1(n_482),
.B2(n_481),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1131),
.A2(n_470),
.B1(n_482),
.B2(n_481),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1131),
.A2(n_514),
.B1(n_470),
.B2(n_482),
.Y(n_1142)
);

XNOR2xp5_ASAP7_75t_L g1143 ( 
.A(n_1131),
.B(n_103),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1131),
.A2(n_514),
.B1(n_470),
.B2(n_481),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1131),
.A2(n_466),
.B1(n_481),
.B2(n_473),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1134),
.B(n_104),
.Y(n_1146)
);

OAI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1136),
.A2(n_466),
.B1(n_473),
.B2(n_524),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1135),
.Y(n_1148)
);

INVx1_ASAP7_75t_SL g1149 ( 
.A(n_1138),
.Y(n_1149)
);

XNOR2xp5_ASAP7_75t_L g1150 ( 
.A(n_1138),
.B(n_105),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1137),
.B(n_106),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1139),
.A2(n_473),
.B1(n_498),
.B2(n_524),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1143),
.A2(n_473),
.B1(n_498),
.B2(n_524),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1142),
.A2(n_498),
.B1(n_524),
.B2(n_110),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1149),
.A2(n_1144),
.B(n_1145),
.Y(n_1155)
);

AOI322xp5_ASAP7_75t_R g1156 ( 
.A1(n_1148),
.A2(n_107),
.A3(n_108),
.B1(n_111),
.B2(n_112),
.C1(n_113),
.C2(n_114),
.Y(n_1156)
);

XOR2xp5_ASAP7_75t_L g1157 ( 
.A(n_1150),
.B(n_1141),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_1151),
.Y(n_1158)
);

XOR2xp5_ASAP7_75t_L g1159 ( 
.A(n_1154),
.B(n_1140),
.Y(n_1159)
);

AOI222xp33_ASAP7_75t_L g1160 ( 
.A1(n_1153),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.C1(n_122),
.C2(n_124),
.Y(n_1160)
);

AO22x2_ASAP7_75t_L g1161 ( 
.A1(n_1152),
.A2(n_125),
.B1(n_126),
.B2(n_127),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1158),
.A2(n_1146),
.B(n_1147),
.Y(n_1162)
);

A2O1A1O1Ixp25_ASAP7_75t_L g1163 ( 
.A1(n_1155),
.A2(n_128),
.B(n_129),
.C(n_131),
.D(n_132),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1159),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_1164),
.A2(n_1157),
.B1(n_1161),
.B2(n_1156),
.C1(n_1160),
.C2(n_142),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1165),
.B(n_1162),
.Y(n_1166)
);

OR2x6_ASAP7_75t_L g1167 ( 
.A(n_1166),
.B(n_1163),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1167),
.A2(n_135),
.B1(n_137),
.B2(n_140),
.C(n_141),
.Y(n_1168)
);

AOI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1168),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1169),
.A2(n_150),
.B1(n_153),
.B2(n_155),
.Y(n_1170)
);

AOI211xp5_ASAP7_75t_L g1171 ( 
.A1(n_1170),
.A2(n_943),
.B(n_157),
.C(n_158),
.Y(n_1171)
);

AOI211xp5_ASAP7_75t_L g1172 ( 
.A1(n_1171),
.A2(n_156),
.B(n_159),
.C(n_160),
.Y(n_1172)
);


endmodule