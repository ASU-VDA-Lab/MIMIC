module fake_jpeg_12004_n_233 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_233);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_233;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_1),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_0),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_55),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_29),
.Y(n_74)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_18),
.B(n_1),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_63),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_26),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_57),
.Y(n_79)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_59),
.Y(n_95)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_62),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_35),
.B1(n_45),
.B2(n_57),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_64),
.A2(n_69),
.B1(n_83),
.B2(n_52),
.Y(n_102)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_35),
.B1(n_25),
.B2(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_32),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_73),
.B(n_74),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_25),
.B1(n_36),
.B2(n_34),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_65),
.B1(n_33),
.B2(n_18),
.Y(n_111)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_22),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_92),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_41),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_106),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_19),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_119),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_70),
.B(n_42),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_104),
.B(n_118),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_110),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_80),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_80),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_69),
.A2(n_40),
.B1(n_20),
.B2(n_28),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g117 ( 
.A1(n_83),
.A2(n_22),
.B1(n_19),
.B2(n_30),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_70),
.B(n_22),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_67),
.B(n_19),
.C(n_30),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_21),
.B1(n_30),
.B2(n_4),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_90),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_75),
.B1(n_90),
.B2(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_72),
.Y(n_134)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_79),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_126),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_118),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_108),
.C(n_66),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_98),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_147),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_114),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_77),
.B1(n_93),
.B2(n_76),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_76),
.B1(n_71),
.B2(n_68),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_95),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_71),
.B1(n_59),
.B2(n_81),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_149),
.A2(n_116),
.B1(n_115),
.B2(n_91),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_119),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_100),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_131),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_154),
.C(n_170),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_118),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_104),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_155),
.B(n_156),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_104),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_148),
.B(n_113),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_167),
.Y(n_183)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_159),
.B(n_166),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_163),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_161),
.A2(n_123),
.B1(n_144),
.B2(n_91),
.Y(n_188)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_141),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_165),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_110),
.B1(n_101),
.B2(n_126),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_148),
.B(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_169),
.C(n_143),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_108),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_182),
.Y(n_196)
);

AOI322xp5_ASAP7_75t_SL g173 ( 
.A1(n_171),
.A2(n_139),
.A3(n_129),
.B1(n_138),
.B2(n_130),
.C1(n_6),
.C2(n_7),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_178),
.A3(n_184),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_192)
);

AOI221xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_135),
.B1(n_137),
.B2(n_132),
.C(n_140),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_SL g178 ( 
.A(n_155),
.B(n_160),
.C(n_153),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_132),
.B(n_105),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_179),
.A2(n_136),
.B(n_21),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_152),
.Y(n_182)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_2),
.C(n_3),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_144),
.C(n_127),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_170),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_163),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_161),
.B1(n_166),
.B2(n_165),
.Y(n_189)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_154),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_193),
.C(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_9),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_175),
.C(n_21),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_181),
.A3(n_187),
.B1(n_182),
.B2(n_186),
.C1(n_178),
.C2(n_188),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_187),
.A3(n_174),
.B1(n_185),
.B2(n_177),
.C1(n_175),
.C2(n_21),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_183),
.B(n_157),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_158),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_21),
.C(n_9),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_136),
.B(n_127),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_198),
.A2(n_201),
.B(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_202),
.A2(n_208),
.B(n_201),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_5),
.B(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_10),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_214),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_199),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_204),
.B(n_199),
.Y(n_216)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_216),
.Y(n_222)
);

NAND4xp25_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_209),
.C(n_191),
.D(n_197),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_193),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_10),
.B(n_11),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_203),
.C(n_195),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_203),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_224),
.C(n_226),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_219),
.B(n_211),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_10),
.C(n_11),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_220),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_224),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g230 ( 
.A1(n_229),
.A2(n_222),
.B(n_221),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_228),
.C(n_13),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_232),
.B(n_231),
.Y(n_233)
);


endmodule