module fake_netlist_5_1466_n_1699 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1699);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1699;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_86),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_52),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_50),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_8),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_56),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_16),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_106),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_34),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_28),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_46),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_35),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_145),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_61),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_12),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_26),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_41),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_65),
.Y(n_179)
);

BUFx10_ASAP7_75t_L g180 ( 
.A(n_16),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_125),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_34),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_36),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_73),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_4),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_31),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_5),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_49),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_123),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_19),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_38),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_109),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_60),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_8),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_51),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_15),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_144),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_53),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_26),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_66),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_46),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_149),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_95),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_9),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_118),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_31),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_49),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_57),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_21),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_75),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_83),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_39),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_91),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_7),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_41),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_62),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_38),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_30),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_80),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_32),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_45),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_108),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_71),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_147),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_98),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_93),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_112),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_58),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_67),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_7),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_151),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_146),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_39),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_94),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_122),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_100),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_72),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_82),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_102),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_32),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_97),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_115),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_59),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_107),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_134),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_4),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_148),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_48),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_63),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_84),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_79),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_42),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_116),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_18),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_88),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_2),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_47),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_23),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_85),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_126),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_22),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_138),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_20),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_14),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_47),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_10),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_129),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_23),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_14),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_150),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_76),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_99),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_121),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_15),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_165),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_204),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_215),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_245),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_165),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_177),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_184),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_154),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_184),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_267),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_210),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_234),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_160),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_157),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_158),
.Y(n_324)
);

INVxp33_ASAP7_75t_SL g325 ( 
.A(n_155),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_162),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_176),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_176),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_170),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_182),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_152),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_245),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_178),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_182),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_189),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_189),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_191),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_191),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_194),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_171),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_200),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_172),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_200),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g347 ( 
.A(n_156),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_258),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_261),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_194),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_202),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_173),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_202),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_222),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_222),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_175),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_228),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_228),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_239),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_179),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_261),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_239),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_241),
.Y(n_363)
);

INVxp67_ASAP7_75t_SL g364 ( 
.A(n_301),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_241),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_252),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_252),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_288),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_227),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_288),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_181),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_260),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_292),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_292),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_185),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_306),
.B(n_161),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_307),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_304),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_287),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_318),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_190),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_318),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_305),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_369),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_311),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_369),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_348),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_322),
.B(n_192),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_301),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_328),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_334),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g400 ( 
.A(n_336),
.B(n_260),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_364),
.B(n_193),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_315),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_344),
.A2(n_283),
.B1(n_273),
.B2(n_296),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_303),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_346),
.A2(n_242),
.B1(n_275),
.B2(n_169),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_328),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_317),
.A2(n_300),
.B1(n_302),
.B2(n_167),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_329),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_329),
.A2(n_187),
.B(n_159),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_372),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_361),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_323),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_330),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_331),
.B(n_199),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_303),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_324),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_308),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_308),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_331),
.B(n_201),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_309),
.Y(n_420)
);

AND2x6_ASAP7_75t_L g421 ( 
.A(n_333),
.B(n_227),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_333),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_337),
.B(n_207),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_337),
.B(n_159),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_338),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_309),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_338),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_339),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g429 ( 
.A1(n_310),
.A2(n_300),
.B(n_166),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_310),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_312),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_312),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_314),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_339),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_314),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_316),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_316),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_341),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_342),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_319),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_319),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_384),
.B(n_327),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_384),
.B(n_332),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_429),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_379),
.B(n_325),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_401),
.B(n_347),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_411),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_385),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_385),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_429),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_401),
.B(n_343),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_411),
.B(n_320),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_399),
.Y(n_466)
);

BUFx6f_ASAP7_75t_SL g467 ( 
.A(n_416),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_394),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_416),
.B(n_152),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_380),
.B(n_345),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_385),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_404),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_400),
.A2(n_231),
.B1(n_295),
.B2(n_293),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_397),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_402),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_404),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_380),
.B(n_352),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_414),
.B(n_356),
.Y(n_482)
);

INVx4_ASAP7_75t_L g483 ( 
.A(n_385),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_414),
.B(n_360),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

NAND2xp33_ASAP7_75t_SL g486 ( 
.A(n_396),
.B(n_410),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_397),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_419),
.B(n_371),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_398),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_419),
.B(n_375),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_395),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_395),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_R g497 ( 
.A(n_391),
.B(n_211),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_389),
.B(n_412),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_406),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

BUFx3_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_402),
.B(n_163),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_408),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_422),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_402),
.B(n_163),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_422),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_377),
.Y(n_512)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_342),
.Y(n_513)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_410),
.B(n_350),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_394),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_395),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_440),
.B(n_425),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_377),
.B(n_153),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_393),
.B(n_208),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_418),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_423),
.B(n_400),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_381),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_394),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_423),
.A2(n_250),
.B1(n_203),
.B2(n_196),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_425),
.Y(n_525)
);

INVx6_ASAP7_75t_L g526 ( 
.A(n_394),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_418),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_427),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_427),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_407),
.B(n_208),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_440),
.B(n_320),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_428),
.B(n_195),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_407),
.B(n_297),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_428),
.B(n_226),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_434),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_434),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_405),
.A2(n_186),
.B1(n_255),
.B2(n_244),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_405),
.B(n_297),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_424),
.B(n_297),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_424),
.B(n_213),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_424),
.B(n_214),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_437),
.B(n_249),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_391),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_439),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_439),
.B(n_321),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_441),
.Y(n_547)
);

AOI22x1_ASAP7_75t_L g548 ( 
.A1(n_424),
.A2(n_238),
.B1(n_236),
.B2(n_221),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_418),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_387),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_409),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_424),
.A2(n_236),
.B1(n_238),
.B2(n_188),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_441),
.B(n_168),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_409),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_442),
.B(n_321),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_L g556 ( 
.A(n_421),
.B(n_227),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_403),
.B(n_216),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_442),
.B(n_197),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_409),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_376),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_387),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_421),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_381),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_381),
.B(n_383),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_376),
.B(n_198),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_378),
.A2(n_243),
.B1(n_233),
.B2(n_232),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_378),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_417),
.A2(n_188),
.B1(n_221),
.B2(n_187),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_417),
.A2(n_209),
.B1(n_298),
.B2(n_282),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_382),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_403),
.B(n_223),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_382),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_418),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_431),
.Y(n_574)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_421),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_381),
.B(n_224),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_386),
.B(n_166),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_417),
.B(n_205),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_431),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_383),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_417),
.B(n_350),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_431),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_431),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_417),
.A2(n_229),
.B1(n_218),
.B2(n_225),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_432),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_420),
.B(n_351),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_432),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_432),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_420),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_451),
.B(n_420),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_462),
.B(n_420),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g594 ( 
.A(n_491),
.B(n_351),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_512),
.B(n_206),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_462),
.B(n_420),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_426),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_521),
.B(n_227),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_518),
.B(n_284),
.C(n_285),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_445),
.B(n_426),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_560),
.Y(n_601)
);

AOI221xp5_ASAP7_75t_L g602 ( 
.A1(n_538),
.A2(n_259),
.B1(n_212),
.B2(n_217),
.C(n_290),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_469),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_550),
.B(n_174),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_482),
.B(n_227),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_472),
.A2(n_263),
.B1(n_235),
.B2(n_247),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_461),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_484),
.B(n_254),
.Y(n_608)
);

BUFx2_ASAP7_75t_L g609 ( 
.A(n_550),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_496),
.A2(n_388),
.B(n_390),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_502),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_488),
.B(n_254),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_463),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_463),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_446),
.B(n_426),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_458),
.B(n_426),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_466),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_481),
.B(n_220),
.Y(n_618)
);

INVxp33_ASAP7_75t_L g619 ( 
.A(n_450),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_493),
.B(n_254),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_466),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_551),
.B(n_254),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_497),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_452),
.B(n_426),
.Y(n_625)
);

INVx4_ASAP7_75t_L g626 ( 
.A(n_526),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_515),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_513),
.B(n_291),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_452),
.B(n_430),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_468),
.B(n_430),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_517),
.B(n_180),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_513),
.B(n_353),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_551),
.B(n_248),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g634 ( 
.A(n_498),
.B(n_251),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_523),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_523),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_551),
.B(n_254),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_479),
.B(n_353),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_526),
.Y(n_639)
);

INVx2_ASAP7_75t_SL g640 ( 
.A(n_514),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_473),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_526),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_514),
.B(n_174),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_551),
.B(n_209),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_517),
.B(n_183),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_471),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_473),
.B(n_430),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_470),
.A2(n_250),
.B1(n_298),
.B2(n_196),
.Y(n_648)
);

BUFx5_ASAP7_75t_L g649 ( 
.A(n_447),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_486),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_544),
.B(n_354),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_478),
.B(n_430),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_531),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_471),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_475),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_557),
.B(n_183),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_571),
.B(n_203),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_560),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_447),
.A2(n_280),
.B1(n_219),
.B2(n_230),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_487),
.B(n_430),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_487),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_475),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_489),
.B(n_490),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_489),
.B(n_430),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_490),
.B(n_430),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_495),
.Y(n_667)
);

NOR3xp33_ASAP7_75t_L g668 ( 
.A(n_530),
.B(n_280),
.C(n_230),
.Y(n_668)
);

AOI221xp5_ASAP7_75t_L g669 ( 
.A1(n_533),
.A2(n_359),
.B1(n_354),
.B2(n_374),
.C(n_373),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_495),
.B(n_430),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_531),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_500),
.B(n_436),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_500),
.B(n_436),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_449),
.B(n_253),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_501),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_501),
.B(n_436),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_449),
.B(n_256),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_464),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_567),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_477),
.B(n_219),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_453),
.B(n_262),
.Y(n_681)
);

BUFx10_ASAP7_75t_L g682 ( 
.A(n_544),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_506),
.B(n_436),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_453),
.B(n_265),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_457),
.A2(n_460),
.B(n_459),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_506),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_508),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_457),
.B(n_266),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_467),
.B(n_413),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_477),
.B(n_237),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_508),
.B(n_436),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_561),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_L g693 ( 
.A(n_459),
.B(n_268),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_511),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_511),
.B(n_436),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_460),
.B(n_270),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_525),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_525),
.B(n_436),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_476),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_503),
.B(n_237),
.C(n_240),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_575),
.B(n_271),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_528),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_464),
.B(n_355),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_546),
.Y(n_704)
);

NOR3xp33_ASAP7_75t_L g705 ( 
.A(n_509),
.B(n_282),
.C(n_246),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_528),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_546),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_553),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_529),
.B(n_436),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_529),
.B(n_246),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_535),
.B(n_257),
.Y(n_711)
);

CKINVDCx20_ASAP7_75t_R g712 ( 
.A(n_561),
.Y(n_712)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_558),
.B(n_274),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_535),
.B(n_257),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_536),
.B(n_264),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_566),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_536),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_540),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_578),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_540),
.B(n_545),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_575),
.B(n_276),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_470),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_565),
.B(n_277),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_545),
.B(n_264),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_575),
.B(n_278),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_524),
.A2(n_272),
.B1(n_269),
.B2(n_367),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_547),
.B(n_269),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_272),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_555),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_524),
.A2(n_368),
.B1(n_355),
.B2(n_357),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_582),
.B(n_383),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_590),
.B(n_286),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_582),
.B(n_383),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_590),
.B(n_289),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_587),
.B(n_388),
.Y(n_735)
);

BUFx5_ASAP7_75t_L g736 ( 
.A(n_559),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_470),
.A2(n_294),
.B1(n_443),
.B2(n_438),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_587),
.B(n_388),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_554),
.B(n_432),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_467),
.A2(n_421),
.B1(n_443),
.B2(n_438),
.Y(n_740)
);

INVx3_ASAP7_75t_L g741 ( 
.A(n_581),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_555),
.Y(n_742)
);

INVx4_ASAP7_75t_L g743 ( 
.A(n_494),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_505),
.B(n_388),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_SL g745 ( 
.A(n_467),
.B(n_413),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_567),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_505),
.B(n_390),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_470),
.A2(n_421),
.B1(n_443),
.B2(n_438),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_570),
.Y(n_749)
);

OAI22xp33_ASAP7_75t_L g750 ( 
.A1(n_470),
.A2(n_585),
.B1(n_532),
.B2(n_534),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_570),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_543),
.B(n_519),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_572),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_581),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_537),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_708),
.B(n_752),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_649),
.B(n_572),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_752),
.B(n_585),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_601),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_624),
.Y(n_760)
);

INVx6_ASAP7_75t_L g761 ( 
.A(n_682),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_712),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_649),
.B(n_576),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_659),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_594),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_679),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_649),
.B(n_576),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_680),
.A2(n_578),
.B1(n_548),
.B2(n_569),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_618),
.A2(n_541),
.B1(n_542),
.B2(n_577),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_639),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_632),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_654),
.B(n_539),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_704),
.B(n_578),
.Y(n_773)
);

OAI22xp5_ASAP7_75t_SL g774 ( 
.A1(n_755),
.A2(n_537),
.B1(n_552),
.B2(n_370),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_635),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_649),
.B(n_554),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_SL g777 ( 
.A1(n_619),
.A2(n_367),
.B1(n_357),
.B2(n_358),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_649),
.B(n_505),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_707),
.B(n_578),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_749),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_749),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_649),
.B(n_559),
.Y(n_782)
);

AND2x6_ASAP7_75t_SL g783 ( 
.A(n_680),
.B(n_358),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_678),
.B(n_494),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_682),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_685),
.B(n_448),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_720),
.B(n_448),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_720),
.B(n_448),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_740),
.B(n_455),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_753),
.Y(n_790)
);

NOR2x1p5_ASAP7_75t_L g791 ( 
.A(n_599),
.B(n_359),
.Y(n_791)
);

INVx8_ASAP7_75t_L g792 ( 
.A(n_604),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_618),
.A2(n_578),
.B1(n_516),
.B2(n_494),
.Y(n_793)
);

INVx4_ASAP7_75t_L g794 ( 
.A(n_635),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_753),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_746),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_591),
.B(n_455),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_660),
.B(n_455),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_729),
.B(n_494),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_741),
.Y(n_800)
);

O2A1O1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_690),
.A2(n_568),
.B(n_589),
.C(n_586),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_660),
.A2(n_548),
.B1(n_362),
.B2(n_365),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_742),
.B(n_494),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_750),
.A2(n_516),
.B1(n_456),
.B2(n_465),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_638),
.B(n_362),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_639),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_623),
.A2(n_564),
.B(n_474),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_741),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_609),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_627),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_736),
.B(n_456),
.Y(n_811)
);

INVx5_ASAP7_75t_L g812 ( 
.A(n_626),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_754),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_751),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_690),
.B(n_456),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_638),
.B(n_703),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_736),
.B(n_664),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_703),
.B(n_516),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_754),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_692),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_627),
.B(n_363),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_641),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_607),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_736),
.B(n_465),
.Y(n_824)
);

NOR3x1_ASAP7_75t_L g825 ( 
.A(n_640),
.B(n_368),
.C(n_374),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_642),
.Y(n_826)
);

HB1xp67_ASAP7_75t_SL g827 ( 
.A(n_671),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_651),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_652),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_628),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_713),
.B(n_516),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_657),
.A2(n_516),
.B1(n_588),
.B2(n_586),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_631),
.B(n_628),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_736),
.B(n_465),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_604),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_613),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_614),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_604),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_595),
.B(n_180),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_716),
.B(n_562),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_736),
.B(n_485),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_617),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_650),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_736),
.B(n_485),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_606),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_662),
.B(n_363),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_600),
.B(n_485),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_SL g848 ( 
.A1(n_595),
.A2(n_365),
.B1(n_366),
.B2(n_370),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_667),
.B(n_366),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_642),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_723),
.B(n_562),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_675),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_710),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_643),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_657),
.B(n_562),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_622),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_615),
.B(n_589),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_643),
.B(n_454),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_645),
.B(n_454),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_658),
.B(n_562),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_658),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_689),
.B(n_562),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_686),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_711),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_592),
.A2(n_522),
.B1(n_563),
.B2(n_483),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_SL g866 ( 
.A1(n_726),
.A2(n_373),
.B1(n_180),
.B2(n_3),
.Y(n_866)
);

AOI21x1_ASAP7_75t_L g867 ( 
.A1(n_739),
.A2(n_588),
.B(n_584),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_616),
.B(n_584),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_602),
.B(n_556),
.C(n_435),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_687),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_722),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_694),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_697),
.B(n_583),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_603),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_745),
.B(n_562),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_611),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_702),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_706),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_717),
.B(n_522),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_645),
.B(n_454),
.Y(n_880)
);

AND2x6_ASAP7_75t_L g881 ( 
.A(n_620),
.B(n_480),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_718),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_636),
.Y(n_883)
);

INVx8_ASAP7_75t_L g884 ( 
.A(n_719),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_630),
.Y(n_885)
);

AND2x6_ASAP7_75t_L g886 ( 
.A(n_748),
.B(n_583),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_647),
.Y(n_887)
);

BUFx4f_ASAP7_75t_L g888 ( 
.A(n_656),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_714),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_731),
.B(n_580),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_653),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_SL g892 ( 
.A(n_669),
.B(n_0),
.C(n_1),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_646),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_655),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_732),
.B(n_483),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_634),
.B(n_563),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_733),
.B(n_580),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_735),
.B(n_574),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_715),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_663),
.Y(n_900)
);

BUFx4f_ASAP7_75t_L g901 ( 
.A(n_699),
.Y(n_901)
);

OR2x2_ASAP7_75t_SL g902 ( 
.A(n_668),
.B(n_728),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_661),
.Y(n_903)
);

OR2x2_ASAP7_75t_SL g904 ( 
.A(n_700),
.B(n_433),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_732),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_626),
.B(n_421),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_598),
.A2(n_574),
.B1(n_573),
.B2(n_549),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_665),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_666),
.Y(n_909)
);

CKINVDCx11_ASAP7_75t_R g910 ( 
.A(n_648),
.Y(n_910)
);

INVx5_ASAP7_75t_L g911 ( 
.A(n_743),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_743),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_670),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_738),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_734),
.A2(n_573),
.B1(n_549),
.B2(n_527),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_724),
.B(n_527),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_724),
.B(n_520),
.Y(n_917)
);

NAND2x1p5_ASAP7_75t_L g918 ( 
.A(n_739),
.B(n_480),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_727),
.B(n_520),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_593),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_727),
.B(n_510),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_734),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_SL g923 ( 
.A1(n_726),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_674),
.B(n_5),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_625),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_672),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_673),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_605),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_705),
.B(n_444),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_676),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_SL g931 ( 
.A(n_737),
.B(n_421),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_596),
.B(n_510),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_597),
.B(n_507),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_744),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_623),
.B(n_507),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_674),
.B(n_499),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_758),
.A2(n_598),
.B(n_681),
.C(n_677),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_812),
.A2(n_693),
.B(n_644),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_854),
.B(n_677),
.Y(n_939)
);

OAI221xp5_ASAP7_75t_L g940 ( 
.A1(n_830),
.A2(n_730),
.B1(n_684),
.B2(n_681),
.C(n_688),
.Y(n_940)
);

BUFx12f_ASAP7_75t_L g941 ( 
.A(n_762),
.Y(n_941)
);

OAI22xp5_ASAP7_75t_L g942 ( 
.A1(n_861),
.A2(n_688),
.B1(n_684),
.B2(n_696),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_816),
.B(n_696),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_816),
.B(n_701),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_775),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_833),
.B(n_605),
.Y(n_946)
);

BUFx12f_ASAP7_75t_L g947 ( 
.A(n_761),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_827),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_809),
.Y(n_949)
);

NAND3xp33_ASAP7_75t_L g950 ( 
.A(n_839),
.B(n_730),
.C(n_633),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_817),
.A2(n_637),
.B1(n_725),
.B2(n_721),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_759),
.Y(n_952)
);

BUFx6f_ASAP7_75t_L g953 ( 
.A(n_806),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_905),
.B(n_701),
.Y(n_954)
);

O2A1O1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_924),
.A2(n_612),
.B(n_608),
.C(n_621),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_853),
.B(n_608),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_SL g957 ( 
.A(n_923),
.B(n_621),
.C(n_612),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_756),
.A2(n_637),
.B(n_698),
.C(n_709),
.Y(n_958)
);

OR2x6_ASAP7_75t_SL g959 ( 
.A(n_760),
.B(n_845),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_817),
.A2(n_725),
.B1(n_721),
.B2(n_629),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_775),
.B(n_812),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_812),
.A2(n_911),
.B(n_776),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_771),
.B(n_765),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_792),
.B(n_695),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_859),
.A2(n_747),
.B1(n_691),
.B2(n_683),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_764),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_864),
.B(n_610),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_820),
.B(n_9),
.C(n_10),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_843),
.B(n_11),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_805),
.B(n_444),
.Y(n_970)
);

INVx1_ASAP7_75t_SL g971 ( 
.A(n_761),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_889),
.B(n_504),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_810),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_769),
.A2(n_492),
.B(n_444),
.C(n_443),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_766),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_911),
.A2(n_390),
.B(n_438),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_899),
.B(n_444),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_780),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_858),
.B(n_435),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_880),
.B(n_435),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_SL g981 ( 
.A(n_785),
.B(n_433),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_757),
.A2(n_435),
.B1(n_433),
.B2(n_390),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_802),
.A2(n_787),
.B(n_788),
.C(n_916),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_775),
.B(n_143),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_911),
.A2(n_90),
.B(n_136),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_776),
.A2(n_87),
.B(n_130),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_781),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_778),
.A2(n_77),
.B(n_127),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_796),
.Y(n_989)
);

CKINVDCx16_ASAP7_75t_R g990 ( 
.A(n_871),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_914),
.B(n_421),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_783),
.B(n_11),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_768),
.A2(n_895),
.B(n_877),
.C(n_882),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_814),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_810),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_821),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_757),
.A2(n_124),
.B1(n_114),
.B2(n_104),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_778),
.A2(n_74),
.B(n_70),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_790),
.B(n_68),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_826),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_914),
.B(n_421),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_782),
.A2(n_64),
.B(n_54),
.Y(n_1002)
);

INVx3_ASAP7_75t_L g1003 ( 
.A(n_826),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_774),
.B(n_13),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_795),
.B(n_17),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_821),
.B(n_421),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_782),
.A2(n_19),
.B(n_20),
.Y(n_1007)
);

CKINVDCx16_ASAP7_75t_R g1008 ( 
.A(n_838),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_922),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_826),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_773),
.B(n_779),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_805),
.B(n_822),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_763),
.A2(n_24),
.B(n_25),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_761),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_829),
.B(n_27),
.Y(n_1015)
);

INVx1_ASAP7_75t_SL g1016 ( 
.A(n_828),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_852),
.B(n_28),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_863),
.A2(n_872),
.B(n_878),
.C(n_801),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_846),
.B(n_29),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_773),
.B(n_29),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_823),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_835),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_836),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_802),
.A2(n_33),
.B(n_35),
.C(n_36),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_770),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_846),
.B(n_849),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_873),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_763),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_1028)
);

OAI21xp33_ASAP7_75t_L g1029 ( 
.A1(n_870),
.A2(n_40),
.B(n_42),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_849),
.B(n_50),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_767),
.A2(n_43),
.B1(n_44),
.B2(n_798),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_787),
.A2(n_43),
.B(n_44),
.C(n_788),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_837),
.Y(n_1033)
);

O2A1O1Ixp5_ASAP7_75t_SL g1034 ( 
.A1(n_936),
.A2(n_896),
.B(n_831),
.C(n_772),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_873),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_806),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_916),
.A2(n_921),
.B(n_919),
.C(n_917),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_885),
.B(n_887),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_SL g1039 ( 
.A(n_779),
.B(n_874),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_917),
.A2(n_921),
.B(n_919),
.C(n_892),
.Y(n_1040)
);

BUFx6f_ASAP7_75t_L g1041 ( 
.A(n_806),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_767),
.A2(n_824),
.B(n_841),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_792),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_874),
.B(n_876),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_874),
.B(n_876),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_884),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_792),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_798),
.A2(n_819),
.B1(n_793),
.B2(n_770),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_811),
.A2(n_834),
.B(n_824),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_804),
.A2(n_928),
.B1(n_922),
.B2(n_794),
.Y(n_1050)
);

BUFx4f_ASAP7_75t_L g1051 ( 
.A(n_884),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_884),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_891),
.B(n_903),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_908),
.B(n_909),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_800),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_876),
.B(n_883),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_842),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_R g1058 ( 
.A(n_910),
.B(n_850),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_794),
.A2(n_813),
.B1(n_808),
.B2(n_786),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_786),
.A2(n_888),
.B1(n_901),
.B2(n_927),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_913),
.B(n_926),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_811),
.A2(n_844),
.B(n_841),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_930),
.B(n_925),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_920),
.A2(n_934),
.B(n_869),
.C(n_888),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_815),
.A2(n_883),
.B1(n_818),
.B2(n_866),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_834),
.A2(n_844),
.B(n_912),
.Y(n_1066)
);

NOR2xp67_ASAP7_75t_SL g1067 ( 
.A(n_912),
.B(n_883),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_847),
.A2(n_933),
.B(n_857),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_SL g1069 ( 
.A(n_901),
.B(n_879),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_815),
.B(n_920),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_856),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_815),
.B(n_797),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_850),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_879),
.B(n_848),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_929),
.B(n_875),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_847),
.A2(n_933),
.B(n_857),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_815),
.B(n_797),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_929),
.B(n_862),
.Y(n_1078)
);

INVx3_ASAP7_75t_L g1079 ( 
.A(n_881),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1066),
.A2(n_867),
.B(n_807),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_989),
.Y(n_1081)
);

INVx3_ASAP7_75t_SL g1082 ( 
.A(n_1043),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1068),
.A2(n_868),
.B(n_898),
.Y(n_1083)
);

OR2x2_ASAP7_75t_L g1084 ( 
.A(n_949),
.B(n_902),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_957),
.A2(n_897),
.B1(n_898),
.B2(n_890),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1038),
.B(n_791),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_994),
.Y(n_1087)
);

NAND2xp33_ASAP7_75t_L g1088 ( 
.A(n_957),
.B(n_886),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1053),
.B(n_868),
.Y(n_1089)
);

OA21x2_ASAP7_75t_L g1090 ( 
.A1(n_993),
.A2(n_1062),
.B(n_1049),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_1026),
.B(n_825),
.Y(n_1091)
);

AOI221x1_ASAP7_75t_L g1092 ( 
.A1(n_942),
.A2(n_807),
.B1(n_932),
.B2(n_897),
.C(n_890),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_950),
.A2(n_840),
.B(n_799),
.C(n_803),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1027),
.B(n_900),
.Y(n_1094)
);

OAI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1042),
.A2(n_918),
.B(n_935),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_937),
.A2(n_983),
.B(n_1037),
.Y(n_1096)
);

OR2x2_ASAP7_75t_L g1097 ( 
.A(n_1012),
.B(n_893),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_938),
.A2(n_918),
.B(n_907),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_1035),
.B(n_894),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_1067),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_981),
.B(n_777),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1054),
.B(n_886),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_937),
.A2(n_983),
.B(n_1037),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_L g1104 ( 
.A1(n_962),
.A2(n_915),
.B(n_832),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1040),
.A2(n_886),
.B(n_789),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1061),
.B(n_886),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_1051),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_970),
.B(n_784),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1064),
.A2(n_855),
.B(n_860),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_960),
.A2(n_851),
.B(n_906),
.Y(n_1110)
);

NAND2x1p5_ASAP7_75t_L g1111 ( 
.A(n_953),
.B(n_865),
.Y(n_1111)
);

NOR2xp67_ASAP7_75t_SL g1112 ( 
.A(n_947),
.B(n_906),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1063),
.B(n_881),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1004),
.A2(n_931),
.B(n_904),
.C(n_881),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1040),
.A2(n_940),
.B(n_1077),
.Y(n_1115)
);

NOR2x1_ASAP7_75t_L g1116 ( 
.A(n_1014),
.B(n_881),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_980),
.A2(n_789),
.B(n_979),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_1072),
.A2(n_789),
.B(n_955),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1011),
.B(n_789),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_941),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_965),
.A2(n_955),
.B(n_967),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1070),
.A2(n_1059),
.B(n_982),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_939),
.A2(n_1004),
.B(n_946),
.C(n_1018),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1034),
.A2(n_1048),
.B(n_976),
.Y(n_1124)
);

AOI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1050),
.A2(n_1060),
.B(n_943),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_944),
.A2(n_958),
.B(n_1078),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_958),
.A2(n_1075),
.B(n_973),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_974),
.A2(n_1031),
.A3(n_997),
.B(n_1028),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_963),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_948),
.B(n_1065),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1055),
.Y(n_1131)
);

O2A1O1Ixp5_ASAP7_75t_L g1132 ( 
.A1(n_954),
.A2(n_999),
.B(n_1045),
.C(n_1044),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_996),
.B(n_969),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_952),
.B(n_966),
.Y(n_1134)
);

BUFx12f_ASAP7_75t_L g1135 ( 
.A(n_1047),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_971),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_975),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_L g1138 ( 
.A1(n_1056),
.A2(n_1015),
.B(n_1017),
.C(n_1005),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_969),
.B(n_1055),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1046),
.Y(n_1140)
);

AO21x2_ASAP7_75t_L g1141 ( 
.A1(n_956),
.A2(n_1002),
.B(n_998),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1074),
.B(n_1039),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_1022),
.B(n_1016),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_984),
.A2(n_1024),
.B(n_1069),
.C(n_1030),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1009),
.A2(n_1024),
.B1(n_1019),
.B2(n_972),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1052),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_978),
.Y(n_1147)
);

AO32x2_ASAP7_75t_L g1148 ( 
.A1(n_1032),
.A2(n_945),
.A3(n_1029),
.B1(n_968),
.B2(n_1013),
.Y(n_1148)
);

OA21x2_ASAP7_75t_L g1149 ( 
.A1(n_988),
.A2(n_1007),
.B(n_986),
.Y(n_1149)
);

NAND3xp33_ASAP7_75t_SL g1150 ( 
.A(n_992),
.B(n_1058),
.C(n_968),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1032),
.A2(n_973),
.B1(n_995),
.B2(n_987),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1020),
.A2(n_992),
.B1(n_1071),
.B2(n_1033),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_1079),
.A2(n_995),
.B(n_1001),
.Y(n_1153)
);

NAND2x1p5_ASAP7_75t_L g1154 ( 
.A(n_953),
.B(n_1041),
.Y(n_1154)
);

NOR2xp67_ASAP7_75t_L g1155 ( 
.A(n_945),
.B(n_1021),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_961),
.A2(n_977),
.B(n_991),
.Y(n_1156)
);

AOI211x1_ASAP7_75t_L g1157 ( 
.A1(n_1057),
.A2(n_1006),
.B(n_985),
.C(n_1025),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_959),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_964),
.A2(n_1025),
.B(n_1073),
.Y(n_1159)
);

OA21x2_ASAP7_75t_L g1160 ( 
.A1(n_1023),
.A2(n_964),
.B(n_1073),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_964),
.A2(n_1010),
.B(n_1000),
.Y(n_1161)
);

NOR2x1_ASAP7_75t_SL g1162 ( 
.A(n_953),
.B(n_1041),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1000),
.A2(n_1010),
.B(n_1003),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1008),
.B(n_1058),
.Y(n_1164)
);

NAND2x1p5_ASAP7_75t_L g1165 ( 
.A(n_953),
.B(n_1036),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_1036),
.Y(n_1166)
);

AO32x2_ASAP7_75t_L g1167 ( 
.A1(n_1051),
.A2(n_1036),
.A3(n_1041),
.B1(n_1003),
.B2(n_990),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1036),
.B(n_1041),
.Y(n_1168)
);

O2A1O1Ixp5_ASAP7_75t_SL g1169 ( 
.A1(n_942),
.A2(n_598),
.B(n_758),
.C(n_608),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1027),
.B(n_1035),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1027),
.B(n_1035),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_957),
.A2(n_861),
.B1(n_660),
.B2(n_1065),
.Y(n_1172)
);

AO21x1_ASAP7_75t_L g1173 ( 
.A1(n_942),
.A2(n_924),
.B(n_937),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_937),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_950),
.A2(n_758),
.B(n_618),
.C(n_861),
.Y(n_1175)
);

OA21x2_ASAP7_75t_L g1176 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_993),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_941),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_941),
.Y(n_1178)
);

AO31x2_ASAP7_75t_L g1179 ( 
.A1(n_951),
.A2(n_960),
.A3(n_1048),
.B(n_942),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1038),
.B(n_854),
.Y(n_1180)
);

NOR2xp67_ASAP7_75t_L g1181 ( 
.A(n_947),
.B(n_491),
.Y(n_1181)
);

BUFx10_ASAP7_75t_L g1182 ( 
.A(n_969),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1038),
.B(n_854),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_954),
.A2(n_861),
.B1(n_305),
.B2(n_330),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_948),
.B(n_491),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1066),
.A2(n_867),
.B(n_1049),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1066),
.A2(n_867),
.B(n_1049),
.Y(n_1187)
);

AO32x2_ASAP7_75t_L g1188 ( 
.A1(n_1031),
.A2(n_942),
.A3(n_923),
.B1(n_1028),
.B2(n_1048),
.Y(n_1188)
);

AO31x2_ASAP7_75t_L g1189 ( 
.A1(n_951),
.A2(n_960),
.A3(n_1048),
.B(n_942),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_950),
.A2(n_758),
.B(n_618),
.C(n_861),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_L g1191 ( 
.A1(n_942),
.A2(n_758),
.B(n_658),
.C(n_657),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1026),
.B(n_491),
.Y(n_1192)
);

INVx4_ASAP7_75t_L g1193 ( 
.A(n_947),
.Y(n_1193)
);

INVx2_ASAP7_75t_SL g1194 ( 
.A(n_963),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1026),
.B(n_861),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1038),
.B(n_854),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_947),
.B(n_491),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1026),
.B(n_491),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1026),
.B(n_491),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1051),
.Y(n_1200)
);

OA21x2_ASAP7_75t_L g1201 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_993),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_937),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1027),
.B(n_1035),
.Y(n_1203)
);

AO22x2_ASAP7_75t_L g1204 ( 
.A1(n_942),
.A2(n_1031),
.B1(n_758),
.B2(n_950),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_947),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1027),
.B(n_1035),
.Y(n_1206)
);

AND2x6_ASAP7_75t_SL g1207 ( 
.A(n_1004),
.B(n_992),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_937),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1068),
.A2(n_1076),
.B(n_937),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_957),
.A2(n_861),
.B1(n_660),
.B2(n_1065),
.Y(n_1210)
);

AOI221x1_ASAP7_75t_L g1211 ( 
.A1(n_942),
.A2(n_1004),
.B1(n_1031),
.B2(n_924),
.C(n_951),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_957),
.A2(n_861),
.B1(n_660),
.B2(n_1065),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_948),
.B(n_491),
.Y(n_1213)
);

O2A1O1Ixp5_ASAP7_75t_SL g1214 ( 
.A1(n_942),
.A2(n_598),
.B(n_758),
.C(n_608),
.Y(n_1214)
);

NAND3xp33_ASAP7_75t_L g1215 ( 
.A(n_1004),
.B(n_518),
.C(n_861),
.Y(n_1215)
);

AND2x2_ASAP7_75t_L g1216 ( 
.A(n_1026),
.B(n_491),
.Y(n_1216)
);

INVx1_ASAP7_75t_SL g1217 ( 
.A(n_1129),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1191),
.A2(n_1215),
.B(n_1190),
.Y(n_1218)
);

INVx4_ASAP7_75t_L g1219 ( 
.A(n_1107),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1172),
.A2(n_1212),
.B1(n_1210),
.B2(n_1173),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1139),
.B(n_1086),
.Y(n_1221)
);

NOR2x1_ASAP7_75t_SL g1222 ( 
.A(n_1151),
.B(n_1125),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1175),
.A2(n_1211),
.B(n_1126),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1123),
.A2(n_1138),
.B(n_1127),
.Y(n_1224)
);

INVx3_ASAP7_75t_L g1225 ( 
.A(n_1166),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1081),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1137),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1087),
.Y(n_1228)
);

OR2x2_ASAP7_75t_L g1229 ( 
.A(n_1180),
.B(n_1183),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1193),
.B(n_1181),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1114),
.A2(n_1103),
.B(n_1096),
.C(n_1212),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1153),
.A2(n_1095),
.B(n_1098),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1133),
.B(n_1192),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1198),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1172),
.A2(n_1210),
.B(n_1093),
.C(n_1102),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1134),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1199),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1216),
.B(n_1091),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_1177),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1119),
.B(n_1161),
.Y(n_1240)
);

OAI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1115),
.A2(n_1132),
.B(n_1121),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1116),
.B(n_1112),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1104),
.A2(n_1122),
.B(n_1110),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1147),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1106),
.B(n_1102),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1174),
.A2(n_1209),
.B(n_1208),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_SL g1247 ( 
.A1(n_1105),
.A2(n_1142),
.B(n_1145),
.C(n_1085),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1108),
.B(n_1194),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1184),
.A2(n_1150),
.B1(n_1185),
.B2(n_1213),
.Y(n_1249)
);

HB1xp67_ASAP7_75t_L g1250 ( 
.A(n_1160),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1196),
.A2(n_1152),
.B1(n_1130),
.B2(n_1084),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1101),
.B(n_1170),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1174),
.A2(n_1209),
.B(n_1208),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_SL g1254 ( 
.A1(n_1161),
.A2(n_1159),
.B(n_1105),
.Y(n_1254)
);

OA21x2_ASAP7_75t_L g1255 ( 
.A1(n_1096),
.A2(n_1103),
.B(n_1202),
.Y(n_1255)
);

CKINVDCx6p67_ASAP7_75t_R g1256 ( 
.A(n_1082),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1205),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1178),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1134),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1171),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1167),
.Y(n_1261)
);

AO21x2_ASAP7_75t_L g1262 ( 
.A1(n_1115),
.A2(n_1124),
.B(n_1083),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1146),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1203),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1169),
.B(n_1214),
.Y(n_1265)
);

AO21x2_ASAP7_75t_L g1266 ( 
.A1(n_1141),
.A2(n_1118),
.B(n_1085),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1206),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1206),
.B(n_1089),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1094),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1204),
.A2(n_1100),
.B1(n_1195),
.B2(n_1113),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1094),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1099),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1143),
.A2(n_1158),
.B1(n_1204),
.B2(n_1088),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1156),
.A2(n_1090),
.B(n_1201),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1119),
.B(n_1163),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1135),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1197),
.A2(n_1145),
.B1(n_1182),
.B2(n_1164),
.Y(n_1277)
);

BUFx2_ASAP7_75t_R g1278 ( 
.A(n_1120),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1176),
.A2(n_1201),
.B(n_1149),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1099),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1097),
.B(n_1131),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1168),
.B(n_1136),
.Y(n_1282)
);

AOI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1144),
.A2(n_1193),
.B1(n_1155),
.B2(n_1200),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1200),
.Y(n_1284)
);

BUFx2_ASAP7_75t_SL g1285 ( 
.A(n_1166),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1092),
.A2(n_1109),
.B(n_1111),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1179),
.A2(n_1189),
.A3(n_1157),
.B(n_1188),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1140),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1154),
.A2(n_1165),
.B(n_1189),
.Y(n_1289)
);

OA21x2_ASAP7_75t_L g1290 ( 
.A1(n_1179),
.A2(n_1128),
.B(n_1188),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1154),
.A2(n_1165),
.B(n_1128),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1128),
.A2(n_1148),
.B(n_1162),
.Y(n_1292)
);

OAI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1207),
.A2(n_1191),
.B(n_1215),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1140),
.B(n_1180),
.Y(n_1294)
);

INVx4_ASAP7_75t_L g1295 ( 
.A(n_1107),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1096),
.A2(n_1103),
.B(n_1174),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1129),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1116),
.B(n_1067),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1177),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1191),
.A2(n_1215),
.B(n_830),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1133),
.B(n_1216),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1081),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1139),
.B(n_1086),
.Y(n_1303)
);

CKINVDCx11_ASAP7_75t_R g1304 ( 
.A(n_1082),
.Y(n_1304)
);

AOI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1215),
.A2(n_305),
.B1(n_330),
.B2(n_317),
.Y(n_1305)
);

OAI22xp5_ASAP7_75t_L g1306 ( 
.A1(n_1215),
.A2(n_861),
.B1(n_1184),
.B2(n_830),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1096),
.A2(n_1103),
.B(n_1174),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1080),
.A2(n_1187),
.B(n_1186),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1215),
.B(n_861),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1081),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1173),
.A2(n_1211),
.A3(n_1121),
.B(n_1092),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1119),
.B(n_1161),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1081),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1191),
.A2(n_1004),
.B(n_690),
.C(n_680),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1080),
.A2(n_1187),
.B(n_1186),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1215),
.A2(n_1004),
.B1(n_690),
.B2(n_680),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1116),
.B(n_1067),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1215),
.A2(n_1004),
.B1(n_690),
.B2(n_680),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1080),
.A2(n_1187),
.B(n_1186),
.Y(n_1319)
);

OR2x2_ASAP7_75t_L g1320 ( 
.A(n_1139),
.B(n_1086),
.Y(n_1320)
);

INVx4_ASAP7_75t_L g1321 ( 
.A(n_1107),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1081),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1081),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1081),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1107),
.Y(n_1325)
);

INVx8_ASAP7_75t_L g1326 ( 
.A(n_1107),
.Y(n_1326)
);

AOI222xp33_ASAP7_75t_L g1327 ( 
.A1(n_1215),
.A2(n_1004),
.B1(n_538),
.B2(n_866),
.C1(n_755),
.C2(n_923),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1215),
.A2(n_305),
.B1(n_330),
.B2(n_317),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1096),
.A2(n_1103),
.B(n_1174),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1249),
.B2(n_1314),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1240),
.B(n_1312),
.Y(n_1331)
);

AND2x2_ASAP7_75t_L g1332 ( 
.A(n_1248),
.B(n_1233),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1229),
.B(n_1252),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1314),
.B2(n_1220),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1279),
.A2(n_1265),
.B(n_1241),
.Y(n_1335)
);

AND2x2_ASAP7_75t_SL g1336 ( 
.A(n_1255),
.B(n_1296),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1301),
.B(n_1221),
.Y(n_1337)
);

A2O1A1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1231),
.A2(n_1223),
.B(n_1218),
.C(n_1293),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1303),
.B(n_1320),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1252),
.B(n_1268),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_1326),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1275),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1238),
.B(n_1282),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1281),
.B(n_1245),
.Y(n_1344)
);

NOR2xp67_ASAP7_75t_L g1345 ( 
.A(n_1294),
.B(n_1288),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1220),
.A2(n_1309),
.B1(n_1273),
.B2(n_1277),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1234),
.B(n_1237),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1309),
.A2(n_1306),
.B1(n_1328),
.B2(n_1305),
.Y(n_1348)
);

OA21x2_ASAP7_75t_L g1349 ( 
.A1(n_1274),
.A2(n_1246),
.B(n_1253),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1231),
.A2(n_1251),
.B1(n_1283),
.B2(n_1217),
.Y(n_1350)
);

INVx2_ASAP7_75t_SL g1351 ( 
.A(n_1228),
.Y(n_1351)
);

BUFx8_ASAP7_75t_SL g1352 ( 
.A(n_1258),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1236),
.B(n_1259),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_SL g1354 ( 
.A1(n_1255),
.A2(n_1329),
.B(n_1296),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1245),
.B(n_1297),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1242),
.A2(n_1270),
.B1(n_1317),
.B2(n_1298),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1260),
.B(n_1264),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1250),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1255),
.A2(n_1329),
.B(n_1296),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1307),
.A2(n_1329),
.B(n_1222),
.Y(n_1360)
);

CKINVDCx12_ASAP7_75t_R g1361 ( 
.A(n_1278),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1312),
.B(n_1227),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1263),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1260),
.B(n_1264),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1253),
.A2(n_1286),
.B(n_1243),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1300),
.B(n_1327),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1235),
.A2(n_1247),
.B(n_1242),
.C(n_1254),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_SL g1369 ( 
.A1(n_1276),
.A2(n_1299),
.B1(n_1239),
.B2(n_1284),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1275),
.B(n_1244),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1244),
.B(n_1302),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1298),
.A2(n_1317),
.B1(n_1307),
.B2(n_1325),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_1313),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1226),
.B(n_1324),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1304),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1269),
.A2(n_1272),
.B(n_1280),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1269),
.B(n_1272),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1325),
.A2(n_1257),
.B1(n_1219),
.B2(n_1321),
.Y(n_1379)
);

AOI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1262),
.A2(n_1230),
.B1(n_1266),
.B2(n_1261),
.C(n_1276),
.Y(n_1380)
);

O2A1O1Ixp5_ASAP7_75t_L g1381 ( 
.A1(n_1225),
.A2(n_1219),
.B(n_1321),
.C(n_1295),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1290),
.A2(n_1295),
.B(n_1262),
.Y(n_1382)
);

O2A1O1Ixp5_ASAP7_75t_L g1383 ( 
.A1(n_1225),
.A2(n_1311),
.B(n_1287),
.C(n_1292),
.Y(n_1383)
);

AOI221xp5_ASAP7_75t_L g1384 ( 
.A1(n_1239),
.A2(n_1299),
.B1(n_1326),
.B2(n_1311),
.C(n_1285),
.Y(n_1384)
);

CKINVDCx16_ASAP7_75t_R g1385 ( 
.A(n_1258),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1289),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1287),
.B(n_1311),
.Y(n_1387)
);

A2O1A1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1292),
.A2(n_1243),
.B(n_1291),
.C(n_1289),
.Y(n_1388)
);

OA21x2_ASAP7_75t_L g1389 ( 
.A1(n_1308),
.A2(n_1319),
.B(n_1315),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1287),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1256),
.A2(n_1304),
.B1(n_1311),
.B2(n_1287),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1232),
.B(n_1308),
.Y(n_1392)
);

OA21x2_ASAP7_75t_L g1393 ( 
.A1(n_1319),
.A2(n_1279),
.B(n_1265),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1229),
.B(n_1252),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1314),
.A2(n_1318),
.B(n_1316),
.C(n_1293),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1215),
.B2(n_861),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1248),
.B(n_1233),
.Y(n_1397)
);

NAND4xp25_ASAP7_75t_L g1398 ( 
.A(n_1316),
.B(n_1215),
.C(n_1318),
.D(n_400),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1215),
.B2(n_861),
.Y(n_1399)
);

AOI221xp5_ASAP7_75t_L g1400 ( 
.A1(n_1316),
.A2(n_1318),
.B1(n_1215),
.B2(n_1004),
.C(n_1314),
.Y(n_1400)
);

O2A1O1Ixp5_ASAP7_75t_L g1401 ( 
.A1(n_1314),
.A2(n_1173),
.B(n_1224),
.C(n_1241),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_SL g1402 ( 
.A1(n_1314),
.A2(n_467),
.B(n_1211),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1314),
.A2(n_1318),
.B(n_1316),
.C(n_1293),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1229),
.B(n_1252),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1248),
.B(n_1233),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1314),
.A2(n_1318),
.B(n_1316),
.C(n_1293),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1250),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_1358),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1358),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1342),
.B(n_1331),
.Y(n_1410)
);

BUFx6f_ASAP7_75t_L g1411 ( 
.A(n_1336),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1354),
.B(n_1359),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1407),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1407),
.Y(n_1415)
);

BUFx4f_ASAP7_75t_SL g1416 ( 
.A(n_1375),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1401),
.A2(n_1388),
.B(n_1383),
.Y(n_1417)
);

AO21x2_ASAP7_75t_L g1418 ( 
.A1(n_1360),
.A2(n_1338),
.B(n_1382),
.Y(n_1418)
);

INVx3_ASAP7_75t_L g1419 ( 
.A(n_1392),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1387),
.B(n_1344),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1351),
.Y(n_1421)
);

AO21x2_ASAP7_75t_L g1422 ( 
.A1(n_1360),
.A2(n_1338),
.B(n_1382),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1333),
.B(n_1394),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1386),
.A2(n_1402),
.B(n_1330),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1340),
.B(n_1404),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1335),
.B(n_1370),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1392),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1370),
.B(n_1362),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1335),
.B(n_1390),
.Y(n_1430)
);

OR2x6_ASAP7_75t_L g1431 ( 
.A(n_1376),
.B(n_1368),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1366),
.A2(n_1400),
.B1(n_1334),
.B2(n_1399),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1349),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1355),
.Y(n_1434)
);

OR2x6_ASAP7_75t_L g1435 ( 
.A(n_1376),
.B(n_1372),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1348),
.B(n_1337),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1377),
.B(n_1353),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1395),
.B(n_1406),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1377),
.B(n_1367),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1357),
.B(n_1364),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1391),
.B(n_1335),
.Y(n_1441)
);

BUFx2_ASAP7_75t_L g1442 ( 
.A(n_1365),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1365),
.B(n_1339),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1366),
.B(n_1373),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1373),
.B(n_1380),
.Y(n_1445)
);

INVxp67_ASAP7_75t_L g1446 ( 
.A(n_1408),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1416),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1433),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1427),
.B(n_1419),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1432),
.A2(n_1396),
.B1(n_1403),
.B2(n_1346),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1418),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1408),
.Y(n_1452)
);

INVxp67_ASAP7_75t_L g1453 ( 
.A(n_1444),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1412),
.B(n_1393),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1412),
.B(n_1393),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1443),
.B(n_1441),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1426),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1432),
.A2(n_1398),
.B1(n_1350),
.B2(n_1384),
.C(n_1356),
.Y(n_1458)
);

HB1xp67_ASAP7_75t_L g1459 ( 
.A(n_1426),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1412),
.B(n_1389),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1413),
.B(n_1442),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1414),
.Y(n_1462)
);

INVx4_ASAP7_75t_L g1463 ( 
.A(n_1431),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1414),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1428),
.B(n_1371),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1418),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1411),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1457),
.Y(n_1468)
);

AOI222xp33_ASAP7_75t_L g1469 ( 
.A1(n_1450),
.A2(n_1436),
.B1(n_1423),
.B2(n_1445),
.C1(n_1444),
.C2(n_1425),
.Y(n_1469)
);

AOI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1450),
.A2(n_1438),
.B(n_1431),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1450),
.A2(n_1438),
.B1(n_1425),
.B2(n_1345),
.C(n_1445),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1456),
.B(n_1420),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1448),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1458),
.A2(n_1438),
.B1(n_1418),
.B2(n_1422),
.Y(n_1474)
);

OAI31xp33_ASAP7_75t_L g1475 ( 
.A1(n_1458),
.A2(n_1438),
.A3(n_1441),
.B(n_1379),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1467),
.A2(n_1438),
.B1(n_1418),
.B2(n_1422),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1457),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1453),
.A2(n_1434),
.B1(n_1437),
.B2(n_1439),
.C(n_1343),
.Y(n_1478)
);

OAI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1453),
.A2(n_1438),
.B1(n_1435),
.B2(n_1434),
.C(n_1437),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1451),
.B(n_1347),
.C(n_1417),
.Y(n_1480)
);

AOI33xp33_ASAP7_75t_L g1481 ( 
.A1(n_1461),
.A2(n_1332),
.A3(n_1397),
.B1(n_1405),
.B2(n_1413),
.B3(n_1415),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_L g1482 ( 
.A1(n_1451),
.A2(n_1439),
.B1(n_1440),
.B2(n_1422),
.C(n_1378),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1449),
.B(n_1411),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1463),
.A2(n_1431),
.B1(n_1424),
.B2(n_1422),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1459),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1459),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_R g1487 ( 
.A(n_1447),
.B(n_1361),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1465),
.B(n_1429),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1465),
.B(n_1429),
.Y(n_1489)
);

NOR2xp67_ASAP7_75t_L g1490 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1456),
.B(n_1461),
.Y(n_1491)
);

OAI221xp5_ASAP7_75t_SL g1492 ( 
.A1(n_1456),
.A2(n_1431),
.B1(n_1435),
.B2(n_1420),
.C(n_1430),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1462),
.Y(n_1493)
);

CKINVDCx14_ASAP7_75t_R g1494 ( 
.A(n_1447),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1449),
.B(n_1411),
.Y(n_1495)
);

AOI21xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1461),
.A2(n_1385),
.B(n_1369),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1462),
.Y(n_1497)
);

AOI221xp5_ASAP7_75t_L g1498 ( 
.A1(n_1451),
.A2(n_1440),
.B1(n_1374),
.B2(n_1421),
.C(n_1409),
.Y(n_1498)
);

OAI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1446),
.A2(n_1381),
.B(n_1435),
.Y(n_1499)
);

HB1xp67_ASAP7_75t_L g1500 ( 
.A(n_1493),
.Y(n_1500)
);

AOI31xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1469),
.A2(n_1482),
.A3(n_1474),
.B(n_1470),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1483),
.B(n_1461),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1497),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1449),
.Y(n_1504)
);

INVx4_ASAP7_75t_SL g1505 ( 
.A(n_1468),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1468),
.Y(n_1506)
);

OA21x2_ASAP7_75t_L g1507 ( 
.A1(n_1480),
.A2(n_1442),
.B(n_1454),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1477),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1477),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1480),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1485),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1496),
.B(n_1410),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1485),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1494),
.B(n_1352),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1486),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1473),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1495),
.B(n_1449),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1472),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1472),
.Y(n_1521)
);

NAND3xp33_ASAP7_75t_SL g1522 ( 
.A(n_1475),
.B(n_1454),
.C(n_1455),
.Y(n_1522)
);

NAND3xp33_ASAP7_75t_L g1523 ( 
.A(n_1475),
.B(n_1451),
.C(n_1466),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1495),
.B(n_1467),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1478),
.B(n_1464),
.Y(n_1525)
);

INVx4_ASAP7_75t_SL g1526 ( 
.A(n_1487),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.Y(n_1527)
);

INVx1_ASAP7_75t_SL g1528 ( 
.A(n_1503),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1500),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1506),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1521),
.B(n_1491),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_SL g1532 ( 
.A(n_1526),
.B(n_1496),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1516),
.B(n_1352),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1525),
.B(n_1481),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1506),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1502),
.B(n_1490),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1508),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1490),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1502),
.B(n_1504),
.Y(n_1539)
);

NAND5xp2_ASAP7_75t_SL g1540 ( 
.A(n_1501),
.B(n_1471),
.C(n_1479),
.D(n_1476),
.E(n_1498),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1525),
.B(n_1464),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1521),
.B(n_1452),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1500),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1520),
.B(n_1488),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1526),
.B(n_1363),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1520),
.B(n_1489),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1503),
.B(n_1510),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1519),
.B(n_1527),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1510),
.B(n_1465),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1508),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1509),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1524),
.B(n_1460),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1509),
.Y(n_1554)
);

INVx4_ASAP7_75t_SL g1555 ( 
.A(n_1510),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1511),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1524),
.B(n_1505),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1511),
.B(n_1514),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1514),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1518),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1510),
.B(n_1465),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1505),
.B(n_1460),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1515),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1528),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1534),
.A2(n_1523),
.B(n_1522),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1548),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1528),
.B(n_1510),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1541),
.B(n_1522),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1545),
.B(n_1526),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1543),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1510),
.Y(n_1575)
);

INVx1_ASAP7_75t_SL g1576 ( 
.A(n_1532),
.Y(n_1576)
);

OAI21xp33_ASAP7_75t_L g1577 ( 
.A1(n_1540),
.A2(n_1523),
.B(n_1510),
.Y(n_1577)
);

AND2x4_ASAP7_75t_L g1578 ( 
.A(n_1555),
.B(n_1505),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1512),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1548),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1547),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1546),
.B(n_1513),
.Y(n_1582)
);

OAI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1540),
.A2(n_1513),
.B1(n_1501),
.B2(n_1484),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1555),
.B(n_1517),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1555),
.B(n_1517),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1555),
.B(n_1505),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1555),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1530),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1542),
.B(n_1507),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1542),
.B(n_1507),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1530),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_L g1593 ( 
.A(n_1549),
.B(n_1451),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1550),
.A2(n_1513),
.B(n_1492),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1535),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1549),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1535),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1531),
.B(n_1513),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1558),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1565),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1583),
.B(n_1539),
.Y(n_1601)
);

CKINVDCx16_ASAP7_75t_R g1602 ( 
.A(n_1567),
.Y(n_1602)
);

INVx2_ASAP7_75t_SL g1603 ( 
.A(n_1578),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1539),
.Y(n_1605)
);

CKINVDCx16_ASAP7_75t_R g1606 ( 
.A(n_1570),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1553),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1599),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1570),
.B(n_1549),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.B(n_1563),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1588),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1572),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1591),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1563),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1595),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1568),
.Y(n_1618)
);

OR2x6_ASAP7_75t_L g1619 ( 
.A(n_1586),
.B(n_1513),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1580),
.B(n_1558),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1580),
.B(n_1574),
.Y(n_1621)
);

BUFx2_ASAP7_75t_L g1622 ( 
.A(n_1587),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1596),
.B(n_1536),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1577),
.B(n_1507),
.C(n_1513),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1600),
.B(n_1533),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1624),
.A2(n_1566),
.B(n_1569),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1609),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1622),
.B(n_1581),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1618),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1604),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1611),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1611),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1602),
.B(n_1573),
.C(n_1575),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1604),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1604),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1602),
.B(n_1571),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1611),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1601),
.A2(n_1594),
.B(n_1573),
.Y(n_1638)
);

AOI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1624),
.A2(n_1593),
.B(n_1584),
.C(n_1585),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1614),
.A2(n_1593),
.B1(n_1597),
.B2(n_1589),
.C(n_1590),
.Y(n_1640)
);

NAND2x1p5_ASAP7_75t_L g1641 ( 
.A(n_1622),
.B(n_1507),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_SL g1642 ( 
.A(n_1606),
.B(n_1579),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1606),
.B(n_1598),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1630),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1631),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1636),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1634),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1635),
.Y(n_1648)
);

NOR2x1_ASAP7_75t_L g1649 ( 
.A(n_1632),
.B(n_1621),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1628),
.B(n_1621),
.Y(n_1650)
);

NOR2x1_ASAP7_75t_L g1651 ( 
.A(n_1637),
.B(n_1628),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1627),
.B(n_1603),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1629),
.B(n_1603),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1613),
.Y(n_1654)
);

NAND4xp25_ASAP7_75t_L g1655 ( 
.A(n_1646),
.B(n_1638),
.C(n_1633),
.D(n_1642),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1649),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1650),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_SL g1658 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1653),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1645),
.B(n_1625),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1654),
.A2(n_1607),
.B1(n_1643),
.B2(n_1639),
.C(n_1640),
.Y(n_1661)
);

OAI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1654),
.A2(n_1640),
.B(n_1641),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1652),
.B(n_1610),
.C(n_1613),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1644),
.A2(n_1619),
.B1(n_1610),
.B2(n_1605),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1658),
.A2(n_1647),
.B(n_1648),
.C(n_1615),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1656),
.B(n_1615),
.Y(n_1666)
);

XNOR2xp5_ASAP7_75t_L g1667 ( 
.A(n_1655),
.B(n_1605),
.Y(n_1667)
);

A2O1A1Ixp33_ASAP7_75t_SL g1668 ( 
.A1(n_1662),
.A2(n_1617),
.B(n_1612),
.C(n_1616),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1661),
.A2(n_1608),
.B1(n_1612),
.B2(n_1616),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1657),
.Y(n_1670)
);

INVxp67_ASAP7_75t_L g1671 ( 
.A(n_1667),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1669),
.B(n_1664),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1670),
.B(n_1660),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1666),
.B(n_1659),
.Y(n_1674)
);

NAND2xp33_ASAP7_75t_L g1675 ( 
.A(n_1668),
.B(n_1663),
.Y(n_1675)
);

INVxp67_ASAP7_75t_L g1676 ( 
.A(n_1665),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1669),
.B(n_1623),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_SL g1678 ( 
.A(n_1674),
.B(n_1641),
.C(n_1617),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1675),
.A2(n_1608),
.B(n_1620),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1676),
.A2(n_1619),
.B(n_1590),
.C(n_1608),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1677),
.Y(n_1681)
);

XOR2xp5_ASAP7_75t_L g1682 ( 
.A(n_1672),
.B(n_1608),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1682),
.Y(n_1683)
);

NOR3x1_ASAP7_75t_L g1684 ( 
.A(n_1678),
.B(n_1673),
.C(n_1671),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_1623),
.C(n_1620),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1685),
.Y(n_1686)
);

AOI322xp5_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1683),
.A3(n_1684),
.B1(n_1679),
.B2(n_1680),
.C1(n_1562),
.C2(n_1538),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1687),
.A2(n_1582),
.B1(n_1619),
.B2(n_1592),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1687),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1689),
.Y(n_1690)
);

INVx2_ASAP7_75t_SL g1691 ( 
.A(n_1688),
.Y(n_1691)
);

BUFx2_ASAP7_75t_L g1692 ( 
.A(n_1691),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1690),
.A2(n_1619),
.B1(n_1592),
.B2(n_1559),
.Y(n_1693)
);

OAI22x1_ASAP7_75t_L g1694 ( 
.A1(n_1692),
.A2(n_1560),
.B1(n_1564),
.B2(n_1552),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_SL g1695 ( 
.A1(n_1694),
.A2(n_1693),
.B1(n_1361),
.B2(n_1619),
.Y(n_1695)
);

XOR2xp5_ASAP7_75t_L g1696 ( 
.A(n_1695),
.B(n_1341),
.Y(n_1696)
);

AOI22x1_ASAP7_75t_L g1697 ( 
.A1(n_1696),
.A2(n_1560),
.B1(n_1561),
.B2(n_1564),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1697),
.A2(n_1537),
.B1(n_1551),
.B2(n_1559),
.Y(n_1698)
);

AOI211xp5_ASAP7_75t_L g1699 ( 
.A1(n_1698),
.A2(n_1561),
.B(n_1556),
.C(n_1554),
.Y(n_1699)
);


endmodule