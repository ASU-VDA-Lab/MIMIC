module fake_aes_1058_n_715 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_715);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_715;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_L g79 ( .A(n_64), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_1), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_72), .Y(n_81) );
BUFx6f_ASAP7_75t_L g82 ( .A(n_17), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_67), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_13), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_17), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_32), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_2), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_24), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_11), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_57), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_68), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_59), .Y(n_93) );
CKINVDCx14_ASAP7_75t_R g94 ( .A(n_36), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_46), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_34), .Y(n_96) );
NOR2xp33_ASAP7_75t_L g97 ( .A(n_43), .B(n_1), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_56), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_39), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_52), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_66), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_69), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_21), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_40), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_73), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_33), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_38), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_27), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_62), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_19), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_22), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_26), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_18), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_20), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_10), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_11), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
INVx1_ASAP7_75t_SL g124 ( .A(n_37), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_22), .Y(n_125) );
INVxp33_ASAP7_75t_L g126 ( .A(n_15), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_61), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_111), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_86), .A2(n_29), .B(n_76), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_122), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_94), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_93), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_110), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx3_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
NOR2xp33_ASAP7_75t_R g139 ( .A(n_109), .B(n_28), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_82), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_81), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_101), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_126), .B(n_0), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_91), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_120), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g146 ( .A(n_116), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_91), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_101), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_80), .B(n_0), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_124), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_92), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_106), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_80), .B(n_2), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_112), .B(n_3), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_82), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_98), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_95), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_95), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_108), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_96), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_99), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_82), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_112), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_99), .Y(n_166) );
AND2x4_ASAP7_75t_L g167 ( .A(n_84), .B(n_3), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_100), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_108), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_100), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_82), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_167), .B(n_84), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_152), .B(n_157), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_138), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_138), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
AOI22xp5_ASAP7_75t_L g181 ( .A1(n_158), .A2(n_117), .B1(n_125), .B2(n_90), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_165), .B(n_79), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_130), .B(n_127), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_154), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_167), .B(n_85), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
NAND3xp33_ASAP7_75t_L g187 ( .A(n_159), .B(n_89), .C(n_125), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_130), .B(n_127), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_131), .B(n_123), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_131), .B(n_123), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_129), .Y(n_194) );
OR2x2_ASAP7_75t_L g195 ( .A(n_143), .B(n_104), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
NAND2x1p5_ASAP7_75t_L g200 ( .A(n_167), .B(n_104), .Y(n_200) );
INVx1_ASAP7_75t_SL g201 ( .A(n_146), .Y(n_201) );
NOR2xp33_ASAP7_75t_SL g202 ( .A(n_134), .B(n_121), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_138), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_155), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_167), .B(n_85), .Y(n_205) );
NAND3x1_ASAP7_75t_L g206 ( .A(n_137), .B(n_87), .C(n_119), .Y(n_206) );
OR2x2_ASAP7_75t_L g207 ( .A(n_165), .B(n_90), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_137), .B(n_121), .Y(n_208) );
OR2x2_ASAP7_75t_L g209 ( .A(n_133), .B(n_119), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
AND2x6_ASAP7_75t_L g212 ( .A(n_144), .B(n_118), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_144), .Y(n_213) );
OAI22x1_ASAP7_75t_L g214 ( .A1(n_145), .A2(n_88), .B1(n_117), .B2(n_87), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_147), .B(n_89), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_168), .A2(n_114), .B1(n_82), .B2(n_97), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_128), .Y(n_217) );
NAND3x1_ASAP7_75t_L g218 ( .A(n_147), .B(n_114), .C(n_115), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_140), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_153), .B(n_118), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_140), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_153), .B(n_115), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_160), .B(n_102), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_140), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_162), .B(n_113), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_128), .Y(n_230) );
AOI22xp33_ASAP7_75t_SL g231 ( .A1(n_156), .A2(n_113), .B1(n_107), .B2(n_105), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_128), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_162), .B(n_170), .Y(n_233) );
INVxp33_ASAP7_75t_L g234 ( .A(n_163), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_141), .Y(n_235) );
INVx1_ASAP7_75t_SL g236 ( .A(n_164), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_234), .B(n_135), .Y(n_237) );
OR2x6_ASAP7_75t_L g238 ( .A(n_194), .B(n_170), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_201), .Y(n_239) );
INVxp67_ASAP7_75t_SL g240 ( .A(n_200), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_233), .Y(n_241) );
OR2x2_ASAP7_75t_L g242 ( .A(n_182), .B(n_209), .Y(n_242) );
AOI211xp5_ASAP7_75t_L g243 ( .A1(n_209), .A2(n_150), .B(n_166), .C(n_163), .Y(n_243) );
NOR3xp33_ASAP7_75t_SL g244 ( .A(n_174), .B(n_136), .C(n_166), .Y(n_244) );
NOR2xp33_ASAP7_75t_R g245 ( .A(n_194), .B(n_171), .Y(n_245) );
NAND2xp33_ASAP7_75t_SL g246 ( .A(n_234), .B(n_139), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_236), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_233), .B(n_148), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_200), .B(n_102), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_233), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_230), .Y(n_251) );
NOR3xp33_ASAP7_75t_SL g252 ( .A(n_174), .B(n_103), .C(n_105), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_172), .B(n_148), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
NOR3xp33_ASAP7_75t_SL g255 ( .A(n_187), .B(n_103), .C(n_107), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_182), .Y(n_256) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_173), .A2(n_169), .B1(n_161), .B2(n_142), .Y(n_257) );
INVx3_ASAP7_75t_L g258 ( .A(n_211), .Y(n_258) );
BUFx2_ASAP7_75t_SL g259 ( .A(n_212), .Y(n_259) );
AND2x4_ASAP7_75t_L g260 ( .A(n_172), .B(n_169), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_211), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_212), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_232), .Y(n_263) );
AND3x2_ASAP7_75t_SL g264 ( .A(n_206), .B(n_169), .C(n_161), .Y(n_264) );
INVx1_ASAP7_75t_SL g265 ( .A(n_207), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_195), .B(n_161), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_195), .B(n_213), .Y(n_267) );
CKINVDCx14_ASAP7_75t_R g268 ( .A(n_212), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_219), .B(n_142), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_220), .B(n_142), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_177), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_207), .B(n_141), .Y(n_272) );
NOR3xp33_ASAP7_75t_SL g273 ( .A(n_188), .B(n_208), .C(n_225), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_232), .Y(n_274) );
NOR2xp33_ASAP7_75t_R g275 ( .A(n_202), .B(n_4), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_211), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_212), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_212), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_215), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_227), .B(n_141), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_231), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_172), .B(n_31), .Y(n_282) );
NOR2xp33_ASAP7_75t_R g283 ( .A(n_176), .B(n_5), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_235), .Y(n_284) );
BUFx2_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_215), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_179), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_185), .B(n_35), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_206), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_185), .B(n_6), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_185), .Y(n_291) );
OR2x6_ASAP7_75t_L g292 ( .A(n_214), .B(n_7), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_214), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_205), .B(n_7), .Y(n_294) );
NAND3xp33_ASAP7_75t_SL g295 ( .A(n_181), .B(n_8), .C(n_9), .Y(n_295) );
NOR2xp33_ASAP7_75t_R g296 ( .A(n_180), .B(n_9), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_205), .B(n_190), .Y(n_297) );
BUFx4f_ASAP7_75t_L g298 ( .A(n_226), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_205), .B(n_10), .Y(n_299) );
NOR3xp33_ASAP7_75t_SL g300 ( .A(n_188), .B(n_12), .C(n_13), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_184), .B(n_47), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_186), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_189), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g304 ( .A1(n_218), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_304) );
AND3x2_ASAP7_75t_SL g305 ( .A(n_218), .B(n_14), .C(n_16), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_251), .Y(n_306) );
OR2x2_ASAP7_75t_L g307 ( .A(n_265), .B(n_183), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_251), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_277), .B(n_196), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
BUFx3_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_238), .B(n_217), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_254), .Y(n_313) );
INVx3_ASAP7_75t_SL g314 ( .A(n_238), .Y(n_314) );
INVx1_ASAP7_75t_SL g315 ( .A(n_239), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_290), .A2(n_226), .B1(n_204), .B2(n_197), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_263), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_263), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
BUFx2_ASAP7_75t_L g320 ( .A(n_238), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_249), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_249), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_290), .A2(n_226), .B1(n_198), .B2(n_208), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_249), .Y(n_324) );
INVx2_ASAP7_75t_SL g325 ( .A(n_290), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_261), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_247), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g328 ( .A1(n_267), .A2(n_229), .B(n_192), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_240), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_271), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_287), .A2(n_177), .B(n_191), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_297), .B(n_226), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_301), .A2(n_222), .B(n_235), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_279), .B(n_217), .Y(n_335) );
INVxp67_ASAP7_75t_L g336 ( .A(n_247), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_245), .Y(n_337) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_268), .A2(n_291), .B1(n_250), .B2(n_241), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_276), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_274), .Y(n_340) );
NAND2xp5_ASAP7_75t_SL g341 ( .A(n_278), .B(n_216), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_286), .B(n_217), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_274), .Y(n_343) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_302), .A2(n_177), .B(n_191), .Y(n_344) );
INVx3_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
BUFx4f_ASAP7_75t_SL g346 ( .A(n_242), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_278), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_284), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_256), .B(n_226), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
CKINVDCx20_ASAP7_75t_R g351 ( .A(n_245), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_272), .B(n_226), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_266), .B(n_177), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_271), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_273), .B(n_210), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_303), .A2(n_191), .B1(n_193), .B2(n_210), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g358 ( .A1(n_295), .A2(n_191), .B1(n_193), .B2(n_210), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_268), .B(n_193), .Y(n_359) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_327), .A2(n_243), .B(n_252), .C(n_244), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_307), .B(n_260), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_320), .A2(n_275), .B1(n_293), .B2(n_296), .Y(n_362) );
NAND3xp33_ASAP7_75t_L g363 ( .A(n_358), .B(n_255), .C(n_300), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_307), .B(n_260), .Y(n_364) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_353), .A2(n_301), .B(n_294), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_346), .A2(n_289), .B1(n_293), .B2(n_283), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_336), .A2(n_237), .B1(n_281), .B2(n_246), .C(n_299), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_320), .A2(n_296), .B1(n_283), .B2(n_246), .Y(n_369) );
NAND2xp33_ASAP7_75t_R g370 ( .A(n_329), .B(n_275), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_306), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_315), .B(n_248), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_322), .B(n_276), .Y(n_373) );
OAI22xp33_ASAP7_75t_SL g374 ( .A1(n_314), .A2(n_292), .B1(n_304), .B2(n_305), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g375 ( .A(n_322), .B(n_298), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_314), .A2(n_260), .B1(n_253), .B2(n_258), .Y(n_377) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_331), .A2(n_271), .B(n_298), .Y(n_378) );
AND2x4_ASAP7_75t_SL g379 ( .A(n_321), .B(n_292), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_328), .A2(n_280), .B(n_270), .C(n_269), .Y(n_380) );
NAND2xp33_ASAP7_75t_R g381 ( .A(n_314), .B(n_292), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_322), .B(n_253), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_322), .B(n_321), .Y(n_384) );
INVx4_ASAP7_75t_L g385 ( .A(n_322), .Y(n_385) );
INVx4_ASAP7_75t_SL g386 ( .A(n_324), .Y(n_386) );
AOI21xp5_ASAP7_75t_L g387 ( .A1(n_344), .A2(n_288), .B(n_282), .Y(n_387) );
OAI22xp5_ASAP7_75t_L g388 ( .A1(n_322), .A2(n_253), .B1(n_259), .B2(n_257), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_324), .B(n_258), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_306), .Y(n_390) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_325), .A2(n_285), .B1(n_262), .B2(n_282), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_330), .A2(n_288), .B(n_210), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_361), .B(n_310), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_371), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_351), .B1(n_337), .B2(n_325), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_367), .A2(n_328), .B1(n_323), .B2(n_358), .C(n_349), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_368), .A2(n_316), .B1(n_332), .B2(n_355), .C(n_338), .Y(n_397) );
OAI21xp5_ASAP7_75t_SL g398 ( .A1(n_362), .A2(n_316), .B(n_312), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_369), .A2(n_352), .B1(n_317), .B2(n_348), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_385), .Y(n_400) );
OAI22xp33_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_305), .B1(n_312), .B2(n_348), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
AOI21xp5_ASAP7_75t_L g403 ( .A1(n_387), .A2(n_330), .B(n_356), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_374), .A2(n_264), .B1(n_342), .B2(n_335), .Y(n_404) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_380), .A2(n_353), .B(n_257), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_317), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
OAI332xp33_ASAP7_75t_L g408 ( .A1(n_366), .A2(n_264), .A3(n_350), .B1(n_310), .B2(n_343), .B3(n_326), .C1(n_340), .C2(n_308), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_371), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_363), .A2(n_343), .B(n_350), .C(n_333), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_377), .A2(n_357), .B1(n_306), .B2(n_308), .Y(n_411) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_361), .A2(n_335), .B1(n_342), .B2(n_341), .C(n_345), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_384), .Y(n_413) );
NAND4xp25_ASAP7_75t_L g414 ( .A(n_381), .B(n_342), .C(n_345), .D(n_339), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_364), .A2(n_342), .B1(n_345), .B2(n_339), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_364), .A2(n_339), .B1(n_345), .B2(n_333), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_390), .Y(n_417) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_392), .A2(n_357), .B(n_318), .Y(n_418) );
AOI322xp5_ASAP7_75t_L g419 ( .A1(n_376), .A2(n_340), .A3(n_318), .B1(n_308), .B2(n_21), .C1(n_23), .C2(n_24), .Y(n_419) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_379), .A2(n_334), .B1(n_333), .B2(n_319), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_417), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_401), .A2(n_379), .B1(n_382), .B2(n_383), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_417), .B(n_340), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_393), .B(n_365), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_398), .A2(n_382), .B1(n_388), .B2(n_385), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_402), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_404), .A2(n_385), .B1(n_389), .B2(n_334), .Y(n_428) );
OAI31xp33_ASAP7_75t_L g429 ( .A1(n_414), .A2(n_380), .A3(n_389), .B(n_375), .Y(n_429) );
NOR2xp33_ASAP7_75t_R g430 ( .A(n_402), .B(n_333), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_400), .Y(n_431) );
OAI221xp5_ASAP7_75t_L g432 ( .A1(n_398), .A2(n_391), .B1(n_318), .B2(n_334), .C(n_313), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_406), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_402), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_394), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g436 ( .A1(n_414), .A2(n_334), .B1(n_313), .B2(n_326), .C(n_375), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_394), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_407), .A2(n_389), .B1(n_373), .B2(n_386), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_413), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_393), .A2(n_373), .B1(n_386), .B2(n_193), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_412), .A2(n_373), .B1(n_386), .B2(n_339), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_421), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_421), .Y(n_443) );
INVx3_ASAP7_75t_L g444 ( .A(n_400), .Y(n_444) );
OAI31xp33_ASAP7_75t_L g445 ( .A1(n_396), .A2(n_319), .A3(n_359), .B(n_309), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_394), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_403), .A2(n_378), .B(n_359), .Y(n_448) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_409), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_397), .A2(n_386), .B1(n_319), .B2(n_311), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_406), .B(n_319), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_408), .B(n_356), .Y(n_454) );
INVx4_ASAP7_75t_L g455 ( .A(n_400), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_413), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_449), .B(n_420), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_449), .B(n_399), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_435), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_423), .B(n_395), .C(n_419), .D(n_415), .Y(n_461) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_433), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_431), .Y(n_463) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_433), .A2(n_408), .B1(n_405), .B2(n_416), .C(n_410), .Y(n_464) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_457), .A2(n_405), .B(n_411), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_436), .A2(n_419), .A3(n_311), .B(n_347), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_435), .B(n_418), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_422), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_431), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_430), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_439), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_422), .B(n_418), .Y(n_472) );
XNOR2xp5_ASAP7_75t_L g473 ( .A(n_423), .B(n_16), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_442), .B(n_418), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_442), .Y(n_475) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
OR2x6_ASAP7_75t_L g477 ( .A(n_455), .B(n_356), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_443), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_435), .B(n_18), .Y(n_480) );
BUFx3_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_435), .B(n_20), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_437), .Y(n_483) );
NAND4xp25_ASAP7_75t_L g484 ( .A(n_428), .B(n_432), .C(n_429), .D(n_445), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_437), .B(n_25), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_437), .B(n_25), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_437), .B(n_30), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_450), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_446), .B(n_356), .Y(n_489) );
AOI22xp33_ASAP7_75t_SL g490 ( .A1(n_430), .A2(n_311), .B1(n_347), .B2(n_354), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_446), .B(n_41), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_450), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_446), .B(n_44), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_456), .B(n_45), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_446), .B(n_49), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_457), .Y(n_498) );
NOR2xp67_ASAP7_75t_L g499 ( .A(n_436), .B(n_51), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_452), .B(n_53), .Y(n_500) );
NOR3xp33_ASAP7_75t_SL g501 ( .A(n_432), .B(n_54), .C(n_55), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_431), .B(n_354), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_457), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_447), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_455), .B(n_58), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_425), .A2(n_356), .B1(n_354), .B2(n_330), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_424), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_445), .A2(n_356), .B1(n_354), .B2(n_330), .C(n_199), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_507), .B(n_427), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_462), .B(n_427), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_468), .B(n_425), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_468), .B(n_457), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
INVx5_ASAP7_75t_L g515 ( .A(n_492), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_471), .B(n_427), .Y(n_516) );
OAI33xp33_ASAP7_75t_L g517 ( .A1(n_461), .A2(n_454), .A3(n_456), .B1(n_429), .B2(n_428), .B3(n_438), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_476), .Y(n_518) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_473), .B(n_440), .C(n_438), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_488), .B(n_427), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_478), .B(n_424), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_470), .Y(n_522) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_470), .B(n_455), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_488), .B(n_434), .Y(n_525) );
XNOR2xp5_ASAP7_75t_L g526 ( .A(n_473), .B(n_426), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_463), .B(n_424), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_461), .A2(n_441), .B1(n_454), .B2(n_426), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_493), .B(n_434), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_478), .B(n_448), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_492), .B(n_431), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_479), .B(n_448), .Y(n_532) );
NOR2xp33_ASAP7_75t_R g533 ( .A(n_463), .B(n_434), .Y(n_533) );
BUFx2_ASAP7_75t_L g534 ( .A(n_492), .Y(n_534) );
AOI211xp5_ASAP7_75t_L g535 ( .A1(n_484), .A2(n_453), .B(n_434), .C(n_447), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_469), .B(n_434), .Y(n_536) );
NAND4xp25_ASAP7_75t_SL g537 ( .A(n_466), .B(n_441), .C(n_440), .D(n_451), .Y(n_537) );
NAND4xp25_ASAP7_75t_L g538 ( .A(n_484), .B(n_451), .C(n_453), .D(n_447), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_479), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_493), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_497), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_497), .B(n_455), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_460), .B(n_455), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_492), .B(n_431), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_458), .Y(n_545) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_464), .B(n_453), .C(n_447), .D(n_444), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_469), .B(n_431), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_503), .B(n_448), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_480), .Y(n_549) );
AND2x2_ASAP7_75t_SL g550 ( .A(n_505), .B(n_444), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_505), .B(n_499), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_482), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_482), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_458), .Y(n_554) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_481), .B(n_444), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_485), .Y(n_556) );
NAND2x1p5_ASAP7_75t_SL g557 ( .A(n_485), .B(n_431), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_460), .B(n_444), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_460), .Y(n_559) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_495), .B(n_444), .C(n_199), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_503), .B(n_472), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_486), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_483), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_483), .B(n_448), .Y(n_564) );
NAND2x1_ASAP7_75t_L g565 ( .A(n_505), .B(n_354), .Y(n_565) );
NOR3xp33_ASAP7_75t_L g566 ( .A(n_486), .B(n_178), .C(n_228), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_483), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_481), .B(n_60), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_513), .Y(n_569) );
AO22x1_ASAP7_75t_L g570 ( .A1(n_515), .A2(n_481), .B1(n_505), .B2(n_504), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_534), .Y(n_571) );
NAND2xp5_ASAP7_75t_SL g572 ( .A(n_515), .B(n_499), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_518), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_514), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_517), .A2(n_464), .B1(n_466), .B2(n_459), .Y(n_575) );
AOI33xp33_ASAP7_75t_L g576 ( .A1(n_528), .A2(n_490), .A3(n_500), .B1(n_504), .B2(n_467), .B3(n_496), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_545), .B(n_459), .Y(n_577) );
AOI222xp33_ASAP7_75t_L g578 ( .A1(n_517), .A2(n_472), .B1(n_474), .B2(n_508), .C1(n_467), .C2(n_500), .Y(n_578) );
AOI322xp5_ASAP7_75t_L g579 ( .A1(n_545), .A2(n_501), .A3(n_474), .B1(n_496), .B2(n_494), .C1(n_491), .C2(n_487), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_539), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_559), .Y(n_581) );
OAI21xp33_ASAP7_75t_SL g582 ( .A1(n_550), .A2(n_477), .B(n_502), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_554), .B(n_498), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_554), .B(n_498), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_540), .Y(n_585) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_526), .A2(n_508), .B(n_490), .Y(n_586) );
AO22x2_ASAP7_75t_L g587 ( .A1(n_541), .A2(n_498), .B1(n_494), .B2(n_491), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_510), .B(n_477), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
NAND3x1_ASAP7_75t_L g590 ( .A(n_516), .B(n_506), .C(n_487), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_563), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_519), .A2(n_501), .B1(n_448), .B2(n_477), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_511), .B(n_465), .Y(n_593) );
NOR4xp25_ASAP7_75t_L g594 ( .A(n_537), .B(n_489), .C(n_465), .D(n_506), .Y(n_594) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_515), .B(n_489), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_538), .B(n_465), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_529), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_511), .B(n_465), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_509), .B(n_477), .Y(n_599) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_567), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_564), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_521), .B(n_477), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_530), .B(n_63), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_521), .B(n_65), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_546), .A2(n_537), .B(n_535), .C(n_551), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_530), .B(n_70), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_512), .Y(n_607) );
AOI222xp33_ASAP7_75t_L g608 ( .A1(n_524), .A2(n_221), .B1(n_228), .B2(n_224), .C1(n_175), .C2(n_178), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_543), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_549), .B(n_71), .Y(n_610) );
OAI322xp33_ASAP7_75t_L g611 ( .A1(n_532), .A2(n_224), .A3(n_175), .B1(n_203), .B2(n_223), .C1(n_221), .C2(n_74), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_512), .Y(n_612) );
AOI21xp33_ASAP7_75t_L g613 ( .A1(n_532), .A2(n_78), .B(n_330), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_527), .B(n_354), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_560), .A2(n_330), .B1(n_221), .B2(n_223), .Y(n_615) );
NAND3xp33_ASAP7_75t_L g616 ( .A(n_566), .B(n_221), .C(n_203), .Y(n_616) );
AOI321xp33_ASAP7_75t_L g617 ( .A1(n_552), .A2(n_556), .A3(n_562), .B1(n_553), .B2(n_560), .C(n_548), .Y(n_617) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_548), .B(n_515), .C(n_544), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_561), .B(n_558), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_561), .B(n_522), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_520), .B(n_542), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_589), .B(n_536), .Y(n_622) );
OAI211xp5_ASAP7_75t_L g623 ( .A1(n_582), .A2(n_533), .B(n_565), .C(n_568), .Y(n_623) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_605), .A2(n_531), .B1(n_555), .B2(n_547), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_601), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_612), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_612), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_619), .B(n_531), .Y(n_628) );
INVxp67_ASAP7_75t_SL g629 ( .A(n_600), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_569), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_574), .Y(n_631) );
OA21x2_ASAP7_75t_SL g632 ( .A1(n_572), .A2(n_557), .B(n_523), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_609), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_609), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_620), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_597), .B(n_619), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_583), .B(n_601), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_580), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_577), .B(n_607), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_621), .Y(n_641) );
AOI311xp33_ASAP7_75t_L g642 ( .A1(n_596), .A2(n_573), .A3(n_602), .B(n_571), .C(n_598), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_586), .B(n_599), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_583), .B(n_575), .Y(n_644) );
INVx1_ASAP7_75t_SL g645 ( .A(n_595), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_575), .B(n_578), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_596), .B(n_584), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_594), .B(n_600), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_587), .B(n_588), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_581), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_581), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_590), .A2(n_592), .B1(n_616), .B2(n_606), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_591), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_595), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_591), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_618), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_617), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g658 ( .A1(n_572), .A2(n_615), .B1(n_570), .B2(n_576), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_643), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_629), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_642), .B(n_576), .C(n_579), .Y(n_661) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_623), .A2(n_587), .B1(n_606), .B2(n_603), .Y(n_662) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_650), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_626), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_644), .B(n_593), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_630), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_650), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_630), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_626), .Y(n_669) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_646), .A2(n_603), .A3(n_604), .B1(n_610), .B2(n_614), .C1(n_590), .C2(n_613), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_631), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
INVxp67_ASAP7_75t_SL g673 ( .A(n_648), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_657), .B(n_587), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_658), .B(n_611), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_631), .Y(n_676) );
XOR2x2_ASAP7_75t_L g677 ( .A(n_624), .B(n_608), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_635), .B(n_647), .Y(n_678) );
INVx1_ASAP7_75t_SL g679 ( .A(n_633), .Y(n_679) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_641), .A2(n_656), .B1(n_634), .B2(n_649), .C1(n_640), .C2(n_639), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_638), .B(n_636), .Y(n_681) );
AO22x2_ASAP7_75t_L g682 ( .A1(n_673), .A2(n_656), .B1(n_645), .B2(n_649), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_659), .B(n_628), .Y(n_683) );
O2A1O1Ixp33_ASAP7_75t_L g684 ( .A1(n_675), .A2(n_654), .B(n_632), .C(n_627), .Y(n_684) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_679), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_660), .Y(n_686) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_667), .B(n_652), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_662), .A2(n_628), .B1(n_622), .B2(n_637), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_666), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_668), .Y(n_690) );
NOR4xp25_ASAP7_75t_L g691 ( .A(n_674), .B(n_653), .C(n_655), .D(n_651), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_671), .Y(n_692) );
OAI21xp5_ASAP7_75t_L g693 ( .A1(n_661), .A2(n_637), .B(n_653), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_665), .B(n_625), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_677), .A2(n_625), .B1(n_655), .B2(n_680), .Y(n_695) );
NOR2xp67_ASAP7_75t_L g696 ( .A(n_678), .B(n_681), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_670), .A2(n_677), .B(n_681), .C(n_676), .Y(n_697) );
NAND4xp25_ASAP7_75t_L g698 ( .A(n_664), .B(n_672), .C(n_669), .D(n_663), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_664), .B(n_669), .Y(n_699) );
BUFx6f_ASAP7_75t_L g700 ( .A(n_672), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_679), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g702 ( .A(n_701), .B(n_685), .Y(n_702) );
INVxp33_ASAP7_75t_SL g703 ( .A(n_686), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_683), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_684), .B(n_697), .C(n_695), .D(n_693), .Y(n_705) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_684), .A2(n_687), .B1(n_688), .B2(n_691), .C(n_698), .Y(n_706) );
XNOR2xp5_ASAP7_75t_L g707 ( .A(n_702), .B(n_682), .Y(n_707) );
OR2x2_ASAP7_75t_L g708 ( .A(n_705), .B(n_687), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_703), .A2(n_682), .B1(n_696), .B2(n_700), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_707), .A2(n_706), .B(n_682), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_708), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_709), .B1(n_704), .B2(n_700), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_710), .B(n_694), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_689), .B1(n_690), .B2(n_692), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_712), .B(n_699), .Y(n_715) );
endmodule