module real_aes_8035_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_0), .A2(n_100), .B1(n_109), .B2(n_744), .Y(n_99) );
NAND3xp33_ASAP7_75t_SL g102 ( .A(n_1), .B(n_103), .C(n_104), .Y(n_102) );
INVx1_ASAP7_75t_L g445 ( .A(n_1), .Y(n_445) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_2), .A2(n_138), .B(n_141), .C(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_3), .A2(n_166), .B(n_167), .Y(n_165) );
INVx1_ASAP7_75t_L g495 ( .A(n_4), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_5), .B(n_177), .Y(n_176) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_6), .A2(n_166), .B(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_L g138 ( .A(n_7), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g241 ( .A(n_8), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_9), .B(n_41), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_10), .A2(n_265), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_11), .B(n_150), .Y(n_218) );
INVx1_ASAP7_75t_L g477 ( .A(n_12), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_13), .B(n_171), .Y(n_528) );
INVx1_ASAP7_75t_L g130 ( .A(n_14), .Y(n_130) );
INVx1_ASAP7_75t_L g540 ( .A(n_15), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g225 ( .A1(n_16), .A2(n_185), .B(n_226), .C(n_228), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_17), .B(n_177), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_18), .B(n_466), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_19), .B(n_166), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_20), .B(n_273), .Y(n_272) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_21), .A2(n_171), .B(n_202), .C(n_205), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_22), .B(n_177), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_23), .B(n_150), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_24), .A2(n_204), .B(n_228), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_25), .B(n_150), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g132 ( .A(n_26), .Y(n_132) );
INVx1_ASAP7_75t_L g183 ( .A(n_27), .Y(n_183) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_28), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_29), .Y(n_214) );
AOI222xp33_ASAP7_75t_L g448 ( .A1(n_30), .A2(n_44), .B1(n_449), .B2(n_736), .C1(n_737), .C2(n_740), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_31), .B(n_150), .Y(n_496) );
INVx1_ASAP7_75t_L g270 ( .A(n_32), .Y(n_270) );
INVx1_ASAP7_75t_L g485 ( .A(n_33), .Y(n_485) );
INVx2_ASAP7_75t_L g136 ( .A(n_34), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_35), .Y(n_220) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_36), .A2(n_171), .B(n_172), .C(n_174), .Y(n_170) );
INVxp67_ASAP7_75t_L g271 ( .A(n_37), .Y(n_271) );
CKINVDCx14_ASAP7_75t_R g168 ( .A(n_38), .Y(n_168) );
A2O1A1Ixp33_ASAP7_75t_L g181 ( .A1(n_39), .A2(n_141), .B(n_182), .C(n_189), .Y(n_181) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_40), .A2(n_138), .B(n_141), .C(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g484 ( .A(n_42), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_43), .A2(n_116), .B1(n_437), .B2(n_438), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_43), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_44), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_45), .A2(n_152), .B(n_239), .C(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_46), .B(n_150), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_47), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_48), .Y(n_267) );
INVx1_ASAP7_75t_L g200 ( .A(n_49), .Y(n_200) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_50), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_51), .B(n_166), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_52), .A2(n_141), .B1(n_205), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_53), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_54), .Y(n_492) );
CKINVDCx14_ASAP7_75t_R g237 ( .A(n_55), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_56), .A2(n_174), .B(n_239), .C(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_57), .Y(n_520) );
INVx1_ASAP7_75t_L g474 ( .A(n_58), .Y(n_474) );
INVx1_ASAP7_75t_L g139 ( .A(n_59), .Y(n_139) );
INVx1_ASAP7_75t_L g129 ( .A(n_60), .Y(n_129) );
INVx1_ASAP7_75t_SL g173 ( .A(n_61), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_62), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_63), .B(n_177), .Y(n_207) );
INVx1_ASAP7_75t_L g145 ( .A(n_64), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_65), .A2(n_174), .B(n_466), .C(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_L g468 ( .A(n_66), .Y(n_468) );
INVx1_ASAP7_75t_L g106 ( .A(n_67), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_68), .A2(n_166), .B(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_69), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_70), .A2(n_166), .B(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_71), .Y(n_488) );
INVx1_ASAP7_75t_L g514 ( .A(n_72), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_73), .B(n_441), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_74), .A2(n_265), .B(n_266), .Y(n_264) );
CKINVDCx16_ASAP7_75t_R g180 ( .A(n_75), .Y(n_180) );
INVx1_ASAP7_75t_L g224 ( .A(n_76), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_77), .A2(n_138), .B(n_141), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_78), .A2(n_166), .B(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g227 ( .A(n_79), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_80), .B(n_184), .Y(n_508) );
INVx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
INVx1_ASAP7_75t_L g217 ( .A(n_82), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_83), .B(n_466), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_84), .A2(n_138), .B(n_141), .C(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g103 ( .A(n_85), .Y(n_103) );
OR2x2_ASAP7_75t_L g442 ( .A(n_85), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g735 ( .A(n_85), .B(n_444), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g140 ( .A1(n_86), .A2(n_141), .B(n_144), .C(n_154), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_87), .B(n_159), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_88), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_89), .A2(n_138), .B(n_141), .C(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_90), .Y(n_532) );
INVx1_ASAP7_75t_L g464 ( .A(n_91), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_92), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_93), .B(n_184), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_94), .B(n_125), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_95), .B(n_125), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_96), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g203 ( .A(n_97), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_98), .A2(n_166), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_101), .Y(n_746) );
OR2x2_ASAP7_75t_SL g101 ( .A(n_102), .B(n_107), .Y(n_101) );
OR2x2_ASAP7_75t_L g452 ( .A(n_103), .B(n_444), .Y(n_452) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_103), .B(n_443), .Y(n_739) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVxp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AND2x2_ASAP7_75t_L g444 ( .A(n_108), .B(n_445), .Y(n_444) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_114), .B(n_447), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx3_ASAP7_75t_L g743 ( .A(n_111), .Y(n_743) );
INVx2_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OAI21xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_439), .B(n_446), .Y(n_114) );
INVx3_ASAP7_75t_L g438 ( .A(n_116), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_116), .A2(n_451), .B1(n_734), .B2(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_SL g116 ( .A(n_117), .B(n_392), .Y(n_116) );
NOR4xp25_ASAP7_75t_L g117 ( .A(n_118), .B(n_329), .C(n_363), .D(n_379), .Y(n_117) );
NAND4xp25_ASAP7_75t_SL g118 ( .A(n_119), .B(n_255), .C(n_293), .D(n_309), .Y(n_118) );
AOI222xp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_192), .B1(n_230), .B2(n_243), .C1(n_248), .C2(n_254), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI31xp33_ASAP7_75t_L g425 ( .A1(n_121), .A2(n_426), .A3(n_427), .B(n_429), .Y(n_425) );
OR2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_160), .Y(n_121) );
AND2x2_ASAP7_75t_L g400 ( .A(n_122), .B(n_162), .Y(n_400) );
BUFx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_SL g247 ( .A(n_123), .Y(n_247) );
AND2x2_ASAP7_75t_L g254 ( .A(n_123), .B(n_178), .Y(n_254) );
AND2x2_ASAP7_75t_L g314 ( .A(n_123), .B(n_163), .Y(n_314) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_131), .B(n_156), .Y(n_123) );
INVx3_ASAP7_75t_L g177 ( .A(n_124), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_124), .B(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_124), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_124), .B(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_125), .Y(n_164) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_125), .A2(n_462), .B(n_469), .Y(n_461) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g263 ( .A(n_126), .Y(n_263) );
AND2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_127), .B(n_128), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B(n_140), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_133), .A2(n_159), .B(n_180), .C(n_181), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g213 ( .A1(n_133), .A2(n_214), .B(n_215), .Y(n_213) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_133), .A2(n_155), .B1(n_482), .B2(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_492), .B(n_493), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_133), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
AND2x4_ASAP7_75t_L g166 ( .A(n_134), .B(n_138), .Y(n_166) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g188 ( .A(n_135), .Y(n_188) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx1_ASAP7_75t_L g206 ( .A(n_136), .Y(n_206) );
INVx1_ASAP7_75t_L g143 ( .A(n_137), .Y(n_143) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_137), .Y(n_150) );
INVx3_ASAP7_75t_L g185 ( .A(n_137), .Y(n_185) );
INVx1_ASAP7_75t_L g466 ( .A(n_137), .Y(n_466) );
INVx4_ASAP7_75t_SL g155 ( .A(n_138), .Y(n_155) );
BUFx3_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
INVx5_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx3_ASAP7_75t_L g153 ( .A(n_142), .Y(n_153) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_146), .B(n_149), .C(n_151), .Y(n_144) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_146), .A2(n_151), .B(n_217), .C(n_218), .Y(n_216) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_147), .A2(n_148), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx4_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
INVx4_ASAP7_75t_L g171 ( .A(n_150), .Y(n_171) );
INVx2_ASAP7_75t_L g239 ( .A(n_150), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_151), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_151), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g228 ( .A(n_153), .Y(n_228) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
O2A1O1Ixp33_ASAP7_75t_L g167 ( .A1(n_155), .A2(n_168), .B(n_169), .C(n_170), .Y(n_167) );
O2A1O1Ixp33_ASAP7_75t_SL g199 ( .A1(n_155), .A2(n_169), .B(n_200), .C(n_201), .Y(n_199) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_155), .A2(n_169), .B(n_224), .C(n_225), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_SL g236 ( .A1(n_155), .A2(n_169), .B(n_237), .C(n_238), .Y(n_236) );
O2A1O1Ixp33_ASAP7_75t_SL g266 ( .A1(n_155), .A2(n_169), .B(n_267), .C(n_268), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_155), .A2(n_169), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_155), .A2(n_169), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_155), .A2(n_169), .B(n_537), .C(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
INVx1_ASAP7_75t_L g273 ( .A(n_158), .Y(n_273) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_158), .A2(n_524), .B(n_531), .Y(n_523) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx1_ASAP7_75t_L g212 ( .A(n_159), .Y(n_212) );
OA21x2_ASAP7_75t_L g234 ( .A1(n_159), .A2(n_235), .B(n_242), .Y(n_234) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_159), .A2(n_535), .B(n_541), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_160), .B(n_344), .Y(n_343) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_161), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_161), .B(n_258), .Y(n_304) );
AND2x2_ASAP7_75t_L g397 ( .A(n_161), .B(n_337), .Y(n_397) );
OAI321xp33_ASAP7_75t_L g431 ( .A1(n_161), .A2(n_247), .A3(n_404), .B1(n_432), .B2(n_434), .C(n_435), .Y(n_431) );
NAND4xp25_ASAP7_75t_L g435 ( .A(n_161), .B(n_233), .C(n_344), .D(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g161 ( .A(n_162), .B(n_178), .Y(n_161) );
AND2x2_ASAP7_75t_L g299 ( .A(n_162), .B(n_245), .Y(n_299) );
AND2x2_ASAP7_75t_L g318 ( .A(n_162), .B(n_247), .Y(n_318) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
AND2x2_ASAP7_75t_L g246 ( .A(n_163), .B(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g274 ( .A(n_163), .B(n_178), .Y(n_274) );
AND2x2_ASAP7_75t_L g360 ( .A(n_163), .B(n_245), .Y(n_360) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_176), .Y(n_163) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_164), .A2(n_198), .B(n_207), .Y(n_197) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_222), .B(n_229), .Y(n_221) );
BUFx2_ASAP7_75t_L g265 ( .A(n_166), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_171), .B(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_175), .Y(n_529) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_177), .A2(n_472), .B(n_478), .Y(n_471) );
INVx3_ASAP7_75t_SL g245 ( .A(n_178), .Y(n_245) );
AND2x2_ASAP7_75t_L g292 ( .A(n_178), .B(n_279), .Y(n_292) );
OR2x2_ASAP7_75t_L g325 ( .A(n_178), .B(n_247), .Y(n_325) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_178), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_178), .B(n_246), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_178), .B(n_334), .Y(n_376) );
AND2x2_ASAP7_75t_L g408 ( .A(n_178), .B(n_400), .Y(n_408) );
AND2x2_ASAP7_75t_L g417 ( .A(n_178), .B(n_259), .Y(n_417) );
OR2x6_ASAP7_75t_L g178 ( .A(n_179), .B(n_190), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_184), .A2(n_204), .B1(n_270), .B2(n_271), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_184), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_185), .B(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_185), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_185), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_188), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_208), .Y(n_193) );
INVx1_ASAP7_75t_SL g385 ( .A(n_194), .Y(n_385) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g250 ( .A(n_195), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g232 ( .A(n_196), .B(n_210), .Y(n_232) );
AND2x2_ASAP7_75t_L g321 ( .A(n_196), .B(n_234), .Y(n_321) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g291 ( .A(n_197), .B(n_221), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_197), .B(n_234), .Y(n_302) );
AND2x2_ASAP7_75t_L g328 ( .A(n_197), .B(n_234), .Y(n_328) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_197), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_204), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_204), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g497 ( .A(n_205), .Y(n_497) );
INVx3_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_208), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_208), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_SL g208 ( .A(n_209), .Y(n_208) );
OR2x2_ASAP7_75t_L g301 ( .A(n_209), .B(n_302), .Y(n_301) );
AOI322xp5_ASAP7_75t_L g387 ( .A1(n_209), .A2(n_291), .A3(n_297), .B1(n_328), .B2(n_378), .C1(n_388), .C2(n_390), .Y(n_387) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_210), .B(n_233), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_210), .B(n_234), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_210), .B(n_251), .Y(n_308) );
AND2x2_ASAP7_75t_L g362 ( .A(n_210), .B(n_328), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_210), .Y(n_366) );
AND2x2_ASAP7_75t_L g378 ( .A(n_210), .B(n_221), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_210), .B(n_250), .Y(n_410) );
INVx4_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g275 ( .A(n_211), .B(n_221), .Y(n_275) );
BUFx3_ASAP7_75t_L g289 ( .A(n_211), .Y(n_289) );
AND3x2_ASAP7_75t_L g371 ( .A(n_211), .B(n_351), .C(n_372), .Y(n_371) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_213), .B(n_219), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_212), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_212), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_212), .B(n_532), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g231 ( .A(n_221), .B(n_232), .C(n_233), .Y(n_231) );
INVx1_ASAP7_75t_SL g251 ( .A(n_221), .Y(n_251) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_221), .Y(n_356) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g350 ( .A(n_232), .B(n_351), .Y(n_350) );
INVxp67_ASAP7_75t_L g357 ( .A(n_232), .Y(n_357) );
AND2x2_ASAP7_75t_L g395 ( .A(n_233), .B(n_373), .Y(n_395) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
BUFx3_ASAP7_75t_L g276 ( .A(n_234), .Y(n_276) );
AND2x2_ASAP7_75t_L g351 ( .A(n_234), .B(n_251), .Y(n_351) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
OR2x2_ASAP7_75t_L g295 ( .A(n_245), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g414 ( .A(n_245), .B(n_314), .Y(n_414) );
AND2x2_ASAP7_75t_L g428 ( .A(n_245), .B(n_247), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_246), .B(n_259), .Y(n_369) );
AND2x2_ASAP7_75t_L g416 ( .A(n_246), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g279 ( .A(n_247), .B(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g296 ( .A(n_247), .B(n_259), .Y(n_296) );
INVx1_ASAP7_75t_L g306 ( .A(n_247), .Y(n_306) );
AND2x2_ASAP7_75t_L g337 ( .A(n_247), .B(n_259), .Y(n_337) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_249), .A2(n_380), .B1(n_384), .B2(n_386), .C(n_387), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_250), .B(n_252), .Y(n_249) );
AND2x2_ASAP7_75t_L g283 ( .A(n_250), .B(n_284), .Y(n_283) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_253), .B(n_290), .Y(n_433) );
AOI322xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_275), .A3(n_276), .B1(n_277), .B2(n_283), .C1(n_285), .C2(n_292), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_274), .Y(n_257) );
NAND2x1p5_ASAP7_75t_L g313 ( .A(n_258), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_258), .B(n_324), .Y(n_323) );
O2A1O1Ixp33_ASAP7_75t_L g347 ( .A1(n_258), .A2(n_274), .B(n_348), .C(n_349), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_258), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_258), .B(n_318), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_258), .B(n_400), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_258), .B(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_259), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_259), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g389 ( .A(n_259), .B(n_276), .Y(n_389) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_264), .B(n_272), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_261), .A2(n_281), .B(n_282), .Y(n_280) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_261), .A2(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AOI21xp5_ASAP7_75t_SL g504 ( .A1(n_262), .A2(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_263), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_263), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_263), .A2(n_491), .B(n_498), .Y(n_490) );
INVx1_ASAP7_75t_L g281 ( .A(n_264), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_272), .Y(n_282) );
INVx1_ASAP7_75t_L g364 ( .A(n_274), .Y(n_364) );
OAI31xp33_ASAP7_75t_L g374 ( .A1(n_274), .A2(n_299), .A3(n_375), .B(n_377), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_274), .B(n_280), .Y(n_426) );
INVx1_ASAP7_75t_SL g287 ( .A(n_275), .Y(n_287) );
AND2x2_ASAP7_75t_L g320 ( .A(n_275), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g401 ( .A(n_275), .B(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g286 ( .A(n_276), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g311 ( .A(n_276), .Y(n_311) );
AND2x2_ASAP7_75t_L g338 ( .A(n_276), .B(n_291), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_276), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g430 ( .A(n_276), .B(n_378), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_278), .B(n_348), .Y(n_421) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g317 ( .A(n_280), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g335 ( .A(n_280), .Y(n_335) );
NAND2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
OAI211xp5_ASAP7_75t_SL g329 ( .A1(n_287), .A2(n_330), .B(n_336), .C(n_352), .Y(n_329) );
OR2x2_ASAP7_75t_L g404 ( .A(n_287), .B(n_385), .Y(n_404) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
CKINVDCx16_ASAP7_75t_R g341 ( .A(n_289), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_289), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g310 ( .A(n_291), .B(n_311), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_297), .B(n_300), .C(n_303), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g344 ( .A(n_296), .Y(n_344) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_299), .B(n_337), .Y(n_342) );
INVx1_ASAP7_75t_L g348 ( .A(n_299), .Y(n_348) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g307 ( .A(n_302), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g340 ( .A(n_302), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g402 ( .A(n_302), .Y(n_402) );
AOI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_305), .B(n_307), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_305), .A2(n_316), .B(n_319), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B(n_315), .C(n_322), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_310), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_313), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g326 ( .A(n_314), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g381 ( .A1(n_316), .A2(n_382), .B(n_383), .Y(n_381) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_321), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g346 ( .A(n_321), .Y(n_346) );
AOI21xp33_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_326), .B(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g377 ( .A(n_328), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_334), .B(n_360), .Y(n_386) );
AND2x2_ASAP7_75t_L g399 ( .A(n_334), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g413 ( .A(n_334), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g423 ( .A(n_334), .B(n_361), .Y(n_423) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_339), .C(n_347), .Y(n_336) );
INVx1_ASAP7_75t_L g383 ( .A(n_337), .Y(n_383) );
OAI22xp33_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_342), .B1(n_343), .B2(n_345), .Y(n_339) );
OR2x2_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_341), .B(n_402), .Y(n_424) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g418 ( .A(n_351), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_358), .B1(n_361), .B2(n_362), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g436 ( .A(n_356), .Y(n_436) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g382 ( .A(n_360), .Y(n_382) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B(n_367), .C(n_374), .Y(n_363) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_382), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR5xp2_ASAP7_75t_L g392 ( .A(n_393), .B(n_411), .C(n_419), .D(n_425), .E(n_431), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_396), .B(n_398), .C(n_405), .Y(n_393) );
INVxp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AOI21xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B(n_403), .Y(n_398) );
OAI21xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_408), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_408), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_415), .B(n_418), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g434 ( .A(n_414), .Y(n_434) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_422), .B(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_438), .A2(n_451), .B1(n_453), .B2(n_734), .Y(n_450) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI21xp33_ASAP7_75t_L g447 ( .A1(n_446), .A2(n_448), .B(n_743), .Y(n_447) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g742 ( .A(n_453), .Y(n_742) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND4x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_652), .C(n_699), .D(n_719), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_582), .C(n_607), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_500), .B(n_542), .C(n_572), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_479), .Y(n_458) );
INVx3_ASAP7_75t_SL g624 ( .A(n_459), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_459), .B(n_555), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_459), .B(n_489), .Y(n_705) );
AND2x2_ASAP7_75t_L g728 ( .A(n_459), .B(n_594), .Y(n_728) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g546 ( .A(n_461), .B(n_471), .Y(n_546) );
INVx3_ASAP7_75t_L g559 ( .A(n_461), .Y(n_559) );
AND2x2_ASAP7_75t_L g564 ( .A(n_461), .B(n_470), .Y(n_564) );
OR2x2_ASAP7_75t_L g615 ( .A(n_461), .B(n_556), .Y(n_615) );
BUFx2_ASAP7_75t_L g635 ( .A(n_461), .Y(n_635) );
AND2x2_ASAP7_75t_L g645 ( .A(n_461), .B(n_556), .Y(n_645) );
AND2x2_ASAP7_75t_L g651 ( .A(n_461), .B(n_480), .Y(n_651) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_471), .B(n_556), .Y(n_570) );
INVx2_ASAP7_75t_L g580 ( .A(n_471), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_471), .B(n_559), .Y(n_593) );
OR2x2_ASAP7_75t_L g604 ( .A(n_471), .B(n_556), .Y(n_604) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_471), .B(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g662 ( .A(n_471), .Y(n_662) );
AND2x2_ASAP7_75t_L g708 ( .A(n_471), .B(n_480), .Y(n_708) );
INVx3_ASAP7_75t_SL g581 ( .A(n_479), .Y(n_581) );
OR2x2_ASAP7_75t_L g634 ( .A(n_479), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
INVx3_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
AND2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_490), .Y(n_623) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_480), .Y(n_691) );
AOI33xp33_ASAP7_75t_L g695 ( .A1(n_480), .A2(n_624), .A3(n_631), .B1(n_640), .B2(n_696), .B3(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g544 ( .A(n_489), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_489), .B(n_559), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_489), .B(n_619), .C(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g644 ( .A(n_489), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_489), .B(n_651), .Y(n_654) );
AND2x2_ASAP7_75t_L g707 ( .A(n_489), .B(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g563 ( .A(n_490), .Y(n_563) );
OR2x2_ASAP7_75t_L g657 ( .A(n_490), .B(n_556), .Y(n_657) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_521), .Y(n_500) );
AOI32xp33_ASAP7_75t_L g608 ( .A1(n_501), .A2(n_609), .A3(n_611), .B1(n_613), .B2(n_616), .Y(n_608) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_501), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g711 ( .A(n_501), .Y(n_711) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g643 ( .A(n_502), .B(n_627), .Y(n_643) );
AND2x2_ASAP7_75t_L g663 ( .A(n_502), .B(n_589), .Y(n_663) );
AND2x2_ASAP7_75t_L g731 ( .A(n_502), .B(n_649), .Y(n_731) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx3_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
AND2x2_ASAP7_75t_L g566 ( .A(n_503), .B(n_550), .Y(n_566) );
OR2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_549), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
AND2x2_ASAP7_75t_L g586 ( .A(n_503), .B(n_560), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_503), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_503), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g641 ( .A(n_503), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_503), .B(n_726), .Y(n_725) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
INVx2_ASAP7_75t_L g550 ( .A(n_512), .Y(n_550) );
AND2x2_ASAP7_75t_L g596 ( .A(n_512), .B(n_522), .Y(n_596) );
AND2x2_ASAP7_75t_L g606 ( .A(n_512), .B(n_534), .Y(n_606) );
INVx2_ASAP7_75t_L g726 ( .A(n_521), .Y(n_726) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_533), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_522), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g567 ( .A(n_522), .Y(n_567) );
AND2x2_ASAP7_75t_L g611 ( .A(n_522), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g627 ( .A(n_522), .B(n_590), .Y(n_627) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g640 ( .A(n_523), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_523), .B(n_550), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g551 ( .A(n_533), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_533), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g649 ( .A(n_533), .Y(n_649) );
INVx1_ASAP7_75t_L g682 ( .A(n_533), .Y(n_682) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g560 ( .A(n_534), .B(n_550), .Y(n_560) );
INVx1_ASAP7_75t_L g590 ( .A(n_534), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_547), .B1(n_553), .B2(n_560), .C(n_561), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_544), .B(n_564), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_544), .B(n_627), .Y(n_704) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_546), .B(n_594), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_546), .B(n_555), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_546), .B(n_569), .Y(n_698) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
AND2x2_ASAP7_75t_L g595 ( .A(n_551), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g673 ( .A(n_551), .Y(n_673) );
AND2x2_ASAP7_75t_L g605 ( .A(n_552), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_552), .B(n_575), .Y(n_621) );
AND2x2_ASAP7_75t_L g685 ( .A(n_552), .B(n_611), .Y(n_685) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g594 ( .A(n_556), .B(n_563), .Y(n_594) );
AND2x2_ASAP7_75t_L g690 ( .A(n_557), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_560), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_560), .B(n_567), .Y(n_655) );
AND2x2_ASAP7_75t_L g675 ( .A(n_560), .B(n_575), .Y(n_675) );
AND2x2_ASAP7_75t_L g696 ( .A(n_560), .B(n_640), .Y(n_696) );
OAI32xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .A3(n_567), .B1(n_568), .B2(n_571), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_SL g569 ( .A(n_563), .Y(n_569) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_563), .B(n_593), .Y(n_610) );
OR2x2_ASAP7_75t_L g614 ( .A(n_563), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_563), .B(n_662), .Y(n_715) );
INVx1_ASAP7_75t_L g583 ( .A(n_564), .Y(n_583) );
OAI221xp5_ASAP7_75t_SL g701 ( .A1(n_565), .A2(n_656), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g616 ( .A(n_566), .B(n_589), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_566), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g694 ( .A(n_566), .B(n_627), .Y(n_694) );
INVxp67_ASAP7_75t_L g630 ( .A(n_567), .Y(n_630) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g700 ( .A(n_569), .B(n_687), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_569), .B(n_650), .Y(n_723) );
INVx1_ASAP7_75t_L g598 ( .A(n_571), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_571), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g716 ( .A(n_571), .B(n_717), .Y(n_716) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_576), .B(n_579), .Y(n_572) );
AND2x2_ASAP7_75t_L g585 ( .A(n_574), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g669 ( .A(n_578), .B(n_589), .Y(n_669) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g687 ( .A(n_580), .B(n_645), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_580), .B(n_644), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_581), .B(n_593), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_587), .C(n_597), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_583), .A2(n_618), .B1(n_622), .B2(n_625), .C(n_628), .Y(n_617) );
AOI31xp33_ASAP7_75t_L g712 ( .A1(n_583), .A2(n_713), .A3(n_714), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .B1(n_593), .B2(n_595), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
INVx1_ASAP7_75t_L g676 ( .A(n_594), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_596), .A2(n_720), .B(n_722), .C(n_724), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_601), .B2(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_602), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g692 ( .A1(n_604), .A2(n_638), .B1(n_657), .B2(n_693), .C(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g688 ( .A(n_605), .Y(n_688) );
INVx1_ASAP7_75t_L g642 ( .A(n_606), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g607 ( .A(n_608), .B(n_617), .C(n_632), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_609), .A2(n_659), .B(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_611), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_639), .Y(n_656) );
INVx1_ASAP7_75t_L g631 ( .A(n_620), .Y(n_631) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g629 ( .A(n_623), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_623), .B(n_661), .Y(n_660) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_624), .B(n_629), .C(n_630), .D(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_643), .B2(n_644), .C1(n_646), .C2(n_650), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g730 ( .A(n_634), .Y(n_730) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_646), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_651), .A2(n_707), .B(n_709), .Y(n_706) );
NOR4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_664), .C(n_677), .D(n_692), .Y(n_652) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g733 ( .A(n_654), .Y(n_733) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_661), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
OAI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_670), .B2(n_671), .C1(n_674), .C2(n_676), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_669), .A2(n_700), .B(n_701), .C(n_712), .Y(n_699) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_683), .B1(n_684), .B2(n_686), .C1(n_688), .C2(n_689), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_694), .A2(n_697), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_727), .B(n_729), .C(n_732), .Y(n_724) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
endmodule