module real_aes_8403_n_383 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_383);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_383;
wire n_480;
wire n_1073;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_800;
wire n_778;
wire n_618;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_905;
wire n_1067;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1114;
wire n_580;
wire n_577;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_919;
wire n_857;
wire n_1089;
wire n_1122;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_571;
wire n_549;
wire n_694;
wire n_491;
wire n_1034;
wire n_894;
wire n_923;
wire n_1123;
wire n_952;
wire n_429;
wire n_1110;
wire n_1137;
wire n_448;
wire n_545;
wire n_556;
wire n_752;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_958;
wire n_677;
wire n_1021;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_678;
wire n_427;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_1072;
wire n_994;
wire n_1078;
wire n_384;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_824;
wire n_1098;
wire n_951;
wire n_467;
wire n_875;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_976;
wire n_466;
wire n_559;
wire n_1049;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_746;
wire n_532;
wire n_656;
wire n_1025;
wire n_1148;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_504;
wire n_725;
wire n_960;
wire n_671;
wire n_1081;
wire n_973;
wire n_1084;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1135;
wire n_641;
wire n_1063;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_1149;
wire n_405;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1131;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_1145;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_488;
wire n_1041;
wire n_501;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_1157;
wire n_471;
wire n_902;
wire n_1105;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_1136;
wire n_579;
wire n_1033;
wire n_533;
wire n_1000;
wire n_699;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_1127;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_831;
wire n_487;
wire n_653;
wire n_899;
wire n_526;
wire n_637;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_787;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_1130;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_1090;
wire n_456;
wire n_717;
wire n_982;
wire n_1133;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_546;
wire n_587;
wire n_1010;
wire n_811;
wire n_823;
wire n_459;
wire n_558;
wire n_1015;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1150;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1143;
wire n_929;
wire n_686;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_1045;
wire n_566;
wire n_719;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_1156;
wire n_829;
wire n_1030;
wire n_1088;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1151;
wire n_1036;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_968;
wire n_743;
wire n_710;
wire n_393;
wire n_1040;
wire n_703;
wire n_652;
wire n_500;
wire n_601;
wire n_1101;
wire n_661;
wire n_463;
wire n_1097;
wire n_396;
wire n_804;
wire n_1076;
wire n_447;
wire n_1102;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1144;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_0), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_1), .A2(n_166), .B1(n_470), .B2(n_474), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_2), .A2(n_171), .B1(n_561), .B2(n_769), .Y(n_807) );
INVx1_ASAP7_75t_L g816 ( .A(n_3), .Y(n_816) );
AOI22xp33_ASAP7_75t_SL g996 ( .A1(n_4), .A2(n_354), .B1(n_430), .B2(n_503), .Y(n_996) );
AOI22xp33_ASAP7_75t_SL g579 ( .A1(n_5), .A2(n_137), .B1(n_469), .B2(n_474), .Y(n_579) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_6), .A2(n_193), .B1(n_302), .B2(n_500), .C1(n_517), .C2(n_658), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_7), .A2(n_103), .B1(n_548), .B2(n_705), .Y(n_704) );
AO22x2_ASAP7_75t_L g417 ( .A1(n_8), .A2(n_227), .B1(n_408), .B2(n_413), .Y(n_417) );
INVx1_ASAP7_75t_L g1123 ( .A(n_8), .Y(n_1123) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_9), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_10), .A2(n_154), .B1(n_712), .B2(n_777), .Y(n_1057) );
AOI222xp33_ASAP7_75t_L g585 ( .A1(n_11), .A2(n_327), .B1(n_339), .B2(n_518), .C1(n_586), .C2(n_588), .Y(n_585) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_12), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_13), .Y(n_621) );
CKINVDCx20_ASAP7_75t_R g946 ( .A(n_14), .Y(n_946) );
INVx1_ASAP7_75t_L g1050 ( .A(n_15), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_16), .A2(n_56), .B1(n_773), .B2(n_831), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_17), .A2(n_132), .B1(n_571), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g885 ( .A1(n_18), .A2(n_121), .B1(n_554), .B2(n_886), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_19), .A2(n_201), .B1(n_446), .B2(n_664), .C(n_667), .Y(n_663) );
INVx1_ASAP7_75t_L g1039 ( .A(n_20), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g875 ( .A1(n_21), .A2(n_285), .B1(n_518), .B2(n_588), .Y(n_875) );
INVx1_ASAP7_75t_L g1043 ( .A(n_22), .Y(n_1043) );
INVx1_ASAP7_75t_L g744 ( .A(n_23), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_24), .A2(n_322), .B1(n_775), .B2(n_933), .Y(n_932) );
AOI22xp5_ASAP7_75t_SL g1071 ( .A1(n_25), .A2(n_196), .B1(n_769), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_SL g882 ( .A1(n_26), .A2(n_263), .B1(n_713), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_27), .A2(n_213), .B1(n_711), .B2(n_713), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g817 ( .A1(n_28), .A2(n_197), .B1(n_520), .B2(n_623), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g1089 ( .A1(n_29), .A2(n_112), .B1(n_429), .B2(n_506), .C(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_30), .A2(n_159), .B1(n_552), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_31), .A2(n_114), .B1(n_570), .B2(n_675), .Y(n_736) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_32), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_33), .A2(n_140), .B1(n_666), .B2(n_708), .Y(n_707) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_34), .A2(n_89), .B1(n_473), .B2(n_853), .Y(n_897) );
AO22x2_ASAP7_75t_L g415 ( .A1(n_35), .A2(n_120), .B1(n_408), .B2(n_409), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_36), .A2(n_254), .B1(n_474), .B2(n_853), .Y(n_959) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_37), .A2(n_273), .B1(n_512), .B2(n_712), .Y(n_993) );
AOI222xp33_ASAP7_75t_L g1065 ( .A1(n_38), .A2(n_195), .B1(n_301), .B2(n_473), .C1(n_520), .C2(n_653), .Y(n_1065) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_39), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_40), .B(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_41), .A2(n_318), .B1(n_800), .B2(n_974), .Y(n_973) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_42), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_43), .A2(n_261), .B1(n_552), .B2(n_553), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_44), .Y(n_724) );
AOI221xp5_ASAP7_75t_L g1098 ( .A1(n_45), .A2(n_208), .B1(n_821), .B2(n_899), .C(n_1099), .Y(n_1098) );
CKINVDCx20_ASAP7_75t_R g671 ( .A(n_46), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g1143 ( .A(n_47), .Y(n_1143) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_48), .A2(n_122), .B1(n_506), .B2(n_582), .Y(n_881) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_49), .A2(n_367), .B1(n_584), .B2(n_599), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_50), .A2(n_180), .B1(n_716), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_SL g1009 ( .A1(n_51), .A2(n_133), .B1(n_473), .B2(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_52), .A2(n_84), .B1(n_609), .B2(n_611), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_53), .B(n_697), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_54), .A2(n_101), .B1(n_512), .B2(n_514), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g931 ( .A(n_55), .Y(n_931) );
INVx1_ASAP7_75t_L g1032 ( .A(n_57), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_58), .A2(n_145), .B1(n_675), .B2(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g859 ( .A(n_59), .Y(n_859) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_60), .A2(n_91), .B1(n_711), .B2(n_769), .Y(n_768) );
AOI22x1_ASAP7_75t_L g1153 ( .A1(n_61), .A2(n_1127), .B1(n_1150), .B2(n_1154), .Y(n_1153) );
CKINVDCx20_ASAP7_75t_R g1154 ( .A(n_61), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_62), .A2(n_108), .B1(n_676), .B2(n_800), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g905 ( .A1(n_63), .A2(n_125), .B1(n_602), .B2(n_906), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g606 ( .A(n_64), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_65), .A2(n_281), .B1(n_446), .B2(n_846), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_66), .A2(n_233), .B1(n_512), .B2(n_741), .Y(n_829) );
AO22x1_ASAP7_75t_L g643 ( .A1(n_67), .A2(n_644), .B1(n_683), .B2(n_684), .Y(n_643) );
INVx1_ASAP7_75t_L g683 ( .A(n_67), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_68), .A2(n_181), .B1(n_351), .B2(n_478), .C1(n_479), .C2(n_483), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_69), .A2(n_98), .B1(n_573), .B2(n_574), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_70), .A2(n_317), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_71), .Y(n_617) );
INVx1_ASAP7_75t_L g1096 ( .A(n_72), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_73), .A2(n_369), .B1(n_573), .B2(n_611), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_74), .B(n_543), .Y(n_578) );
INVx1_ASAP7_75t_L g998 ( .A(n_75), .Y(n_998) );
AOI22xp33_ASAP7_75t_SL g715 ( .A1(n_76), .A2(n_381), .B1(n_429), .B2(n_716), .Y(n_715) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_77), .A2(n_167), .B1(n_708), .B2(n_1016), .Y(n_1015) );
AOI22xp33_ASAP7_75t_SL g997 ( .A1(n_78), .A2(n_232), .B1(n_514), .B2(n_800), .Y(n_997) );
AOI22xp33_ASAP7_75t_SL g1020 ( .A1(n_79), .A2(n_300), .B1(n_514), .B2(n_974), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_80), .A2(n_341), .B1(n_439), .B2(n_446), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g972 ( .A1(n_81), .A2(n_335), .B1(n_772), .B2(n_803), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_82), .A2(n_374), .B1(n_473), .B2(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g731 ( .A(n_83), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g938 ( .A(n_85), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_86), .A2(n_204), .B1(n_772), .B2(n_773), .Y(n_771) );
CKINVDCx20_ASAP7_75t_R g600 ( .A(n_87), .Y(n_600) );
AOI22xp33_ASAP7_75t_SL g994 ( .A1(n_88), .A2(n_259), .B1(n_506), .B2(n_827), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_90), .Y(n_790) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_92), .A2(n_110), .B1(n_740), .B2(n_775), .C(n_1094), .Y(n_1093) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_93), .Y(n_418) );
AO22x2_ASAP7_75t_L g412 ( .A1(n_94), .A2(n_260), .B1(n_408), .B2(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g1120 ( .A(n_94), .Y(n_1120) );
CKINVDCx20_ASAP7_75t_R g923 ( .A(n_95), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g1130 ( .A(n_96), .Y(n_1130) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_97), .A2(n_149), .B1(n_547), .B2(n_548), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_99), .A2(n_222), .B1(n_539), .B2(n_548), .Y(n_1079) );
CKINVDCx20_ASAP7_75t_R g1141 ( .A(n_100), .Y(n_1141) );
AOI22xp33_ASAP7_75t_SL g990 ( .A1(n_102), .A2(n_274), .B1(n_470), .B2(n_623), .Y(n_990) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_104), .A2(n_397), .B1(n_487), .B2(n_488), .Y(n_396) );
CKINVDCx16_ASAP7_75t_R g487 ( .A(n_104), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_105), .A2(n_116), .B1(n_184), .B2(n_517), .C1(n_518), .C2(n_521), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1061 ( .A1(n_106), .A2(n_371), .B1(n_469), .B2(n_500), .Y(n_1061) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_107), .Y(n_1007) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_109), .A2(n_954), .B1(n_975), .B2(n_976), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g975 ( .A(n_109), .Y(n_975) );
INVx1_ASAP7_75t_L g1100 ( .A(n_111), .Y(n_1100) );
XOR2x2_ASAP7_75t_L g530 ( .A(n_113), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g1081 ( .A(n_115), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_117), .A2(n_279), .B1(n_434), .B2(n_582), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g985 ( .A(n_118), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_119), .A2(n_270), .B1(n_404), .B2(n_503), .Y(n_1070) );
INVx1_ASAP7_75t_L g1124 ( .A(n_120), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_123), .A2(n_265), .B1(n_1075), .B2(n_1133), .Y(n_1132) );
AOI22xp5_ASAP7_75t_L g1074 ( .A1(n_124), .A2(n_306), .B1(n_429), .B2(n_1075), .Y(n_1074) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_126), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g1144 ( .A(n_127), .Y(n_1144) );
XOR2x2_ASAP7_75t_L g869 ( .A(n_128), .B(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_129), .B(n_545), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_130), .Y(n_647) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_131), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g1140 ( .A(n_134), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_135), .A2(n_151), .B1(n_451), .B2(n_454), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_136), .B(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_138), .A2(n_355), .B1(n_430), .B2(n_443), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g957 ( .A(n_139), .Y(n_957) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_141), .Y(n_1148) );
AOI22xp5_ASAP7_75t_L g1087 ( .A1(n_142), .A2(n_1088), .B1(n_1103), .B2(n_1104), .Y(n_1087) );
INVx1_ASAP7_75t_L g1103 ( .A(n_142), .Y(n_1103) );
OAI22xp5_ASAP7_75t_SL g749 ( .A1(n_143), .A2(n_750), .B1(n_751), .B2(n_778), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_143), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_144), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_146), .A2(n_165), .B1(n_772), .B2(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g1095 ( .A(n_147), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_148), .A2(n_231), .B1(n_802), .B2(n_803), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_150), .A2(n_362), .B1(n_446), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g759 ( .A(n_152), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_153), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_155), .A2(n_202), .B1(n_483), .B2(n_623), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_156), .A2(n_211), .B1(n_469), .B2(n_473), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_157), .A2(n_307), .B1(n_570), .B2(n_571), .Y(n_569) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_158), .A2(n_347), .B1(n_556), .B2(n_908), .Y(n_907) );
AND2x6_ASAP7_75t_L g386 ( .A(n_160), .B(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_160), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_161), .A2(n_284), .B1(n_561), .B2(n_565), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_162), .A2(n_334), .B1(n_500), .B2(n_520), .Y(n_729) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_163), .A2(n_266), .B1(n_694), .B2(n_697), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g949 ( .A(n_164), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_168), .A2(n_338), .B1(n_769), .B2(n_1035), .Y(n_1034) );
AOI222xp33_ASAP7_75t_L g865 ( .A1(n_169), .A2(n_244), .B1(n_258), .B2(n_478), .C1(n_500), .C2(n_697), .Y(n_865) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_170), .Y(n_589) );
INVx1_ASAP7_75t_L g866 ( .A(n_172), .Y(n_866) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_173), .A2(n_343), .B1(n_402), .B2(n_603), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_174), .Y(n_1135) );
AOI22xp33_ASAP7_75t_SL g826 ( .A1(n_175), .A2(n_363), .B1(n_451), .B2(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g682 ( .A(n_176), .Y(n_682) );
INVx1_ASAP7_75t_L g1049 ( .A(n_177), .Y(n_1049) );
AOI22xp5_ASAP7_75t_L g1076 ( .A1(n_178), .A2(n_321), .B1(n_603), .B2(n_664), .Y(n_1076) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_179), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_182), .A2(n_256), .B1(n_711), .B2(n_713), .Y(n_1137) );
AOI22xp5_ASAP7_75t_L g559 ( .A1(n_183), .A2(n_250), .B1(n_560), .B2(n_561), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_185), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_186), .A2(n_353), .B1(n_434), .B2(n_743), .Y(n_742) );
AO22x2_ASAP7_75t_L g407 ( .A1(n_187), .A2(n_251), .B1(n_408), .B2(n_409), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_187), .B(n_1122), .Y(n_1121) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_188), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_189), .A2(n_219), .B1(n_564), .B2(n_565), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g576 ( .A(n_190), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_191), .Y(n_894) );
INVx1_ASAP7_75t_L g692 ( .A(n_192), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g874 ( .A(n_194), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_198), .B(n_484), .Y(n_791) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_199), .Y(n_755) );
AOI22xp33_ASAP7_75t_SL g902 ( .A1(n_200), .A2(n_349), .B1(n_769), .B2(n_903), .Y(n_902) );
XOR2x2_ASAP7_75t_L g490 ( .A(n_203), .B(n_491), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_205), .A2(n_278), .B1(n_821), .B2(n_899), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_206), .A2(n_311), .B1(n_494), .B2(n_700), .Y(n_1078) );
CKINVDCx20_ASAP7_75t_R g1066 ( .A(n_207), .Y(n_1066) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_209), .Y(n_467) );
OA22x2_ASAP7_75t_L g1028 ( .A1(n_210), .A2(n_1029), .B1(n_1030), .B2(n_1052), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_210), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_212), .A2(n_298), .B1(n_675), .B2(n_676), .C(n_679), .Y(n_674) );
INVx1_ASAP7_75t_L g861 ( .A(n_214), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g969 ( .A(n_215), .Y(n_969) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_216), .A2(n_305), .B1(n_494), .B2(n_497), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g988 ( .A(n_217), .B(n_494), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_218), .B(n_483), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_220), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g1145 ( .A(n_221), .Y(n_1145) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_223), .A2(n_269), .B1(n_430), .B2(n_451), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_224), .B(n_700), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_225), .A2(n_296), .B1(n_506), .B2(n_508), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_226), .A2(n_247), .B1(n_484), .B2(n_705), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_228), .A2(n_320), .B1(n_474), .B2(n_1046), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_229), .A2(n_283), .B1(n_666), .B2(n_827), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_230), .A2(n_299), .B1(n_521), .B2(n_853), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_234), .A2(n_370), .B1(n_454), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g1131 ( .A(n_235), .Y(n_1131) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_236), .Y(n_427) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_237), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g1005 ( .A(n_238), .Y(n_1005) );
CKINVDCx20_ASAP7_75t_R g632 ( .A(n_239), .Y(n_632) );
INVx1_ASAP7_75t_L g857 ( .A(n_240), .Y(n_857) );
INVx1_ASAP7_75t_L g1101 ( .A(n_241), .Y(n_1101) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_242), .A2(n_337), .B1(n_469), .B2(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_243), .A2(n_264), .B1(n_451), .B2(n_454), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_245), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_246), .A2(n_380), .B1(n_899), .B2(n_1012), .Y(n_1011) );
INVx2_ASAP7_75t_L g391 ( .A(n_248), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_249), .A2(n_280), .B1(n_484), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g962 ( .A(n_252), .Y(n_962) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_253), .Y(n_925) );
XNOR2xp5_ASAP7_75t_L g999 ( .A(n_255), .B(n_1000), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_257), .A2(n_303), .B1(n_479), .B2(n_520), .Y(n_1082) );
AOI211xp5_ASAP7_75t_L g383 ( .A1(n_262), .A2(n_384), .B(n_392), .C(n_1125), .Y(n_383) );
INVx1_ASAP7_75t_L g733 ( .A(n_267), .Y(n_733) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_268), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_271), .A2(n_291), .B1(n_602), .B2(n_603), .Y(n_601) );
CKINVDCx20_ASAP7_75t_R g963 ( .A(n_272), .Y(n_963) );
INVx1_ASAP7_75t_L g1033 ( .A(n_275), .Y(n_1033) );
AOI22xp33_ASAP7_75t_SL g887 ( .A1(n_276), .A2(n_378), .B1(n_777), .B2(n_802), .Y(n_887) );
XOR2x2_ASAP7_75t_L g687 ( .A(n_277), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g408 ( .A(n_282), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_282), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g968 ( .A(n_286), .Y(n_968) );
CKINVDCx20_ASAP7_75t_R g958 ( .A(n_287), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_288), .A2(n_368), .B1(n_711), .B2(n_713), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_289), .B(n_543), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_290), .A2(n_345), .B1(n_553), .B2(n_886), .Y(n_1041) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_292), .Y(n_786) );
INVx1_ASAP7_75t_L g1092 ( .A(n_293), .Y(n_1092) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_294), .B(n_497), .Y(n_819) );
INVx1_ASAP7_75t_L g1051 ( .A(n_295), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g918 ( .A1(n_297), .A2(n_919), .B1(n_950), .B2(n_951), .Y(n_918) );
INVx1_ASAP7_75t_L g950 ( .A(n_297), .Y(n_950) );
CKINVDCx20_ASAP7_75t_R g1003 ( .A(n_304), .Y(n_1003) );
CKINVDCx20_ASAP7_75t_R g936 ( .A(n_308), .Y(n_936) );
INVx1_ASAP7_75t_L g1044 ( .A(n_309), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_310), .Y(n_793) );
AOI22xp5_ASAP7_75t_L g1126 ( .A1(n_312), .A2(n_1127), .B1(n_1149), .B2(n_1150), .Y(n_1126) );
CKINVDCx20_ASAP7_75t_R g1149 ( .A(n_312), .Y(n_1149) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_313), .Y(n_432) );
INVx1_ASAP7_75t_L g680 ( .A(n_314), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_315), .B(n_821), .Y(n_820) );
OA22x2_ASAP7_75t_L g889 ( .A1(n_316), .A2(n_890), .B1(n_891), .B2(n_910), .Y(n_889) );
CKINVDCx20_ASAP7_75t_R g890 ( .A(n_316), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_319), .A2(n_376), .B1(n_498), .B2(n_543), .Y(n_1060) );
INVx1_ASAP7_75t_L g390 ( .A(n_323), .Y(n_390) );
CKINVDCx20_ASAP7_75t_R g929 ( .A(n_324), .Y(n_929) );
CKINVDCx20_ASAP7_75t_R g789 ( .A(n_325), .Y(n_789) );
INVx1_ASAP7_75t_L g387 ( .A(n_326), .Y(n_387) );
INVx1_ASAP7_75t_L g1083 ( .A(n_328), .Y(n_1083) );
CKINVDCx20_ASAP7_75t_R g1147 ( .A(n_329), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_330), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_331), .A2(n_336), .B1(n_503), .B2(n_800), .Y(n_1063) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_332), .Y(n_728) );
INVx1_ASAP7_75t_L g863 ( .A(n_333), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_340), .Y(n_795) );
INVx1_ASAP7_75t_L g1091 ( .A(n_342), .Y(n_1091) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_344), .A2(n_364), .B1(n_561), .B2(n_1018), .Y(n_1017) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_346), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g965 ( .A(n_348), .Y(n_965) );
CKINVDCx20_ASAP7_75t_R g1136 ( .A(n_350), .Y(n_1136) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_352), .Y(n_614) );
INVx1_ASAP7_75t_L g849 ( .A(n_356), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g948 ( .A(n_357), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_358), .B(n_497), .Y(n_989) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_359), .B(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_360), .A2(n_373), .B1(n_678), .B2(n_743), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_361), .B(n_700), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_365), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_366), .B(n_851), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_372), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g781 ( .A1(n_375), .A2(n_782), .B1(n_808), .B2(n_809), .Y(n_781) );
INVx1_ASAP7_75t_L g808 ( .A(n_375), .Y(n_808) );
INVx1_ASAP7_75t_L g1040 ( .A(n_377), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_379), .A2(n_593), .B1(n_638), .B2(n_639), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_379), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g726 ( .A(n_382), .Y(n_726) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_386), .B(n_388), .Y(n_385) );
HB1xp67_ASAP7_75t_L g1116 ( .A(n_387), .Y(n_1116) );
OA21x2_ASAP7_75t_L g1156 ( .A1(n_388), .A2(n_1115), .B(n_1157), .Y(n_1156) );
NOR2xp33_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_838), .B1(n_1110), .B2(n_1111), .C(n_1112), .Y(n_392) );
INVx1_ASAP7_75t_L g1110 ( .A(n_393), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_524), .B1(n_836), .B2(n_837), .Y(n_393) );
INVx1_ASAP7_75t_L g836 ( .A(n_394), .Y(n_836) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_489), .B1(n_522), .B2(n_523), .Y(n_395) );
INVx1_ASAP7_75t_L g522 ( .A(n_396), .Y(n_522) );
INVx2_ASAP7_75t_SL g488 ( .A(n_397), .Y(n_488) );
AND4x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_437), .C(n_457), .D(n_477), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_399), .B(n_426), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_418), .B2(n_419), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_401), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_401), .A2(n_513), .B1(n_1039), .B2(n_1040), .C(n_1041), .Y(n_1038) );
OAI221xp5_ASAP7_75t_SL g1134 ( .A1(n_401), .A2(n_419), .B1(n_1135), .B2(n_1136), .C(n_1137), .Y(n_1134) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g560 ( .A(n_403), .Y(n_560) );
INVx3_ASAP7_75t_L g741 ( .A(n_403), .Y(n_741) );
INVx2_ASAP7_75t_L g803 ( .A(n_403), .Y(n_803) );
INVx6_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g514 ( .A(n_404), .Y(n_514) );
BUFx3_ASAP7_75t_L g584 ( .A(n_404), .Y(n_584) );
BUFx3_ASAP7_75t_L g777 ( .A(n_404), .Y(n_777) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_414), .Y(n_404) );
AND2x2_ASAP7_75t_L g431 ( .A(n_405), .B(n_424), .Y(n_431) );
AND2x6_ASAP7_75t_L g443 ( .A(n_405), .B(n_444), .Y(n_443) );
AND2x6_ASAP7_75t_L g478 ( .A(n_405), .B(n_476), .Y(n_478) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_411), .Y(n_405) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_412), .Y(n_436) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g422 ( .A(n_407), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_407), .B(n_412), .Y(n_449) );
AND2x2_ASAP7_75t_L g472 ( .A(n_407), .B(n_417), .Y(n_472) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_410), .Y(n_413) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g423 ( .A(n_412), .Y(n_423) );
INVx1_ASAP7_75t_L g482 ( .A(n_412), .Y(n_482) );
AND2x2_ASAP7_75t_L g453 ( .A(n_414), .B(n_422), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g466 ( .A(n_414), .B(n_436), .Y(n_466) );
AND2x6_ASAP7_75t_L g498 ( .A(n_414), .B(n_436), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_414), .B(n_422), .Y(n_670) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx2_ASAP7_75t_L g425 ( .A(n_415), .Y(n_425) );
OR2x2_ASAP7_75t_L g445 ( .A(n_415), .B(n_416), .Y(n_445) );
INVx1_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AND2x2_ASAP7_75t_L g476 ( .A(n_415), .B(n_417), .Y(n_476) );
AND2x2_ASAP7_75t_L g424 ( .A(n_416), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI221xp5_ASAP7_75t_SL g604 ( .A1(n_419), .A2(n_605), .B1(n_606), .B2(n_607), .C(n_608), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_419), .A2(n_857), .B1(n_858), .B2(n_859), .Y(n_856) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g922 ( .A(n_420), .Y(n_922) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_422), .B(n_424), .Y(n_421) );
AND2x2_ASAP7_75t_L g504 ( .A(n_422), .B(n_424), .Y(n_504) );
INVx1_ASAP7_75t_L g475 ( .A(n_423), .Y(n_475) );
AND2x4_ASAP7_75t_L g435 ( .A(n_424), .B(n_436), .Y(n_435) );
AND2x4_ASAP7_75t_L g447 ( .A(n_424), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g481 ( .A(n_425), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g631 ( .A(n_425), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_432), .B2(n_433), .Y(n_426) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g596 ( .A(n_430), .Y(n_596) );
BUFx3_ASAP7_75t_L g772 ( .A(n_430), .Y(n_772) );
BUFx3_ASAP7_75t_L g933 ( .A(n_430), .Y(n_933) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g557 ( .A(n_431), .Y(n_557) );
BUFx2_ASAP7_75t_SL g582 ( .A(n_431), .Y(n_582) );
BUFx2_ASAP7_75t_SL g675 ( .A(n_431), .Y(n_675) );
INVxp67_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g599 ( .A(n_434), .Y(n_599) );
BUFx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g507 ( .A(n_435), .Y(n_507) );
BUFx3_ASAP7_75t_L g564 ( .A(n_435), .Y(n_564) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_435), .Y(n_666) );
BUFx3_ASAP7_75t_L g773 ( .A(n_435), .Y(n_773) );
INVx1_ASAP7_75t_L g461 ( .A(n_436), .Y(n_461) );
AND2x4_ASAP7_75t_L g496 ( .A(n_436), .B(n_444), .Y(n_496) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_450), .Y(n_437) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx5_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g552 ( .A(n_442), .Y(n_552) );
INVx4_ASAP7_75t_L g740 ( .A(n_442), .Y(n_740) );
INVx2_ASAP7_75t_L g1075 ( .A(n_442), .Y(n_1075) );
INVx11_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx11_ASAP7_75t_L g513 ( .A(n_443), .Y(n_513) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g460 ( .A(n_445), .B(n_461), .Y(n_460) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
BUFx3_ASAP7_75t_L g571 ( .A(n_447), .Y(n_571) );
BUFx2_ASAP7_75t_SL g603 ( .A(n_447), .Y(n_603) );
BUFx2_ASAP7_75t_L g743 ( .A(n_447), .Y(n_743) );
BUFx3_ASAP7_75t_L g800 ( .A(n_447), .Y(n_800) );
BUFx2_ASAP7_75t_SL g886 ( .A(n_447), .Y(n_886) );
BUFx3_ASAP7_75t_L g909 ( .A(n_447), .Y(n_909) );
AND2x2_ASAP7_75t_L g827 ( .A(n_448), .B(n_631), .Y(n_827) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g455 ( .A(n_449), .B(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_451), .Y(n_903) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g562 ( .A(n_452), .Y(n_562) );
INVx3_ASAP7_75t_L g573 ( .A(n_452), .Y(n_573) );
INVx1_ASAP7_75t_L g610 ( .A(n_452), .Y(n_610) );
INVx5_ASAP7_75t_L g712 ( .A(n_452), .Y(n_712) );
INVx4_ASAP7_75t_L g1037 ( .A(n_452), .Y(n_1037) );
INVx8_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g565 ( .A(n_454), .Y(n_565) );
BUFx2_ASAP7_75t_L g574 ( .A(n_454), .Y(n_574) );
BUFx4f_ASAP7_75t_SL g673 ( .A(n_454), .Y(n_673) );
BUFx2_ASAP7_75t_L g713 ( .A(n_454), .Y(n_713) );
BUFx2_ASAP7_75t_L g769 ( .A(n_454), .Y(n_769) );
INVx6_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g611 ( .A(n_455), .Y(n_611) );
INVx1_ASAP7_75t_SL g1018 ( .A(n_455), .Y(n_1018) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_455), .A2(n_669), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
INVx1_ASAP7_75t_L g471 ( .A(n_456), .Y(n_471) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
OAI221xp5_ASAP7_75t_SL g458 ( .A1(n_459), .A2(n_462), .B1(n_463), .B2(n_467), .C(n_468), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g784 ( .A1(n_459), .A2(n_650), .B1(n_785), .B2(n_786), .Y(n_784) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g616 ( .A(n_460), .Y(n_616) );
BUFx3_ASAP7_75t_L g725 ( .A(n_460), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g753 ( .A1(n_463), .A2(n_648), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx3_ASAP7_75t_L g577 ( .A(n_465), .Y(n_577) );
BUFx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g619 ( .A(n_466), .Y(n_619) );
BUFx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g548 ( .A(n_470), .Y(n_548) );
INVx1_ASAP7_75t_L g854 ( .A(n_470), .Y(n_854) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_470), .Y(n_1010) );
AND2x4_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
AND2x4_ASAP7_75t_L g480 ( .A(n_472), .B(n_481), .Y(n_480) );
AND2x4_ASAP7_75t_L g485 ( .A(n_472), .B(n_486), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g630 ( .A(n_472), .B(n_631), .Y(n_630) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_SL g521 ( .A(n_474), .Y(n_521) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
BUFx2_ASAP7_75t_SL g705 ( .A(n_474), .Y(n_705) );
AND2x4_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g637 ( .A(n_475), .Y(n_637) );
INVx1_ASAP7_75t_L g636 ( .A(n_476), .Y(n_636) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_478), .Y(n_517) );
INVx2_ASAP7_75t_SL g534 ( .A(n_478), .Y(n_534) );
INVx4_ASAP7_75t_L g587 ( .A(n_478), .Y(n_587) );
BUFx3_ASAP7_75t_L g653 ( .A(n_478), .Y(n_653) );
INVx2_ASAP7_75t_L g984 ( .A(n_478), .Y(n_984) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_480), .Y(n_500) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_480), .Y(n_547) );
BUFx4f_ASAP7_75t_SL g623 ( .A(n_480), .Y(n_623) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_480), .Y(n_696) );
INVx1_ASAP7_75t_L g486 ( .A(n_482), .Y(n_486) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx3_ASAP7_75t_L g945 ( .A(n_484), .Y(n_945) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx12f_ASAP7_75t_L g520 ( .A(n_485), .Y(n_520) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_485), .Y(n_697) );
INVx1_ASAP7_75t_L g1006 ( .A(n_485), .Y(n_1006) );
INVxp67_ASAP7_75t_L g523 ( .A(n_489), .Y(n_523) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND4xp75_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .C(n_510), .D(n_516), .Y(n_491) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_493), .B(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx5_ASAP7_75t_L g543 ( .A(n_495), .Y(n_543) );
INVx2_ASAP7_75t_L g703 ( .A(n_495), .Y(n_703) );
INVx2_ASAP7_75t_L g821 ( .A(n_495), .Y(n_821) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx4f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g545 ( .A(n_498), .Y(n_545) );
INVx1_ASAP7_75t_SL g701 ( .A(n_498), .Y(n_701) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_500), .Y(n_588) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_505), .Y(n_501) );
INVx1_ASAP7_75t_L g717 ( .A(n_503), .Y(n_717) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx3_ASAP7_75t_L g554 ( .A(n_504), .Y(n_554) );
BUFx3_ASAP7_75t_L g570 ( .A(n_504), .Y(n_570) );
BUFx3_ASAP7_75t_L g678 ( .A(n_504), .Y(n_678) );
INVx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_515), .Y(n_510) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g602 ( .A(n_513), .Y(n_602) );
INVx3_ASAP7_75t_L g767 ( .A(n_513), .Y(n_767) );
INVx2_ASAP7_75t_SL g802 ( .A(n_513), .Y(n_802) );
INVx2_ASAP7_75t_SL g873 ( .A(n_517), .Y(n_873) );
INVx2_ASAP7_75t_L g942 ( .A(n_517), .Y(n_942) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx4f_ASAP7_75t_SL g658 ( .A(n_520), .Y(n_658) );
INVx1_ASAP7_75t_L g837 ( .A(n_524), .Y(n_837) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_526), .B1(n_746), .B2(n_835), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B1(n_640), .B2(n_641), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
XNOR2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_592), .Y(n_528) );
AO22x2_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_566), .B1(n_590), .B2(n_591), .Y(n_529) );
INVx2_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_532), .B(n_549), .Y(n_531) );
NOR2xp33_ASAP7_75t_SL g532 ( .A(n_533), .B(n_540), .Y(n_532) );
OAI21xp5_ASAP7_75t_SL g533 ( .A1(n_534), .A2(n_535), .B(n_536), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_534), .A2(n_621), .B1(n_622), .B2(n_624), .C(n_625), .Y(n_620) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .C(n_546), .Y(n_540) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx6f_ASAP7_75t_L g1012 ( .A(n_543), .Y(n_1012) );
CKINVDCx20_ASAP7_75t_R g961 ( .A(n_547), .Y(n_961) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_555), .Y(n_550) );
INVx1_ASAP7_75t_L g709 ( .A(n_552), .Y(n_709) );
BUFx4f_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx3_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx3_ASAP7_75t_L g831 ( .A(n_557), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
INVx3_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_564), .Y(n_806) );
INVx3_ASAP7_75t_SL g591 ( .A(n_566), .Y(n_591) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_589), .Y(n_566) );
NAND4xp75_ASAP7_75t_L g567 ( .A(n_568), .B(n_575), .C(n_580), .D(n_585), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
BUFx3_ASAP7_75t_L g906 ( .A(n_570), .Y(n_906) );
INVxp67_ASAP7_75t_L g858 ( .A(n_571), .Y(n_858) );
OA211x2_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_577), .B(n_578), .C(n_579), .Y(n_575) );
OA211x2_ASAP7_75t_L g848 ( .A1(n_577), .A2(n_849), .B(n_850), .C(n_852), .Y(n_848) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
INVx1_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
INVx2_ASAP7_75t_L g691 ( .A(n_586), .Y(n_691) );
INVx4_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
BUFx2_ASAP7_75t_L g788 ( .A(n_587), .Y(n_788) );
OAI222xp33_ASAP7_75t_L g1047 ( .A1(n_587), .A2(n_964), .B1(n_1048), .B2(n_1049), .C1(n_1050), .C2(n_1051), .Y(n_1047) );
INVx2_ASAP7_75t_SL g655 ( .A(n_588), .Y(n_655) );
INVx2_ASAP7_75t_SL g758 ( .A(n_588), .Y(n_758) );
INVx2_ASAP7_75t_L g639 ( .A(n_593), .Y(n_639) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_594), .B(n_612), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_604), .Y(n_594) );
OAI221xp5_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_597), .B1(n_598), .B2(n_600), .C(n_601), .Y(n_595) );
INVx2_ASAP7_75t_L g1016 ( .A(n_596), .Y(n_1016) );
OAI221xp5_ASAP7_75t_SL g1031 ( .A1(n_596), .A2(n_665), .B1(n_1032), .B2(n_1033), .C(n_1034), .Y(n_1031) );
OAI221xp5_ASAP7_75t_SL g1129 ( .A1(n_596), .A2(n_930), .B1(n_1130), .B2(n_1131), .C(n_1132), .Y(n_1129) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g681 ( .A(n_602), .Y(n_681) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR3xp33_ASAP7_75t_L g612 ( .A(n_613), .B(n_620), .C(n_626), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_617), .B2(n_618), .Y(n_613) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g648 ( .A(n_616), .Y(n_648) );
INVx2_ASAP7_75t_L g937 ( .A(n_616), .Y(n_937) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_618), .A2(n_724), .B1(n_725), .B2(n_726), .Y(n_723) );
OAI221xp5_ASAP7_75t_SL g956 ( .A1(n_618), .A2(n_937), .B1(n_957), .B2(n_958), .C(n_959), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g1042 ( .A1(n_618), .A2(n_937), .B1(n_1043), .B2(n_1044), .C(n_1045), .Y(n_1042) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_SL g650 ( .A(n_619), .Y(n_650) );
INVx2_ASAP7_75t_L g939 ( .A(n_619), .Y(n_939) );
OAI221xp5_ASAP7_75t_SL g787 ( .A1(n_622), .A2(n_788), .B1(n_789), .B2(n_790), .C(n_791), .Y(n_787) );
OAI222xp33_ASAP7_75t_L g1142 ( .A1(n_622), .A2(n_942), .B1(n_964), .B2(n_1143), .C1(n_1144), .C2(n_1145), .Y(n_1142) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_628), .B1(n_632), .B2(n_633), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_628), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_628), .A2(n_633), .B1(n_948), .B2(n_949), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_628), .A2(n_633), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx3_ASAP7_75t_SL g794 ( .A(n_629), .Y(n_794) );
INVx4_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
BUFx3_ASAP7_75t_L g732 ( .A(n_630), .Y(n_732) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_L g662 ( .A(n_634), .Y(n_662) );
CKINVDCx16_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_635), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
BUFx2_ASAP7_75t_L g796 ( .A(n_635), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_635), .A2(n_732), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
OR2x6_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_643), .B1(n_685), .B2(n_686), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g684 ( .A(n_644), .Y(n_684) );
AND3x1_ASAP7_75t_L g644 ( .A(n_645), .B(n_663), .C(n_674), .Y(n_644) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_651), .C(n_659), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_651) );
OAI21xp33_ASAP7_75t_L g727 ( .A1(n_652), .A2(n_728), .B(n_729), .Y(n_727) );
OAI21xp5_ASAP7_75t_SL g815 ( .A1(n_652), .A2(n_816), .B(n_817), .Y(n_815) );
OAI21xp5_ASAP7_75t_SL g893 ( .A1(n_652), .A2(n_894), .B(n_895), .Y(n_893) );
INVx3_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g964 ( .A(n_658), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_662), .A2(n_732), .B1(n_762), .B2(n_763), .Y(n_761) );
INVx4_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx3_ASAP7_75t_L g846 ( .A(n_665), .Y(n_846) );
OAI221xp5_ASAP7_75t_SL g967 ( .A1(n_665), .A2(n_928), .B1(n_968), .B2(n_969), .C(n_970), .Y(n_967) );
INVx4_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_667) );
BUFx2_ASAP7_75t_R g669 ( .A(n_670), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx2_ASAP7_75t_L g974 ( .A(n_678), .Y(n_974) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_719), .B1(n_720), .B2(n_745), .Y(n_686) );
INVx2_ASAP7_75t_L g745 ( .A(n_687), .Y(n_745) );
NAND3x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_706), .C(n_714), .Y(n_688) );
NOR2x1_ASAP7_75t_SL g689 ( .A(n_690), .B(n_698), .Y(n_689) );
OAI21xp5_ASAP7_75t_SL g690 ( .A1(n_691), .A2(n_692), .B(n_693), .Y(n_690) );
OAI221xp5_ASAP7_75t_SL g756 ( .A1(n_691), .A2(n_757), .B1(n_758), .B2(n_759), .C(n_760), .Y(n_756) );
OAI222xp33_ASAP7_75t_L g960 ( .A1(n_691), .A2(n_961), .B1(n_962), .B2(n_963), .C1(n_964), .C2(n_965), .Y(n_960) );
INVx1_ASAP7_75t_L g1048 ( .A(n_694), .Y(n_1048) );
INVx3_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx4_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g1004 ( .A(n_696), .Y(n_1004) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_702), .C(n_704), .Y(n_698) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g899 ( .A(n_701), .Y(n_899) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_712), .Y(n_883) );
AND2x2_ASAP7_75t_L g714 ( .A(n_715), .B(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AO22x1_ASAP7_75t_L g811 ( .A1(n_719), .A2(n_720), .B1(n_812), .B2(n_833), .Y(n_811) );
INVx2_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
XOR2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_744), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_734), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_723), .B(n_727), .C(n_730), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_742), .Y(n_738) );
INVx1_ASAP7_75t_SL g928 ( .A(n_740), .Y(n_928) );
INVx1_ASAP7_75t_L g864 ( .A(n_741), .Y(n_864) );
INVx1_ASAP7_75t_L g835 ( .A(n_746), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B1(n_779), .B2(n_834), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_764), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .C(n_761), .Y(n_752) );
OAI222xp33_ASAP7_75t_L g940 ( .A1(n_758), .A2(n_941), .B1(n_942), .B2(n_943), .C1(n_944), .C2(n_946), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_770), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx1_ASAP7_75t_L g862 ( .A(n_767), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_774), .Y(n_770) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g834 ( .A(n_779), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_780), .A2(n_781), .B1(n_810), .B2(n_811), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g809 ( .A(n_782), .Y(n_809) );
AND2x2_ASAP7_75t_SL g782 ( .A(n_783), .B(n_797), .Y(n_782) );
NOR3xp33_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .C(n_792), .Y(n_783) );
OAI21xp5_ASAP7_75t_SL g1080 ( .A1(n_788), .A2(n_1081), .B(n_1082), .Y(n_1080) );
OAI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_795), .B2(n_796), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_798), .B(n_804), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .Y(n_798) );
INVx2_ASAP7_75t_L g924 ( .A(n_800), .Y(n_924) );
HB1xp67_ASAP7_75t_L g1133 ( .A(n_800), .Y(n_1133) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g930 ( .A(n_806), .Y(n_930) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx3_ASAP7_75t_SL g833 ( .A(n_812), .Y(n_833) );
XOR2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_832), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g813 ( .A(n_814), .B(n_823), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g814 ( .A(n_815), .B(n_818), .Y(n_814) );
NAND3xp33_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .C(n_822), .Y(n_818) );
BUFx2_ASAP7_75t_L g851 ( .A(n_821), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_824), .B(n_828), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_829), .B(n_830), .Y(n_828) );
INVxp67_ASAP7_75t_L g1111 ( .A(n_838), .Y(n_1111) );
XNOR2xp5_ASAP7_75t_L g838 ( .A(n_839), .B(n_1024), .Y(n_838) );
XNOR2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_913), .Y(n_839) );
BUFx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_867), .B1(n_868), .B2(n_912), .Y(n_841) );
INVx2_ASAP7_75t_L g912 ( .A(n_842), .Y(n_912) );
XOR2x2_ASAP7_75t_L g842 ( .A(n_843), .B(n_866), .Y(n_842) );
NAND4xp75_ASAP7_75t_L g843 ( .A(n_844), .B(n_848), .C(n_855), .D(n_865), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_845), .B(n_847), .Y(n_844) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g1046 ( .A(n_854), .Y(n_1046) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_856), .B(n_860), .Y(n_855) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
OAI22xp5_ASAP7_75t_SL g868 ( .A1(n_869), .A2(n_888), .B1(n_889), .B2(n_911), .Y(n_868) );
INVx1_ASAP7_75t_L g911 ( .A(n_869), .Y(n_911) );
NAND3xp33_ASAP7_75t_L g870 ( .A(n_871), .B(n_880), .C(n_884), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_876), .Y(n_871) );
OAI21xp5_ASAP7_75t_SL g872 ( .A1(n_873), .A2(n_874), .B(n_875), .Y(n_872) );
OAI222xp33_ASAP7_75t_L g1002 ( .A1(n_873), .A2(n_1003), .B1(n_1004), .B2(n_1005), .C1(n_1006), .C2(n_1007), .Y(n_1002) );
NAND3xp33_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .C(n_879), .Y(n_876) );
AND2x2_ASAP7_75t_L g880 ( .A(n_881), .B(n_882), .Y(n_880) );
AND2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_887), .Y(n_884) );
INVx1_ASAP7_75t_SL g1097 ( .A(n_886), .Y(n_1097) );
INVx1_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
INVx1_ASAP7_75t_SL g910 ( .A(n_891), .Y(n_910) );
NAND3x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_900), .C(n_904), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_898), .Y(n_896) );
AND2x2_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
AND2x2_ASAP7_75t_L g904 ( .A(n_905), .B(n_907), .Y(n_904) );
BUFx2_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_915), .B1(n_978), .B2(n_1023), .Y(n_913) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_916), .A2(n_917), .B1(n_952), .B2(n_977), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g951 ( .A(n_919), .Y(n_951) );
AND2x2_ASAP7_75t_L g919 ( .A(n_920), .B(n_934), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_921), .B(n_927), .Y(n_920) );
OAI221xp5_ASAP7_75t_SL g921 ( .A1(n_922), .A2(n_923), .B1(n_924), .B2(n_925), .C(n_926), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_922), .A2(n_1095), .B1(n_1096), .B2(n_1097), .Y(n_1094) );
OAI221xp5_ASAP7_75t_SL g927 ( .A1(n_928), .A2(n_929), .B1(n_930), .B2(n_931), .C(n_932), .Y(n_927) );
NOR3xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_940), .C(n_947), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_939), .Y(n_935) );
OAI22xp5_ASAP7_75t_L g1139 ( .A1(n_937), .A2(n_939), .B1(n_1140), .B2(n_1141), .Y(n_1139) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g977 ( .A(n_952), .Y(n_977) );
INVx1_ASAP7_75t_SL g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g976 ( .A(n_954), .Y(n_976) );
AND2x2_ASAP7_75t_L g954 ( .A(n_955), .B(n_966), .Y(n_954) );
NOR2xp33_ASAP7_75t_SL g955 ( .A(n_956), .B(n_960), .Y(n_955) );
NOR2xp33_ASAP7_75t_L g966 ( .A(n_967), .B(n_971), .Y(n_966) );
NAND2xp33_ASAP7_75t_SL g971 ( .A(n_972), .B(n_973), .Y(n_971) );
INVx2_ASAP7_75t_L g1023 ( .A(n_978), .Y(n_1023) );
OA22x2_ASAP7_75t_SL g978 ( .A1(n_979), .A2(n_980), .B1(n_999), .B2(n_1022), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_979), .A2(n_980), .B1(n_1067), .B2(n_1107), .Y(n_1106) );
INVx1_ASAP7_75t_L g979 ( .A(n_980), .Y(n_979) );
XOR2x2_ASAP7_75t_L g980 ( .A(n_981), .B(n_998), .Y(n_980) );
NAND2x1_ASAP7_75t_L g981 ( .A(n_982), .B(n_991), .Y(n_981) );
NOR2xp33_ASAP7_75t_L g982 ( .A(n_983), .B(n_987), .Y(n_982) );
OAI21xp5_ASAP7_75t_SL g983 ( .A1(n_984), .A2(n_985), .B(n_986), .Y(n_983) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_989), .C(n_990), .Y(n_987) );
NOR2x1_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_996), .B(n_997), .Y(n_995) );
INVx1_ASAP7_75t_L g1022 ( .A(n_999), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1013), .Y(n_1000) );
NOR2xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1008), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1011), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1019), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1017), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
HB1xp67_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1027), .B1(n_1086), .B2(n_1109), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_1027), .Y(n_1026) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_1028), .A2(n_1053), .B1(n_1084), .B2(n_1085), .Y(n_1027) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1028), .Y(n_1084) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1030), .Y(n_1052) );
OR4x1_ASAP7_75t_L g1030 ( .A(n_1031), .B(n_1038), .C(n_1042), .D(n_1047), .Y(n_1030) );
INVx3_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
BUFx6f_ASAP7_75t_L g1072 ( .A(n_1037), .Y(n_1072) );
INVx1_ASAP7_75t_L g1085 ( .A(n_1053), .Y(n_1085) );
XNOR2xp5_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1067), .Y(n_1053) );
XOR2x2_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1066), .Y(n_1054) );
NAND4xp75_ASAP7_75t_L g1055 ( .A(n_1056), .B(n_1059), .C(n_1062), .D(n_1065), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1058), .Y(n_1056) );
AND2x2_ASAP7_75t_SL g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1064), .Y(n_1062) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_1067), .Y(n_1107) );
XOR2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1083), .Y(n_1067) );
NOR4xp75_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1073), .C(n_1077), .D(n_1080), .Y(n_1068) );
NAND2xp5_ASAP7_75t_SL g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
NAND2x1_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1076), .Y(n_1073) );
NAND2xp5_ASAP7_75t_SL g1077 ( .A(n_1078), .B(n_1079), .Y(n_1077) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_1086), .Y(n_1109) );
OA22x2_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1105), .B1(n_1106), .B2(n_1108), .Y(n_1086) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1087), .Y(n_1108) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1088), .Y(n_1104) );
AND4x1_ASAP7_75t_L g1088 ( .A(n_1089), .B(n_1093), .C(n_1098), .D(n_1102), .Y(n_1088) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
NOR2x1_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1118), .Y(n_1113) );
OR2x2_ASAP7_75t_SL g1155 ( .A(n_1114), .B(n_1119), .Y(n_1155) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_1115), .B(n_1117), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1151 ( .A(n_1115), .B(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1116), .B(n_1152), .Y(n_1157) );
CKINVDCx16_ASAP7_75t_R g1152 ( .A(n_1117), .Y(n_1152) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_1119), .Y(n_1118) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1122 ( .A(n_1123), .B(n_1124), .Y(n_1122) );
OAI222xp33_ASAP7_75t_L g1125 ( .A1(n_1126), .A2(n_1151), .B1(n_1153), .B2(n_1154), .C1(n_1155), .C2(n_1156), .Y(n_1125) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1127), .Y(n_1150) );
AND2x2_ASAP7_75t_SL g1127 ( .A(n_1128), .B(n_1138), .Y(n_1127) );
NOR2xp33_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1134), .Y(n_1128) );
NOR3xp33_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1142), .C(n_1146), .Y(n_1138) );
endmodule