module fake_aes_3447_n_464 (n_53, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_464);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_464;
wire n_117;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_455;
wire n_137;
wire n_277;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_442;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_69;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_245;
wire n_70;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_458;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_68;
wire n_123;
wire n_457;
wire n_223;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g66 ( .A(n_34), .Y(n_66) );
CKINVDCx5p33_ASAP7_75t_R g67 ( .A(n_7), .Y(n_67) );
INVx1_ASAP7_75t_L g68 ( .A(n_9), .Y(n_68) );
INVxp67_ASAP7_75t_SL g69 ( .A(n_50), .Y(n_69) );
INVxp67_ASAP7_75t_SL g70 ( .A(n_36), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_22), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_24), .Y(n_72) );
INVxp67_ASAP7_75t_L g73 ( .A(n_0), .Y(n_73) );
INVxp67_ASAP7_75t_L g74 ( .A(n_29), .Y(n_74) );
INVxp67_ASAP7_75t_SL g75 ( .A(n_6), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_65), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_57), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_64), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_3), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_2), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_43), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_60), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_53), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_63), .Y(n_85) );
INVxp33_ASAP7_75t_SL g86 ( .A(n_32), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_28), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_51), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_25), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_49), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_45), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_39), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_38), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_8), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_27), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_21), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_42), .Y(n_98) );
BUFx3_ASAP7_75t_L g99 ( .A(n_66), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_66), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_67), .Y(n_101) );
INVxp67_ASAP7_75t_L g102 ( .A(n_96), .Y(n_102) );
INVx3_ASAP7_75t_L g103 ( .A(n_79), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_71), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_87), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_71), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_73), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_68), .B(n_0), .Y(n_111) );
OA21x2_ASAP7_75t_L g112 ( .A1(n_72), .A2(n_98), .B(n_97), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_74), .B(n_1), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_79), .B(n_1), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_86), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_95), .Y(n_118) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_80), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_119) );
AND2x4_ASAP7_75t_L g120 ( .A(n_80), .B(n_4), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_82), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_106), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_99), .B(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_106), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_120), .B(n_93), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_106), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_102), .B(n_88), .Y(n_127) );
NOR2x1p5_ASAP7_75t_L g128 ( .A(n_105), .B(n_75), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_106), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_120), .B(n_93), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_106), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_106), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_100), .A2(n_98), .B1(n_97), .B2(n_94), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_102), .B(n_83), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_99), .B(n_84), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_121), .B(n_89), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_112), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_116), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_120), .A2(n_94), .B1(n_92), .B2(n_91), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_120), .B(n_92), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_112), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_116), .Y(n_144) );
INVxp67_ASAP7_75t_SL g145 ( .A(n_108), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_112), .Y(n_146) );
BUFx2_ASAP7_75t_L g147 ( .A(n_145), .Y(n_147) );
OAI21xp5_ASAP7_75t_L g148 ( .A1(n_138), .A2(n_112), .B(n_108), .Y(n_148) );
NOR3xp33_ASAP7_75t_SL g149 ( .A(n_135), .B(n_118), .C(n_117), .Y(n_149) );
BUFx2_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_125), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_139), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_128), .Y(n_153) );
NOR2x1_ASAP7_75t_L g154 ( .A(n_128), .B(n_107), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_125), .Y(n_155) );
INVx5_ASAP7_75t_L g156 ( .A(n_144), .Y(n_156) );
INVx2_ASAP7_75t_SL g157 ( .A(n_125), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_140), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_127), .B(n_107), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_129), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_140), .B(n_116), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_144), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_127), .B(n_100), .Y(n_163) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_137), .A2(n_110), .B1(n_101), .B2(n_114), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_139), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_125), .B(n_130), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_142), .B(n_115), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_125), .B(n_114), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_130), .B(n_111), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
AND2x4_ASAP7_75t_L g173 ( .A(n_130), .B(n_119), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
OR2x2_ASAP7_75t_L g176 ( .A(n_137), .B(n_111), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_142), .A2(n_130), .B1(n_144), .B2(n_141), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_130), .B(n_104), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_149), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_148), .A2(n_146), .B(n_143), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
AOI22xp5_ASAP7_75t_L g184 ( .A1(n_173), .A2(n_142), .B1(n_144), .B2(n_141), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_147), .B(n_144), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_156), .B(n_142), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_173), .A2(n_142), .B1(n_141), .B2(n_133), .Y(n_187) );
AOI221xp5_ASAP7_75t_L g188 ( .A1(n_173), .A2(n_133), .B1(n_113), .B2(n_104), .C(n_115), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_166), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_166), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g191 ( .A1(n_147), .A2(n_141), .B1(n_146), .B2(n_143), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_152), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_168), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_176), .B(n_141), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_150), .B(n_176), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
AND2x2_ASAP7_75t_L g198 ( .A(n_150), .B(n_123), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_168), .B(n_119), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_153), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_168), .B(n_123), .Y(n_203) );
INVxp67_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_156), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_153), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_163), .B(n_143), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_177), .B(n_146), .Y(n_208) );
BUFx2_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_158), .Y(n_210) );
INVxp67_ASAP7_75t_L g211 ( .A(n_161), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_197), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_197), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_200), .A2(n_158), .B1(n_171), .B2(n_169), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_189), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_196), .B(n_151), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_192), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_197), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_192), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_197), .Y(n_220) );
OR2x2_ASAP7_75t_L g221 ( .A(n_196), .B(n_204), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_184), .B(n_162), .Y(n_222) );
CKINVDCx11_ASAP7_75t_R g223 ( .A(n_201), .Y(n_223) );
AOI22xp33_ASAP7_75t_L g224 ( .A1(n_200), .A2(n_165), .B1(n_172), .B2(n_175), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_189), .Y(n_225) );
NAND3xp33_ASAP7_75t_L g226 ( .A(n_188), .B(n_164), .C(n_170), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_198), .B(n_151), .Y(n_227) );
OR2x6_ASAP7_75t_L g228 ( .A(n_194), .B(n_155), .Y(n_228) );
NAND3xp33_ASAP7_75t_L g229 ( .A(n_188), .B(n_154), .C(n_113), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_198), .B(n_155), .Y(n_230) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_209), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_189), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_200), .A2(n_172), .B1(n_165), .B2(n_175), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_193), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_187), .B(n_157), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_200), .B1(n_187), .B2(n_184), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g237 ( .A1(n_221), .A2(n_210), .B1(n_180), .B2(n_211), .Y(n_237) );
OAI221xp5_ASAP7_75t_L g238 ( .A1(n_221), .A2(n_195), .B1(n_194), .B2(n_206), .C(n_203), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_221), .B(n_203), .Y(n_239) );
OAI21x1_ASAP7_75t_L g240 ( .A1(n_215), .A2(n_182), .B(n_183), .Y(n_240) );
AOI221xp5_ASAP7_75t_L g241 ( .A1(n_226), .A2(n_185), .B1(n_178), .B2(n_99), .C(n_208), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_223), .Y(n_242) );
AOI221xp5_ASAP7_75t_L g243 ( .A1(n_214), .A2(n_185), .B1(n_208), .B2(n_136), .C(n_103), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_216), .B(n_207), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_216), .B(n_207), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_222), .A2(n_209), .B1(n_186), .B2(n_193), .Y(n_246) );
OA21x2_ASAP7_75t_L g247 ( .A1(n_215), .A2(n_181), .B(n_202), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_157), .B1(n_191), .B2(n_136), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_235), .A2(n_109), .B1(n_189), .B2(n_179), .Y(n_249) );
OAI221xp5_ASAP7_75t_L g250 ( .A1(n_214), .A2(n_109), .B1(n_205), .B2(n_103), .C(n_162), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_231), .Y(n_251) );
INVxp33_ASAP7_75t_L g252 ( .A(n_231), .Y(n_252) );
OAI22xp33_ASAP7_75t_L g253 ( .A1(n_235), .A2(n_156), .B1(n_167), .B2(n_179), .Y(n_253) );
OAI22xp33_ASAP7_75t_L g254 ( .A1(n_228), .A2(n_156), .B1(n_167), .B2(n_179), .Y(n_254) );
AOI33xp33_ASAP7_75t_L g255 ( .A1(n_224), .A2(n_109), .A3(n_77), .B1(n_78), .B2(n_81), .B3(n_91), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_244), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_244), .B(n_217), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_247), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_245), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_245), .Y(n_260) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_242), .Y(n_261) );
AND2x2_ASAP7_75t_L g262 ( .A(n_239), .B(n_217), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_247), .Y(n_263) );
INVxp67_ASAP7_75t_SL g264 ( .A(n_249), .Y(n_264) );
OAI31xp33_ASAP7_75t_L g265 ( .A1(n_238), .A2(n_222), .A3(n_216), .B(n_229), .Y(n_265) );
INVxp67_ASAP7_75t_SL g266 ( .A(n_249), .Y(n_266) );
AND2x4_ASAP7_75t_L g267 ( .A(n_240), .B(n_212), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_247), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_236), .B(n_219), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_239), .B(n_219), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_240), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_251), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_236), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
NAND3xp33_ASAP7_75t_SL g276 ( .A(n_243), .B(n_220), .C(n_212), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_248), .B(n_234), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_257), .B(n_234), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_258), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_258), .Y(n_280) );
OAI31xp33_ASAP7_75t_L g281 ( .A1(n_265), .A2(n_237), .A3(n_222), .B(n_229), .Y(n_281) );
OAI211xp5_ASAP7_75t_SL g282 ( .A1(n_265), .A2(n_103), .B(n_90), .C(n_77), .Y(n_282) );
NAND2x1_ASAP7_75t_L g283 ( .A(n_267), .B(n_212), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_273), .Y(n_284) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_273), .B(n_78), .C(n_81), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g286 ( .A1(n_274), .A2(n_222), .B1(n_246), .B2(n_252), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_270), .B(n_248), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_257), .B(n_112), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_258), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_268), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_261), .B(n_69), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_257), .B(n_220), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g294 ( .A1(n_275), .A2(n_250), .B1(n_103), .B2(n_224), .C(n_233), .Y(n_294) );
NAND4xp25_ASAP7_75t_L g295 ( .A(n_275), .B(n_233), .C(n_241), .D(n_227), .Y(n_295) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
AND3x2_ASAP7_75t_L g297 ( .A(n_261), .B(n_70), .C(n_227), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_270), .B(n_218), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_268), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_267), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_273), .A2(n_228), .B1(n_212), .B2(n_213), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_256), .B(n_227), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_263), .Y(n_303) );
INVx1_ASAP7_75t_SL g304 ( .A(n_263), .Y(n_304) );
OAI22xp33_ASAP7_75t_SL g305 ( .A1(n_256), .A2(n_212), .B1(n_213), .B2(n_228), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_267), .B(n_213), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_269), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_269), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_259), .A2(n_228), .B1(n_213), .B2(n_218), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_290), .B(n_269), .Y(n_310) );
NOR2xp33_ASAP7_75t_R g311 ( .A(n_297), .B(n_259), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_300), .B(n_270), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_306), .Y(n_313) );
OAI33xp33_ASAP7_75t_L g314 ( .A1(n_305), .A2(n_282), .A3(n_299), .B1(n_285), .B2(n_309), .B3(n_287), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_296), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_289), .B(n_274), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_278), .B(n_277), .Y(n_317) );
NOR3xp33_ASAP7_75t_L g318 ( .A(n_291), .B(n_276), .C(n_213), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_289), .Y(n_319) );
BUFx3_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_283), .B(n_267), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_293), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_304), .B(n_277), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g324 ( .A(n_281), .B(n_267), .C(n_260), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_287), .B(n_277), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_284), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_302), .B(n_262), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_289), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_288), .B(n_262), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
OAI211xp5_ASAP7_75t_L g332 ( .A1(n_281), .A2(n_271), .B(n_262), .C(n_266), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_298), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVxp67_ASAP7_75t_SL g336 ( .A(n_280), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_305), .B(n_271), .Y(n_337) );
OAI33xp33_ASAP7_75t_L g338 ( .A1(n_295), .A2(n_253), .A3(n_6), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_295), .B(n_271), .Y(n_339) );
NAND3xp33_ASAP7_75t_SL g340 ( .A(n_301), .B(n_5), .C(n_10), .Y(n_340) );
NAND5xp2_ASAP7_75t_SL g341 ( .A(n_286), .B(n_5), .C(n_10), .D(n_11), .E(n_12), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_292), .B(n_272), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
OAI21xp5_ASAP7_75t_L g345 ( .A1(n_288), .A2(n_266), .B(n_264), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_306), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_303), .B(n_307), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_306), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_307), .B(n_272), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_313), .B(n_308), .Y(n_350) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_335), .Y(n_351) );
INVx1_ASAP7_75t_SL g352 ( .A(n_325), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g353 ( .A1(n_340), .A2(n_294), .B(n_306), .Y(n_353) );
AO22x1_ASAP7_75t_L g354 ( .A1(n_321), .A2(n_264), .B1(n_272), .B2(n_218), .Y(n_354) );
NAND3xp33_ASAP7_75t_L g355 ( .A(n_318), .B(n_129), .C(n_134), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_337), .A2(n_228), .B1(n_254), .B2(n_232), .Y(n_356) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_337), .A2(n_228), .B1(n_232), .B2(n_225), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_348), .B(n_12), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_339), .A2(n_225), .B1(n_215), .B2(n_230), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_348), .B(n_13), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_315), .A2(n_13), .B(n_14), .Y(n_361) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_320), .B(n_225), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_230), .B(n_134), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_199), .B1(n_190), .B2(n_183), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_322), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_310), .B(n_15), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_333), .B(n_15), .Y(n_367) );
NAND2xp33_ASAP7_75t_SL g368 ( .A(n_311), .B(n_16), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_325), .Y(n_369) );
INVxp67_ASAP7_75t_L g370 ( .A(n_310), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_346), .B(n_16), .Y(n_371) );
NAND2xp33_ASAP7_75t_L g372 ( .A(n_327), .B(n_189), .Y(n_372) );
INVx1_ASAP7_75t_SL g373 ( .A(n_320), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_314), .A2(n_122), .B1(n_124), .B2(n_126), .C(n_131), .Y(n_374) );
AOI21xp33_ASAP7_75t_L g375 ( .A1(n_345), .A2(n_17), .B(n_18), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_338), .A2(n_202), .B1(n_199), .B2(n_190), .Y(n_376) );
OAI32xp33_ASAP7_75t_L g377 ( .A1(n_312), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_202), .Y(n_377) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_312), .A2(n_19), .B(n_134), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_323), .Y(n_379) );
OAI21xp33_ASAP7_75t_SL g380 ( .A1(n_336), .A2(n_199), .B(n_190), .Y(n_380) );
OAI32xp33_ASAP7_75t_L g381 ( .A1(n_323), .A2(n_183), .A3(n_181), .B1(n_132), .B2(n_131), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_347), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_319), .Y(n_383) );
AND2x4_ASAP7_75t_L g384 ( .A(n_347), .B(n_20), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_330), .B(n_23), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_317), .B(n_132), .Y(n_386) );
OAI22xp33_ASAP7_75t_L g387 ( .A1(n_328), .A2(n_189), .B1(n_181), .B2(n_179), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
AND3x2_ASAP7_75t_L g389 ( .A(n_341), .B(n_26), .C(n_30), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_344), .B(n_126), .C(n_124), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_382), .B(n_316), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_368), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_360), .Y(n_393) );
NOR3xp33_ASAP7_75t_SL g394 ( .A(n_353), .B(n_326), .C(n_341), .Y(n_394) );
NAND4xp25_ASAP7_75t_SL g395 ( .A(n_353), .B(n_343), .C(n_334), .D(n_331), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_379), .B(n_316), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_370), .B(n_349), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g398 ( .A1(n_354), .A2(n_343), .B(n_334), .C(n_331), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_365), .B(n_349), .Y(n_399) );
XOR2x2_ASAP7_75t_L g400 ( .A(n_389), .B(n_342), .Y(n_400) );
NAND2xp33_ASAP7_75t_SL g401 ( .A(n_360), .B(n_342), .Y(n_401) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_380), .B(n_122), .Y(n_402) );
NAND2x1_ASAP7_75t_L g403 ( .A(n_357), .B(n_31), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_351), .B(n_33), .Y(n_404) );
XOR2x2_ASAP7_75t_L g405 ( .A(n_358), .B(n_35), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_352), .B(n_37), .Y(n_406) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_373), .B(n_40), .Y(n_407) );
NOR3xp33_ASAP7_75t_L g408 ( .A(n_355), .B(n_174), .C(n_160), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g409 ( .A(n_373), .B(n_44), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_383), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_350), .B(n_46), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_388), .B(n_47), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_366), .B(n_48), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_352), .B(n_52), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_369), .B(n_54), .Y(n_415) );
INVxp67_ASAP7_75t_L g416 ( .A(n_369), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_367), .B(n_55), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_362), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_371), .B(n_56), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g420 ( .A(n_356), .B(n_58), .Y(n_420) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_384), .B(n_59), .Y(n_421) );
AOI211xp5_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_375), .B(n_377), .C(n_359), .Y(n_422) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_420), .A2(n_363), .B(n_361), .Y(n_423) );
AOI221xp5_ASAP7_75t_SL g424 ( .A1(n_416), .A2(n_378), .B1(n_364), .B2(n_386), .C(n_372), .Y(n_424) );
NOR2x1p5_ASAP7_75t_SL g425 ( .A(n_414), .B(n_385), .Y(n_425) );
XNOR2xp5_ASAP7_75t_L g426 ( .A(n_405), .B(n_384), .Y(n_426) );
AOI221xp5_ASAP7_75t_SL g427 ( .A1(n_420), .A2(n_397), .B1(n_399), .B2(n_396), .C(n_391), .Y(n_427) );
OAI31xp33_ASAP7_75t_L g428 ( .A1(n_401), .A2(n_387), .A3(n_390), .B(n_381), .Y(n_428) );
OAI22xp33_ASAP7_75t_SL g429 ( .A1(n_393), .A2(n_376), .B1(n_374), .B2(n_62), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_392), .A2(n_160), .B1(n_174), .B2(n_61), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_410), .B(n_393), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_421), .Y(n_432) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_394), .A2(n_401), .B1(n_405), .B2(n_398), .C(n_403), .Y(n_433) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_395), .A2(n_409), .B(n_407), .Y(n_434) );
XOR2x2_ASAP7_75t_L g435 ( .A(n_400), .B(n_407), .Y(n_435) );
NOR2x1_ASAP7_75t_L g436 ( .A(n_409), .B(n_418), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_418), .B(n_402), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_404), .B(n_417), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_400), .B(n_406), .Y(n_440) );
NAND4xp75_ASAP7_75t_L g441 ( .A(n_427), .B(n_419), .C(n_415), .D(n_413), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_433), .A2(n_402), .B(n_411), .C(n_412), .Y(n_442) );
BUFx8_ASAP7_75t_SL g443 ( .A(n_440), .Y(n_443) );
NAND2xp33_ASAP7_75t_R g444 ( .A(n_434), .B(n_408), .Y(n_444) );
AOI211xp5_ASAP7_75t_L g445 ( .A1(n_429), .A2(n_426), .B(n_432), .C(n_428), .Y(n_445) );
OAI21xp5_ASAP7_75t_SL g446 ( .A1(n_437), .A2(n_436), .B(n_423), .Y(n_446) );
AOI211xp5_ASAP7_75t_L g447 ( .A1(n_422), .A2(n_424), .B(n_439), .C(n_435), .Y(n_447) );
AOI211xp5_ASAP7_75t_SL g448 ( .A1(n_439), .A2(n_430), .B(n_431), .C(n_438), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_425), .A2(n_435), .B1(n_392), .B2(n_433), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_433), .B(n_392), .C(n_428), .Y(n_450) );
OA22x2_ASAP7_75t_L g451 ( .A1(n_440), .A2(n_426), .B1(n_432), .B2(n_393), .Y(n_451) );
INVx1_ASAP7_75t_SL g452 ( .A(n_432), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g453 ( .A(n_443), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_444), .Y(n_454) );
CKINVDCx20_ASAP7_75t_R g455 ( .A(n_443), .Y(n_455) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_449), .A2(n_447), .B1(n_446), .B2(n_445), .C(n_450), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_456), .A2(n_449), .B1(n_444), .B2(n_451), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_454), .Y(n_458) );
AND3x4_ASAP7_75t_L g459 ( .A(n_455), .B(n_441), .C(n_442), .Y(n_459) );
NOR2x1p5_ASAP7_75t_L g460 ( .A(n_458), .B(n_453), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_459), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_460), .Y(n_462) );
NAND3x1_ASAP7_75t_L g463 ( .A(n_462), .B(n_461), .C(n_457), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_463), .A2(n_452), .B(n_448), .Y(n_464) );
endmodule