module real_aes_7018_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_716, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_716;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_417;
wire n_182;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_527;
wire n_434;
wire n_505;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_0), .A2(n_172), .B(n_173), .C(n_177), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_1), .B(n_166), .Y(n_179) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g150 ( .A(n_3), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_4), .A2(n_140), .B(n_157), .C(n_467), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_5), .A2(n_160), .B(n_488), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_6), .A2(n_160), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_7), .B(n_166), .Y(n_494) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_8), .A2(n_132), .B(n_219), .Y(n_218) );
AND2x6_ASAP7_75t_L g157 ( .A(n_9), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g236 ( .A1(n_10), .A2(n_140), .B(n_157), .C(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g459 ( .A(n_11), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_12), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_12), .B(n_40), .Y(n_424) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_13), .B(n_176), .Y(n_469) );
INVx1_ASAP7_75t_L g137 ( .A(n_14), .Y(n_137) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_15), .B(n_151), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_16), .A2(n_152), .B(n_478), .C(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_17), .B(n_166), .Y(n_481) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_18), .A2(n_66), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_18), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_19), .B(n_209), .Y(n_528) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_20), .A2(n_140), .B(n_203), .C(n_208), .Y(n_202) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_21), .A2(n_175), .B(n_227), .C(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_22), .B(n_176), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_23), .B(n_176), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g497 ( .A(n_24), .Y(n_497) );
INVx1_ASAP7_75t_L g509 ( .A(n_25), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_26), .A2(n_140), .B(n_208), .C(n_222), .Y(n_221) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_27), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_28), .Y(n_465) );
INVx1_ASAP7_75t_L g526 ( .A(n_29), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_30), .A2(n_160), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g142 ( .A(n_31), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_32), .A2(n_155), .B(n_187), .C(n_188), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_33), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g490 ( .A1(n_34), .A2(n_175), .B(n_491), .C(n_493), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g120 ( .A1(n_35), .A2(n_121), .B1(n_416), .B2(n_417), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_35), .Y(n_416) );
INVxp67_ASAP7_75t_L g527 ( .A(n_36), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_37), .B(n_224), .Y(n_223) );
CKINVDCx14_ASAP7_75t_R g489 ( .A(n_38), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_39), .A2(n_140), .B(n_208), .C(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g113 ( .A(n_40), .Y(n_113) );
AOI222xp33_ASAP7_75t_L g430 ( .A1(n_41), .A2(n_431), .B1(n_699), .B2(n_700), .C1(n_706), .C2(n_710), .Y(n_430) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_42), .A2(n_177), .B(n_457), .C(n_458), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g103 ( .A1(n_43), .A2(n_104), .B1(n_105), .B2(n_114), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_44), .B(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_45), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_46), .B(n_151), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_47), .B(n_160), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_48), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_49), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_50), .A2(n_155), .B(n_187), .C(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g174 ( .A(n_51), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_52), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_52), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_53), .A2(n_84), .B1(n_704), .B2(n_705), .Y(n_703) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_53), .Y(n_705) );
INVx1_ASAP7_75t_L g249 ( .A(n_54), .Y(n_249) );
INVx1_ASAP7_75t_L g447 ( .A(n_55), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_56), .B(n_160), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_57), .Y(n_212) );
CKINVDCx14_ASAP7_75t_R g455 ( .A(n_58), .Y(n_455) );
INVx1_ASAP7_75t_L g158 ( .A(n_59), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_60), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_61), .B(n_166), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_62), .A2(n_147), .B(n_207), .C(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g136 ( .A(n_63), .Y(n_136) );
INVx1_ASAP7_75t_SL g492 ( .A(n_64), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_65), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_66), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_67), .B(n_151), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_68), .B(n_166), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_69), .B(n_152), .Y(n_238) );
INVx1_ASAP7_75t_L g500 ( .A(n_70), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_71), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_72), .B(n_191), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_73), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g263 ( .A(n_74), .Y(n_263) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_76), .A2(n_160), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_77), .B(n_426), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_78), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_79), .A2(n_160), .B(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_80), .A2(n_201), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g476 ( .A(n_81), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g506 ( .A(n_82), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_83), .B(n_190), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_84), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_85), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_86), .A2(n_160), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g479 ( .A(n_87), .Y(n_479) );
INVx2_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx1_ASAP7_75t_L g468 ( .A(n_89), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_90), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_91), .B(n_176), .Y(n_239) );
INVx2_ASAP7_75t_L g108 ( .A(n_92), .Y(n_108) );
OR2x2_ASAP7_75t_L g421 ( .A(n_92), .B(n_422), .Y(n_421) );
OR2x2_ASAP7_75t_L g434 ( .A(n_92), .B(n_423), .Y(n_434) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_93), .A2(n_140), .B(n_155), .C(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_94), .B(n_160), .Y(n_185) );
INVx1_ASAP7_75t_L g189 ( .A(n_95), .Y(n_189) );
INVxp67_ASAP7_75t_L g266 ( .A(n_96), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_97), .B(n_132), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_98), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx1_ASAP7_75t_L g234 ( .A(n_100), .Y(n_234) );
INVx2_ASAP7_75t_L g450 ( .A(n_101), .Y(n_450) );
AND2x2_ASAP7_75t_L g251 ( .A(n_102), .B(n_194), .Y(n_251) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g423 ( .A(n_107), .B(n_424), .Y(n_423) );
OR2x2_ASAP7_75t_L g437 ( .A(n_108), .B(n_423), .Y(n_437) );
NOR2x2_ASAP7_75t_L g712 ( .A(n_108), .B(n_422), .Y(n_712) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B(n_429), .Y(n_114) );
HB1xp67_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g714 ( .A(n_117), .Y(n_714) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
OAI21xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_418), .B(n_425), .Y(n_119) );
INVx1_ASAP7_75t_L g417 ( .A(n_121), .Y(n_417) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
INVx2_ASAP7_75t_L g435 ( .A(n_125), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_125), .A2(n_433), .B1(n_708), .B2(n_709), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g125 ( .A(n_126), .B(n_359), .Y(n_125) );
AND4x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_299), .C(n_314), .D(n_339), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g127 ( .A(n_128), .B(n_272), .Y(n_127) );
OAI21xp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_180), .B(n_252), .Y(n_128) );
AND2x2_ASAP7_75t_L g302 ( .A(n_129), .B(n_198), .Y(n_302) );
AND2x2_ASAP7_75t_L g315 ( .A(n_129), .B(n_197), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_129), .B(n_181), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_129), .Y(n_369) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
INVx2_ASAP7_75t_L g286 ( .A(n_130), .Y(n_286) );
BUFx2_ASAP7_75t_L g313 ( .A(n_130), .Y(n_313) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_138), .B(n_163), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_131), .B(n_164), .Y(n_163) );
INVx3_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_131), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_131), .A2(n_233), .B(n_240), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_131), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_131), .A2(n_496), .B(n_502), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_131), .B(n_512), .Y(n_511) );
INVx4_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_132), .A2(n_220), .B(n_221), .Y(n_219) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_132), .Y(n_260) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_L g242 ( .A(n_133), .Y(n_242) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x2_ASAP7_75t_SL g194 ( .A(n_134), .B(n_135), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_159), .Y(n_138) );
INVx5_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_141), .Y(n_154) );
BUFx3_ASAP7_75t_L g178 ( .A(n_141), .Y(n_178) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
INVx1_ASAP7_75t_L g228 ( .A(n_142), .Y(n_228) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_144), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
AND2x2_ASAP7_75t_L g161 ( .A(n_144), .B(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
INVx1_ASAP7_75t_L g224 ( .A(n_144), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g449 ( .A(n_148), .B(n_450), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_148), .B(n_479), .Y(n_478) );
OAI22xp33_ASAP7_75t_L g525 ( .A1(n_148), .A2(n_151), .B1(n_526), .B2(n_527), .Y(n_525) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g191 ( .A(n_149), .Y(n_191) );
INVx2_ASAP7_75t_L g172 ( .A(n_151), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_151), .B(n_266), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g508 ( .A1(n_151), .A2(n_206), .B(n_509), .C(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_152), .B(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx3_ASAP7_75t_L g493 ( .A(n_154), .Y(n_493) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_156), .A2(n_169), .B(n_170), .C(n_171), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_156), .A2(n_170), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_SL g446 ( .A1(n_156), .A2(n_170), .B(n_447), .C(n_448), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_156), .A2(n_170), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_156), .A2(n_170), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_156), .A2(n_170), .B(n_489), .C(n_490), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_SL g522 ( .A1(n_156), .A2(n_170), .B(n_523), .C(n_524), .Y(n_522) );
INVx4_ASAP7_75t_SL g156 ( .A(n_157), .Y(n_156) );
AND2x4_ASAP7_75t_L g160 ( .A(n_157), .B(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g208 ( .A(n_157), .Y(n_208) );
NAND2x1p5_ASAP7_75t_L g235 ( .A(n_157), .B(n_161), .Y(n_235) );
BUFx2_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
INVx1_ASAP7_75t_L g207 ( .A(n_162), .Y(n_207) );
AND2x2_ASAP7_75t_L g253 ( .A(n_165), .B(n_198), .Y(n_253) );
INVx2_ASAP7_75t_L g269 ( .A(n_165), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_165), .B(n_197), .Y(n_278) );
AND2x2_ASAP7_75t_L g357 ( .A(n_165), .B(n_286), .Y(n_357) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_179), .Y(n_165) );
INVx2_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_175), .B(n_492), .Y(n_491) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g457 ( .A(n_176), .Y(n_457) );
INVx2_ASAP7_75t_L g470 ( .A(n_177), .Y(n_470) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_178), .Y(n_193) );
INVx1_ASAP7_75t_L g480 ( .A(n_178), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_214), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_181), .B(n_284), .Y(n_322) );
INVx1_ASAP7_75t_L g410 ( .A(n_181), .Y(n_410) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
AND2x2_ASAP7_75t_L g268 ( .A(n_182), .B(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g282 ( .A(n_182), .B(n_283), .Y(n_282) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_182), .Y(n_311) );
OR2x2_ASAP7_75t_L g343 ( .A(n_182), .B(n_285), .Y(n_343) );
AND2x2_ASAP7_75t_L g351 ( .A(n_182), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g384 ( .A(n_182), .B(n_353), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_182), .B(n_253), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_182), .B(n_313), .Y(n_409) );
AND2x2_ASAP7_75t_L g415 ( .A(n_182), .B(n_302), .Y(n_415) );
INVx5_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx2_ASAP7_75t_L g275 ( .A(n_183), .Y(n_275) );
AND2x2_ASAP7_75t_L g305 ( .A(n_183), .B(n_285), .Y(n_305) );
AND2x2_ASAP7_75t_L g338 ( .A(n_183), .B(n_298), .Y(n_338) );
AND2x2_ASAP7_75t_L g358 ( .A(n_183), .B(n_198), .Y(n_358) );
AND2x2_ASAP7_75t_L g392 ( .A(n_183), .B(n_258), .Y(n_392) );
OR2x6_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_194), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_192), .C(n_193), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_190), .A2(n_193), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp5_ASAP7_75t_L g467 ( .A1(n_190), .A2(n_468), .B(n_469), .C(n_470), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g499 ( .A1(n_190), .A2(n_470), .B(n_500), .C(n_501), .Y(n_499) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g210 ( .A(n_194), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_194), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_194), .A2(n_246), .B(n_247), .Y(n_245) );
OA21x2_ASAP7_75t_L g452 ( .A1(n_194), .A2(n_453), .B(n_460), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_194), .A2(n_235), .B(n_506), .C(n_507), .Y(n_505) );
AND2x4_ASAP7_75t_L g298 ( .A(n_197), .B(n_269), .Y(n_298) );
AND2x2_ASAP7_75t_L g309 ( .A(n_197), .B(n_305), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_197), .B(n_285), .Y(n_348) );
INVx2_ASAP7_75t_L g363 ( .A(n_197), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_197), .B(n_297), .Y(n_386) );
AND2x2_ASAP7_75t_L g405 ( .A(n_197), .B(n_357), .Y(n_405) );
INVx5_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_198), .Y(n_304) );
AND2x2_ASAP7_75t_L g312 ( .A(n_198), .B(n_313), .Y(n_312) );
AND2x4_ASAP7_75t_L g353 ( .A(n_198), .B(n_269), .Y(n_353) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_211), .Y(n_198) );
AOI21xp5_ASAP7_75t_SL g199 ( .A1(n_200), .A2(n_202), .B(n_209), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_206), .Y(n_203) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_207), .B(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_210), .B(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
AO21x2_ASAP7_75t_L g463 ( .A1(n_213), .A2(n_464), .B(n_471), .Y(n_463) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_229), .Y(n_215) );
AND2x2_ASAP7_75t_L g276 ( .A(n_216), .B(n_259), .Y(n_276) );
INVx1_ASAP7_75t_SL g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_217), .B(n_232), .Y(n_256) );
OR2x2_ASAP7_75t_L g289 ( .A(n_217), .B(n_259), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_217), .B(n_259), .Y(n_294) );
AND2x2_ASAP7_75t_L g321 ( .A(n_217), .B(n_258), .Y(n_321) );
AND2x2_ASAP7_75t_L g373 ( .A(n_217), .B(n_231), .Y(n_373) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_218), .B(n_243), .Y(n_281) );
AND2x2_ASAP7_75t_L g317 ( .A(n_218), .B(n_232), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_225), .B(n_226), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_226), .A2(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_229), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
OR2x2_ASAP7_75t_L g307 ( .A(n_230), .B(n_289), .Y(n_307) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_243), .Y(n_230) );
OAI322xp33_ASAP7_75t_L g272 ( .A1(n_231), .A2(n_273), .A3(n_277), .B1(n_279), .B2(n_282), .C1(n_287), .C2(n_295), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_231), .B(n_258), .Y(n_280) );
OR2x2_ASAP7_75t_L g290 ( .A(n_231), .B(n_244), .Y(n_290) );
AND2x2_ASAP7_75t_L g292 ( .A(n_231), .B(n_244), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_231), .B(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_231), .B(n_259), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_231), .B(n_388), .Y(n_387) );
INVx5_ASAP7_75t_SL g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_232), .B(n_276), .Y(n_402) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_236), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_235), .A2(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_235), .A2(n_497), .B(n_498), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx2_ASAP7_75t_L g520 ( .A(n_242), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_243), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g270 ( .A(n_243), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_243), .B(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g332 ( .A(n_243), .B(n_259), .Y(n_332) );
AOI211xp5_ASAP7_75t_SL g360 ( .A1(n_243), .A2(n_361), .B(n_364), .C(n_376), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_243), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g398 ( .A(n_243), .B(n_373), .Y(n_398) );
INVx5_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g326 ( .A(n_244), .B(n_259), .Y(n_326) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_244), .Y(n_335) );
AND2x2_ASAP7_75t_L g375 ( .A(n_244), .B(n_373), .Y(n_375) );
AND2x2_ASAP7_75t_SL g406 ( .A(n_244), .B(n_276), .Y(n_406) );
AND2x2_ASAP7_75t_L g413 ( .A(n_244), .B(n_372), .Y(n_413) );
OR2x6_ASAP7_75t_L g244 ( .A(n_245), .B(n_251), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B1(n_268), .B2(n_270), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_253), .B(n_275), .Y(n_323) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx1_ASAP7_75t_L g271 ( .A(n_256), .Y(n_271) );
OR2x2_ASAP7_75t_L g331 ( .A(n_256), .B(n_332), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g379 ( .A1(n_256), .A2(n_380), .B1(n_382), .B2(n_383), .C(n_385), .Y(n_379) );
INVx2_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
AND2x2_ASAP7_75t_L g291 ( .A(n_258), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g381 ( .A(n_258), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_258), .B(n_373), .Y(n_394) );
INVx3_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVxp67_ASAP7_75t_L g336 ( .A(n_259), .Y(n_336) );
AND2x2_ASAP7_75t_L g372 ( .A(n_259), .B(n_373), .Y(n_372) );
OA21x2_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_267), .Y(n_259) );
OA21x2_ASAP7_75t_L g444 ( .A1(n_260), .A2(n_445), .B(n_451), .Y(n_444) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_260), .A2(n_474), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_260), .A2(n_487), .B(n_494), .Y(n_486) );
AND2x2_ASAP7_75t_L g374 ( .A(n_268), .B(n_313), .Y(n_374) );
AND2x2_ASAP7_75t_L g284 ( .A(n_269), .B(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_269), .B(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_SL g355 ( .A(n_271), .B(n_318), .Y(n_355) );
INVx1_ASAP7_75t_SL g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g361 ( .A(n_274), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g347 ( .A(n_275), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g412 ( .A(n_275), .B(n_357), .Y(n_412) );
INVx2_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
NAND4xp25_ASAP7_75t_SL g408 ( .A(n_277), .B(n_409), .C(n_410), .D(n_411), .Y(n_408) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_278), .B(n_342), .Y(n_377) );
OR2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
INVx1_ASAP7_75t_SL g414 ( .A(n_281), .Y(n_414) );
O2A1O1Ixp33_ASAP7_75t_SL g376 ( .A1(n_282), .A2(n_345), .B(n_349), .C(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g371 ( .A(n_284), .B(n_363), .Y(n_371) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_285), .Y(n_297) );
INVx1_ASAP7_75t_L g352 ( .A(n_285), .Y(n_352) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_286), .Y(n_329) );
AOI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .B(n_291), .C(n_293), .Y(n_287) );
AND2x2_ASAP7_75t_L g308 ( .A(n_288), .B(n_292), .Y(n_308) );
OAI322xp33_ASAP7_75t_SL g346 ( .A1(n_288), .A2(n_347), .A3(n_349), .B1(n_350), .B2(n_354), .C1(n_355), .C2(n_356), .Y(n_346) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g368 ( .A(n_290), .B(n_294), .Y(n_368) );
INVx1_ASAP7_75t_L g349 ( .A(n_292), .Y(n_349) );
INVx1_ASAP7_75t_SL g367 ( .A(n_294), .Y(n_367) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AOI222xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_308), .B2(n_309), .C1(n_310), .C2(n_716), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_301), .B(n_303), .Y(n_300) );
OAI322xp33_ASAP7_75t_L g389 ( .A1(n_301), .A2(n_363), .A3(n_368), .B1(n_390), .B2(n_391), .C1(n_393), .C2(n_394), .Y(n_389) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_302), .A2(n_316), .B1(n_340), .B2(n_344), .C(n_346), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
OAI222xp33_ASAP7_75t_L g319 ( .A1(n_307), .A2(n_320), .B1(n_322), .B2(n_323), .C1(n_324), .C2(n_327), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_309), .A2(n_316), .B1(n_386), .B2(n_387), .Y(n_385) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
AOI211xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B(n_319), .C(n_330), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g395 ( .A1(n_316), .A2(n_353), .B(n_396), .C(n_399), .Y(n_395) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g325 ( .A(n_317), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g388 ( .A(n_321), .Y(n_388) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_328), .B(n_353), .Y(n_382) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_333), .B(n_337), .Y(n_330) );
OAI221xp5_ASAP7_75t_SL g399 ( .A1(n_331), .A2(n_400), .B1(n_401), .B2(n_402), .C(n_403), .Y(n_399) );
INVxp33_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_335), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_342), .B(n_353), .Y(n_393) );
INVx2_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g404 ( .A(n_357), .B(n_363), .Y(n_404) );
AND4x1_ASAP7_75t_L g359 ( .A(n_360), .B(n_378), .C(n_395), .D(n_407), .Y(n_359) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OAI221xp5_ASAP7_75t_SL g364 ( .A1(n_365), .A2(n_366), .B1(n_368), .B2(n_369), .C(n_370), .Y(n_364) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_374), .B2(n_375), .Y(n_370) );
INVx1_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
INVx1_ASAP7_75t_SL g390 ( .A(n_375), .Y(n_390) );
NOR2xp33_ASAP7_75t_SL g378 ( .A(n_379), .B(n_389), .Y(n_378) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_391), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_398), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_413), .B1(n_414), .B2(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx2_ASAP7_75t_L g428 ( .A(n_421), .Y(n_428) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g429 ( .A1(n_425), .A2(n_430), .B(n_713), .Y(n_429) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_436), .B2(n_438), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx6_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g708 ( .A(n_437), .Y(n_708) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g709 ( .A(n_439), .Y(n_709) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_625), .Y(n_439) );
NOR4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_567), .C(n_597), .D(n_607), .Y(n_440) );
OAI211xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_482), .B(n_530), .C(n_557), .Y(n_441) );
OAI222xp33_ASAP7_75t_L g652 ( .A1(n_442), .A2(n_572), .B1(n_653), .B2(n_654), .C1(n_655), .C2(n_656), .Y(n_652) );
OR2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_461), .Y(n_442) );
AOI33xp33_ASAP7_75t_L g578 ( .A1(n_443), .A2(n_565), .A3(n_566), .B1(n_579), .B2(n_584), .B3(n_586), .Y(n_578) );
OAI211xp5_ASAP7_75t_SL g635 ( .A1(n_443), .A2(n_636), .B(n_638), .C(n_640), .Y(n_635) );
OR2x2_ASAP7_75t_L g651 ( .A(n_443), .B(n_637), .Y(n_651) );
INVx1_ASAP7_75t_L g684 ( .A(n_443), .Y(n_684) );
OR2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_452), .Y(n_443) );
INVx2_ASAP7_75t_L g561 ( .A(n_444), .Y(n_561) );
AND2x2_ASAP7_75t_L g577 ( .A(n_444), .B(n_473), .Y(n_577) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_444), .Y(n_612) );
AND2x2_ASAP7_75t_L g641 ( .A(n_444), .B(n_452), .Y(n_641) );
INVx2_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
BUFx3_ASAP7_75t_L g549 ( .A(n_452), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_452), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g560 ( .A(n_452), .B(n_561), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_452), .B(n_462), .Y(n_589) );
AND2x2_ASAP7_75t_L g658 ( .A(n_452), .B(n_592), .Y(n_658) );
INVx2_ASAP7_75t_SL g552 ( .A(n_461), .Y(n_552) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_462), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g594 ( .A(n_462), .Y(n_594) );
AND2x2_ASAP7_75t_L g605 ( .A(n_462), .B(n_561), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_462), .B(n_590), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_462), .B(n_592), .Y(n_637) );
AND2x2_ASAP7_75t_L g696 ( .A(n_462), .B(n_641), .Y(n_696) );
INVx4_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g566 ( .A(n_463), .B(n_473), .Y(n_566) );
AND2x2_ASAP7_75t_L g576 ( .A(n_463), .B(n_577), .Y(n_576) );
BUFx3_ASAP7_75t_L g598 ( .A(n_463), .Y(n_598) );
AND3x2_ASAP7_75t_L g657 ( .A(n_463), .B(n_658), .C(n_659), .Y(n_657) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
INVx1_ASAP7_75t_SL g592 ( .A(n_473), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_473), .B(n_541), .C(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_483), .B(n_513), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_483), .A2(n_576), .B(n_628), .C(n_630), .Y(n_627) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_485), .B(n_504), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_485), .B(n_634), .Y(n_633) );
INVx2_ASAP7_75t_SL g644 ( .A(n_485), .Y(n_644) );
AND2x2_ASAP7_75t_L g665 ( .A(n_485), .B(n_515), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_485), .B(n_574), .Y(n_693) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
AND2x2_ASAP7_75t_L g538 ( .A(n_486), .B(n_529), .Y(n_538) );
INVx2_ASAP7_75t_L g545 ( .A(n_486), .Y(n_545) );
AND2x2_ASAP7_75t_L g565 ( .A(n_486), .B(n_515), .Y(n_565) );
AND2x2_ASAP7_75t_L g615 ( .A(n_486), .B(n_504), .Y(n_615) );
INVx1_ASAP7_75t_L g619 ( .A(n_486), .Y(n_619) );
INVx2_ASAP7_75t_SL g529 ( .A(n_495), .Y(n_529) );
BUFx2_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
AND2x2_ASAP7_75t_L g682 ( .A(n_495), .B(n_504), .Y(n_682) );
INVx3_ASAP7_75t_SL g515 ( .A(n_504), .Y(n_515) );
AND2x2_ASAP7_75t_L g537 ( .A(n_504), .B(n_538), .Y(n_537) );
AND2x4_ASAP7_75t_L g544 ( .A(n_504), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g574 ( .A(n_504), .B(n_534), .Y(n_574) );
OR2x2_ASAP7_75t_L g583 ( .A(n_504), .B(n_529), .Y(n_583) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_504), .Y(n_601) );
AND2x2_ASAP7_75t_L g606 ( .A(n_504), .B(n_559), .Y(n_606) );
AND2x2_ASAP7_75t_L g634 ( .A(n_504), .B(n_517), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_504), .B(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g672 ( .A(n_504), .B(n_516), .Y(n_672) );
OR2x6_ASAP7_75t_L g504 ( .A(n_505), .B(n_511), .Y(n_504) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
AND2x2_ASAP7_75t_L g596 ( .A(n_515), .B(n_545), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_515), .B(n_538), .Y(n_624) );
AND2x2_ASAP7_75t_L g642 ( .A(n_515), .B(n_559), .Y(n_642) );
OR2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_529), .Y(n_516) );
AND2x2_ASAP7_75t_L g543 ( .A(n_517), .B(n_529), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_517), .B(n_572), .Y(n_571) );
BUFx3_ASAP7_75t_L g581 ( .A(n_517), .Y(n_581) );
OR2x2_ASAP7_75t_L g629 ( .A(n_517), .B(n_549), .Y(n_629) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .B(n_528), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_519), .A2(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g535 ( .A(n_521), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_528), .Y(n_536) );
AND2x2_ASAP7_75t_L g564 ( .A(n_529), .B(n_534), .Y(n_564) );
INVx1_ASAP7_75t_L g572 ( .A(n_529), .Y(n_572) );
AND2x2_ASAP7_75t_L g667 ( .A(n_529), .B(n_545), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_539), .B1(n_542), .B2(n_546), .C1(n_550), .C2(n_553), .Y(n_530) );
INVx1_ASAP7_75t_L g662 ( .A(n_531), .Y(n_662) );
AND2x2_ASAP7_75t_L g531 ( .A(n_532), .B(n_537), .Y(n_531) );
AND2x2_ASAP7_75t_L g558 ( .A(n_532), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g569 ( .A(n_532), .B(n_538), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_532), .B(n_560), .Y(n_585) );
OAI222xp33_ASAP7_75t_L g607 ( .A1(n_532), .A2(n_608), .B1(n_613), .B2(n_614), .C1(n_622), .C2(n_624), .Y(n_607) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g595 ( .A(n_534), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_534), .B(n_615), .Y(n_655) );
AND2x2_ASAP7_75t_L g666 ( .A(n_534), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g674 ( .A(n_537), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_539), .B(n_590), .Y(n_653) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_541), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g611 ( .A(n_541), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
INVx3_ASAP7_75t_L g556 ( .A(n_544), .Y(n_556) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_544), .A2(n_647), .B(n_650), .C(n_652), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_544), .B(n_581), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_544), .B(n_564), .Y(n_686) );
AND2x2_ASAP7_75t_L g559 ( .A(n_545), .B(n_555), .Y(n_559) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_549), .B(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g638 ( .A(n_549), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g677 ( .A(n_549), .B(n_577), .Y(n_677) );
INVx1_ASAP7_75t_L g689 ( .A(n_549), .Y(n_689) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_552), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
INVx1_ASAP7_75t_L g670 ( .A(n_555), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_560), .B(n_562), .C(n_566), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_558), .A2(n_588), .B1(n_603), .B2(n_606), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_559), .B(n_573), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_559), .B(n_581), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_560), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_SL g623 ( .A(n_560), .Y(n_623) );
AND2x2_ASAP7_75t_L g630 ( .A(n_560), .B(n_610), .Y(n_630) );
INVx2_ASAP7_75t_L g591 ( .A(n_561), .Y(n_591) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NOR4xp25_ASAP7_75t_L g568 ( .A(n_565), .B(n_569), .C(n_570), .D(n_573), .Y(n_568) );
INVx1_ASAP7_75t_SL g639 ( .A(n_566), .Y(n_639) );
AND2x2_ASAP7_75t_L g683 ( .A(n_566), .B(n_684), .Y(n_683) );
OAI211xp5_ASAP7_75t_SL g567 ( .A1(n_568), .A2(n_575), .B(n_578), .C(n_587), .Y(n_567) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_574), .B(n_644), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_576), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_694) );
INVx1_ASAP7_75t_SL g649 ( .A(n_577), .Y(n_649) );
AND2x2_ASAP7_75t_L g688 ( .A(n_577), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_581), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_585), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_586), .B(n_611), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_593), .B(n_595), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g663 ( .A(n_590), .Y(n_663) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g691 ( .A(n_591), .Y(n_691) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_592), .Y(n_618) );
OAI21xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_602), .Y(n_597) );
CKINVDCx16_ASAP7_75t_R g610 ( .A(n_598), .Y(n_610) );
OR2x2_ASAP7_75t_L g648 ( .A(n_598), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_601), .A2(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_605), .A2(n_632), .B1(n_635), .B2(n_642), .C(n_643), .Y(n_631) );
INVx1_ASAP7_75t_SL g675 ( .A(n_606), .Y(n_675) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g622 ( .A(n_610), .B(n_623), .Y(n_622) );
INVxp67_ASAP7_75t_L g659 ( .A(n_612), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_616), .B1(n_619), .B2(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g654 ( .A(n_615), .Y(n_654) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_618), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NOR4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_660), .C(n_673), .D(n_685), .Y(n_625) );
NAND3xp33_ASAP7_75t_SL g626 ( .A(n_627), .B(n_631), .C(n_646), .Y(n_626) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_629), .B(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_636), .B(n_641), .Y(n_645) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_648), .A2(n_674), .B1(n_675), .B2(n_676), .C(n_678), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_650), .A2(n_665), .B(n_666), .C(n_668), .Y(n_664) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_651), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_668) );
INVx2_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B(n_663), .C(n_664), .Y(n_660) );
INVx1_ASAP7_75t_L g679 ( .A(n_672), .Y(n_679) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g678 ( .A1(n_679), .A2(n_680), .B(n_683), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI221xp5_ASAP7_75t_SL g685 ( .A1(n_686), .A2(n_687), .B1(n_690), .B2(n_692), .C(n_694), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
INVx3_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
endmodule