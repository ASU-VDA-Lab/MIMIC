module fake_aes_11290_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_8;
wire n_10;
wire n_7;
INVx1_ASAP7_75t_L g3 ( .A(n_0), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
BUFx10_ASAP7_75t_L g5 ( .A(n_0), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
AND2x4_ASAP7_75t_L g7 ( .A(n_4), .B(n_0), .Y(n_7) );
OAI21x1_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_1), .B(n_2), .Y(n_8) );
BUFx2_ASAP7_75t_L g9 ( .A(n_8), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
AOI22xp5_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_7), .B1(n_5), .B2(n_8), .Y(n_11) );
OAI221xp5_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_6), .B1(n_5), .B2(n_7), .C(n_1), .Y(n_12) );
OAI22x1_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_7), .B1(n_1), .B2(n_6), .Y(n_13) );
endmodule