module fake_jpeg_21585_n_324 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_14),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_34),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_14),
.B1(n_19),
.B2(n_18),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_38),
.A2(n_30),
.B1(n_27),
.B2(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_41),
.Y(n_50)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_49),
.A2(n_64),
.B1(n_40),
.B2(n_36),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_44),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_60),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_25),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_40),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_24),
.Y(n_69)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_65),
.A2(n_62),
.B1(n_53),
.B2(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_72),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_36),
.B1(n_45),
.B2(n_46),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_14),
.B1(n_60),
.B2(n_52),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_35),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_59),
.A2(n_37),
.B1(n_39),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_76),
.B1(n_53),
.B2(n_45),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_19),
.B1(n_18),
.B2(n_43),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_58),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_84),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_48),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_36),
.B(n_31),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_90),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_105),
.B(n_78),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_64),
.B1(n_49),
.B2(n_45),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_91),
.A2(n_97),
.B1(n_102),
.B2(n_80),
.Y(n_118)
);

OAI21x1_ASAP7_75t_R g92 ( 
.A1(n_71),
.A2(n_47),
.B(n_12),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_33),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_104),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_66),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_65),
.A2(n_61),
.B1(n_14),
.B2(n_29),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_103),
.A2(n_60),
.B1(n_52),
.B2(n_12),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_31),
.C(n_26),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_20),
.B(n_16),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_89),
.B(n_101),
.Y(n_111)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_70),
.A3(n_72),
.B1(n_84),
.B2(n_77),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_108),
.A2(n_111),
.B(n_126),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_69),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_110),
.B(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_69),
.Y(n_116)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_77),
.A3(n_68),
.B1(n_82),
.B2(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_119),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_118),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_172)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_92),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_127),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_82),
.B1(n_80),
.B2(n_76),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_121),
.A2(n_137),
.B1(n_112),
.B2(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_79),
.C(n_82),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_100),
.C(n_95),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_75),
.B(n_15),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_79),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_31),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_63),
.Y(n_164)
);

OR2x2_ASAP7_75t_SL g129 ( 
.A(n_85),
.B(n_78),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_10),
.C(n_22),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_91),
.A2(n_80),
.B1(n_19),
.B2(n_18),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_19),
.B1(n_18),
.B2(n_16),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_18),
.B1(n_15),
.B2(n_16),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_15),
.B1(n_16),
.B2(n_12),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_137),
.B1(n_98),
.B2(n_97),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_63),
.B(n_20),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_17),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_133),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_140),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_139),
.A2(n_145),
.B1(n_148),
.B2(n_171),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_94),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_142),
.B(n_149),
.Y(n_196)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_143),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_109),
.A2(n_86),
.B1(n_92),
.B2(n_105),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_20),
.B1(n_10),
.B2(n_2),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_147),
.C(n_152),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_106),
.C(n_103),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_112),
.A2(n_103),
.B1(n_106),
.B2(n_15),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_114),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_79),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_23),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_79),
.C(n_57),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_63),
.A3(n_26),
.B1(n_32),
.B2(n_52),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_154),
.A2(n_159),
.B(n_136),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_32),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_155),
.B(n_157),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_63),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_123),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_164),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_116),
.B(n_57),
.C(n_21),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_165),
.B(n_166),
.C(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_115),
.B(n_113),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_60),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_170),
.A2(n_130),
.B(n_118),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_120),
.A2(n_20),
.B1(n_10),
.B2(n_57),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_113),
.B(n_126),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_131),
.C(n_132),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_176),
.B(n_186),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_198),
.B(n_202),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_21),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_135),
.C(n_57),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_188),
.A2(n_192),
.B1(n_193),
.B2(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_156),
.A2(n_23),
.B1(n_21),
.B2(n_13),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_201),
.B1(n_184),
.B2(n_190),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_166),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_192)
);

OAI22x1_ASAP7_75t_SL g193 ( 
.A1(n_153),
.A2(n_22),
.B1(n_17),
.B2(n_10),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_197),
.Y(n_204)
);

AND2x4_ASAP7_75t_SL g198 ( 
.A(n_141),
.B(n_22),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_163),
.B(n_21),
.C(n_13),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_169),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_22),
.B(n_11),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_164),
.C(n_173),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_199),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_147),
.B(n_146),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_174),
.B(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_207),
.A2(n_226),
.B1(n_0),
.B2(n_3),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_186),
.A2(n_165),
.B1(n_157),
.B2(n_155),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_217),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_183),
.B(n_185),
.Y(n_217)
);

AOI221xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_139),
.B1(n_162),
.B2(n_158),
.C(n_11),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_225),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_219),
.B(n_221),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_195),
.Y(n_227)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_174),
.C(n_178),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_237),
.C(n_241),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_232),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_178),
.C(n_200),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_194),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_242),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_223),
.A2(n_177),
.B1(n_194),
.B2(n_198),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_214),
.B1(n_207),
.B2(n_222),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_198),
.C(n_192),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_21),
.Y(n_242)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_245),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_21),
.C(n_13),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_210),
.C(n_221),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_3),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_228),
.B(n_211),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_253),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_230),
.B(n_204),
.Y(n_255)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_224),
.B1(n_216),
.B2(n_226),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_258),
.B1(n_259),
.B2(n_220),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_215),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_261),
.Y(n_272)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_262),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_241),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_265),
.Y(n_278)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_4),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_220),
.B1(n_236),
.B2(n_204),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_268),
.A2(n_271),
.B1(n_263),
.B2(n_259),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_257),
.B(n_232),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_250),
.A2(n_242),
.B1(n_233),
.B2(n_238),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_239),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_276),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_260),
.A2(n_229),
.B(n_240),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_231),
.B(n_258),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_262),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_237),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_251),
.C(n_252),
.Y(n_286)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

FAx1_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_233),
.CI(n_222),
.CON(n_282),
.SN(n_282)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_288),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_7),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_3),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_3),
.Y(n_288)
);

AND2x4_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_4),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_290),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_4),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_269),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_291),
.B(n_292),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_267),
.B1(n_277),
.B2(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_301),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_4),
.C(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_298),
.B(n_300),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_5),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_7),
.B(n_8),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_302),
.B(n_290),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_7),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_307),
.B(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_8),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_8),
.C(n_9),
.Y(n_312)
);

OAI21x1_ASAP7_75t_SL g314 ( 
.A1(n_312),
.A2(n_299),
.B(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_314),
.B(n_310),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_315),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_SL g318 ( 
.A(n_313),
.B(n_305),
.C(n_300),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_316),
.C(n_311),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_304),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_8),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_9),
.B(n_317),
.Y(n_324)
);


endmodule