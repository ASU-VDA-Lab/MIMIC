module fake_jpeg_10577_n_171 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_11),
.B(n_1),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_33),
.B(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_21),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_25),
.B1(n_17),
.B2(n_21),
.Y(n_52)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NAND2x1p5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_24),
.Y(n_45)
);

XNOR2x1_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_33),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_28),
.B1(n_23),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_34),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_30),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_28),
.B1(n_20),
.B2(n_18),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_52),
.B1(n_56),
.B2(n_29),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_14),
.B1(n_18),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_38),
.B1(n_31),
.B2(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_53),
.B(n_19),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_31),
.B1(n_17),
.B2(n_15),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_59),
.B(n_26),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_19),
.B1(n_16),
.B2(n_41),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_29),
.A3(n_36),
.B1(n_34),
.B2(n_32),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_42),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_62),
.A2(n_26),
.B1(n_24),
.B2(n_16),
.Y(n_92)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_65),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_15),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_70),
.Y(n_88)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_30),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_64),
.A2(n_43),
.B1(n_31),
.B2(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_77),
.B1(n_83),
.B2(n_32),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_35),
.B(n_51),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_87),
.B(n_89),
.C(n_26),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_67),
.A2(n_35),
.B1(n_41),
.B2(n_39),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_55),
.B1(n_26),
.B2(n_27),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_69),
.B(n_73),
.C(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_82),
.A2(n_92),
.B1(n_66),
.B2(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_41),
.B1(n_39),
.B2(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_59),
.A2(n_51),
.B(n_39),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_103),
.Y(n_110)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_91),
.Y(n_94)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_97),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_70),
.C(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_51),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_102),
.B1(n_108),
.B2(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_55),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_13),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_81),
.B(n_13),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_0),
.Y(n_122)
);

XOR2x1_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_89),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_88),
.C(n_85),
.Y(n_112)
);

OA21x2_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_99),
.B(n_82),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_83),
.B(n_88),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_113),
.A2(n_114),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_95),
.A2(n_76),
.B(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_97),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_131),
.C(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_100),
.B1(n_108),
.B2(n_95),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_130),
.B(n_94),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_106),
.B(n_99),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_113),
.Y(n_131)
);

OAI321xp33_ASAP7_75t_L g140 ( 
.A1(n_133),
.A2(n_120),
.A3(n_116),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_86),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_84),
.B(n_77),
.C(n_102),
.D(n_39),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_110),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_141),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_132),
.B(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_128),
.A2(n_127),
.B1(n_118),
.B2(n_130),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_139),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_140),
.A2(n_142),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_134),
.B(n_111),
.Y(n_141)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_111),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_143),
.A2(n_135),
.B1(n_129),
.B2(n_131),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_94),
.C(n_91),
.Y(n_145)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_145),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_143),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_153),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_144),
.B(n_6),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_148),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_144),
.C(n_7),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_5),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_8),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_158),
.B(n_148),
.C(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_163),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_164),
.B(n_156),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_165),
.A2(n_160),
.B(n_10),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_166),
.B(n_11),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);


endmodule