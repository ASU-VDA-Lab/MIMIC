module fake_jpeg_1498_n_227 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_227);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_227;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_220;
wire n_137;
wire n_31;
wire n_207;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_10),
.B(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_39),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_58),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_21),
.B(n_13),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_45),
.B(n_55),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_48),
.Y(n_86)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_49),
.B(n_65),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx6p67_ASAP7_75t_R g91 ( 
.A(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_1),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_28),
.B(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_64),
.Y(n_90)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_15),
.B(n_2),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_34),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_93),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_30),
.B(n_19),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_79),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_19),
.B1(n_34),
.B2(n_32),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_87),
.A2(n_97),
.B1(n_29),
.B2(n_8),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_32),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_57),
.A2(n_18),
.B1(n_23),
.B2(n_22),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_87),
.B1(n_80),
.B2(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_18),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_99),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_19),
.B1(n_27),
.B2(n_23),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_42),
.B(n_36),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_16),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_4),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_56),
.B(n_16),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_27),
.B1(n_29),
.B2(n_7),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_59),
.B1(n_29),
.B2(n_7),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_47),
.B(n_4),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_38),
.B(n_29),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_106),
.B(n_54),
.Y(n_111)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_130),
.B1(n_105),
.B2(n_80),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_113),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_124),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_4),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_114),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_5),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_5),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_71),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_11),
.B1(n_29),
.B2(n_91),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_79),
.A2(n_11),
.B1(n_93),
.B2(n_76),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_11),
.B1(n_91),
.B2(n_102),
.Y(n_123)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_126),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_86),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_77),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_134),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_89),
.A2(n_74),
.B1(n_87),
.B2(n_102),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_104),
.B(n_70),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_131),
.B(n_89),
.Y(n_140)
);

NOR2x1_ASAP7_75t_R g133 ( 
.A(n_87),
.B(n_106),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_82),
.Y(n_149)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_73),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_138),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_75),
.B1(n_105),
.B2(n_95),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_151),
.B(n_152),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_118),
.A2(n_82),
.B(n_95),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_122),
.A2(n_111),
.B(n_130),
.Y(n_152)
);

AOI22x1_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_72),
.B1(n_107),
.B2(n_81),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_153),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_111),
.A2(n_108),
.B(n_73),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_160),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_139),
.Y(n_170)
);

O2A1O1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_128),
.A2(n_72),
.B(n_81),
.C(n_85),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_109),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_165),
.B(n_174),
.Y(n_181)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_170),
.Y(n_187)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_138),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_169),
.C(n_148),
.D(n_114),
.Y(n_188)
);

O2A1O1Ixp5_ASAP7_75t_L g169 ( 
.A1(n_140),
.A2(n_139),
.B(n_131),
.C(n_115),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_143),
.B1(n_150),
.B2(n_141),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_128),
.C(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.C(n_176),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_112),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_150),
.B(n_110),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_135),
.C(n_119),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_182),
.Y(n_194)
);

NOR3xp33_ASAP7_75t_SL g182 ( 
.A(n_173),
.B(n_158),
.C(n_146),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_161),
.B1(n_146),
.B2(n_144),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_184),
.B1(n_191),
.B2(n_167),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_162),
.B1(n_147),
.B2(n_153),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_153),
.B(n_160),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

AOI211xp5_ASAP7_75t_SL g186 ( 
.A1(n_178),
.A2(n_160),
.B(n_162),
.C(n_148),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_177),
.B(n_167),
.Y(n_198)
);

OAI322xp33_ASAP7_75t_L g196 ( 
.A1(n_188),
.A2(n_172),
.A3(n_177),
.B1(n_156),
.B2(n_166),
.C1(n_163),
.C2(n_176),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_154),
.B(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_190),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_168),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_182),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

XOR2x2_ASAP7_75t_L g204 ( 
.A(n_196),
.B(n_188),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_198),
.A2(n_181),
.B(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_181),
.B1(n_179),
.B2(n_185),
.Y(n_202)
);

AO221x1_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_183),
.B1(n_124),
.B2(n_187),
.C(n_125),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_202),
.A2(n_207),
.B1(n_205),
.B2(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_180),
.Y(n_203)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_192),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_208),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_205),
.A2(n_197),
.B(n_193),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_189),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_209),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_193),
.B1(n_208),
.B2(n_206),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_197),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_212),
.B(n_204),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_155),
.B(n_159),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_218),
.A2(n_219),
.B(n_209),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_155),
.C(n_125),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_215),
.B(n_211),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_221),
.A2(n_222),
.B(n_223),
.Y(n_225)
);

AOI322xp5_ASAP7_75t_L g223 ( 
.A1(n_215),
.A2(n_159),
.A3(n_145),
.B1(n_124),
.B2(n_132),
.C1(n_71),
.C2(n_136),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_220),
.A2(n_145),
.B(n_132),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_137),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);


endmodule