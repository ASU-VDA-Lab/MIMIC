module fake_jpeg_5898_n_332 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_15),
.B(n_0),
.Y(n_37)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_37),
.B(n_10),
.Y(n_101)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_39),
.B(n_45),
.Y(n_69)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_14),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_48),
.B(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g103 ( 
.A(n_50),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_36),
.B1(n_34),
.B2(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_32),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_62),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_55),
.A2(n_101),
.B(n_22),
.C(n_14),
.Y(n_132)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_26),
.B1(n_33),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_57),
.A2(n_68),
.B1(n_75),
.B2(n_22),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_60),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_25),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_25),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_66),
.Y(n_128)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_72),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_15),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_51),
.A2(n_46),
.B1(n_53),
.B2(n_38),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_17),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_87),
.Y(n_110)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_73),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_44),
.A2(n_26),
.B1(n_21),
.B2(n_36),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_41),
.B(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_23),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_49),
.B(n_29),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_29),
.Y(n_88)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_31),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_92),
.C(n_30),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_95),
.Y(n_135)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_28),
.C(n_31),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_45),
.B(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_45),
.B(n_18),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_81),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_108),
.B(n_103),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_32),
.B1(n_19),
.B2(n_30),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_115),
.A2(n_121),
.B1(n_100),
.B2(n_102),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_30),
.B(n_32),
.C(n_19),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_116),
.A2(n_79),
.B1(n_85),
.B2(n_94),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_30),
.B1(n_32),
.B2(n_19),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_119),
.A2(n_134),
.B1(n_61),
.B2(n_76),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_56),
.A2(n_30),
.B1(n_22),
.B2(n_20),
.Y(n_121)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_30),
.B1(n_22),
.B2(n_20),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_127),
.B(n_130),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_89),
.A2(n_22),
.B(n_1),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_54),
.A2(n_22),
.B(n_1),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_132),
.B(n_92),
.Y(n_145)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_136),
.B(n_137),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g137 ( 
.A(n_121),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_130),
.A2(n_62),
.B(n_63),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_150),
.B(n_107),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_142),
.A2(n_129),
.B1(n_65),
.B2(n_4),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_72),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_145),
.B(n_126),
.Y(n_187)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_146),
.B(n_147),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_121),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_103),
.C(n_82),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_156),
.C(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_91),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_127),
.A2(n_71),
.B(n_60),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_90),
.C(n_64),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_151),
.B(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_58),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_70),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_111),
.Y(n_197)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_155),
.Y(n_195)
);

INVx11_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

OA22x2_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_94),
.B1(n_85),
.B2(n_80),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_167),
.B(n_124),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_110),
.B(n_99),
.C(n_97),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_117),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_163),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_161),
.A2(n_113),
.B1(n_129),
.B2(n_109),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_162),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_69),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_100),
.Y(n_165)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_86),
.B(n_59),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_157),
.B1(n_109),
.B2(n_136),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_169),
.B(n_173),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_112),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_170),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_125),
.B(n_61),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_0),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_135),
.B1(n_105),
.B2(n_123),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_174),
.A2(n_178),
.B1(n_202),
.B2(n_65),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_166),
.A2(n_123),
.B1(n_133),
.B2(n_112),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_150),
.B(n_139),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_194),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_187),
.A2(n_192),
.B(n_153),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_139),
.B1(n_154),
.B2(n_137),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_159),
.C(n_148),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_1),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_152),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_205),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_144),
.B(n_2),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_164),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_158),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_2),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_173),
.Y(n_222)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_157),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_210),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_214),
.A2(n_224),
.B(n_225),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_210),
.A2(n_142),
.B1(n_145),
.B2(n_169),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_228),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_201),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_205),
.B(n_170),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_227),
.C(n_237),
.Y(n_253)
);

NAND2xp33_ASAP7_75t_SL g224 ( 
.A(n_192),
.B(n_156),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_156),
.Y(n_226)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_189),
.A2(n_147),
.B(n_137),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_189),
.B(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_229),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_211),
.A2(n_208),
.B1(n_193),
.B2(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_232),
.B1(n_235),
.B2(n_181),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_179),
.A2(n_161),
.B(n_4),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_8),
.C(n_11),
.Y(n_236)
);

OAI322xp33_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_209),
.A3(n_206),
.B1(n_203),
.B2(n_174),
.C1(n_9),
.C2(n_12),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_238),
.B(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_190),
.B(n_8),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_188),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_241),
.B(n_252),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

NOR3xp33_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_260),
.C(n_262),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_238),
.A2(n_204),
.B1(n_186),
.B2(n_176),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_212),
.B(n_219),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_233),
.B1(n_218),
.B2(n_214),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_255),
.B1(n_258),
.B2(n_213),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_229),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_237),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_257),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_181),
.C(n_191),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_232),
.A2(n_187),
.B1(n_199),
.B2(n_184),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_202),
.Y(n_261)
);

AOI321xp33_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_224),
.A3(n_227),
.B1(n_217),
.B2(n_222),
.C(n_216),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_240),
.A2(n_230),
.B1(n_215),
.B2(n_227),
.Y(n_265)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_250),
.A2(n_233),
.B1(n_242),
.B2(n_244),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_248),
.A2(n_212),
.B1(n_220),
.B2(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_278),
.C(n_257),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_247),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_271),
.B(n_273),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_234),
.B1(n_217),
.B2(n_180),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_274),
.C(n_277),
.Y(n_281)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_250),
.A2(n_234),
.B(n_239),
.Y(n_274)
);

OA21x2_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_176),
.B(n_228),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_246),
.B(n_245),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_244),
.A2(n_196),
.B1(n_236),
.B2(n_177),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_245),
.A2(n_196),
.B1(n_177),
.B2(n_175),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_241),
.C(n_253),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_286),
.C(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_285),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_253),
.C(n_256),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_252),
.C(n_254),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_274),
.B(n_267),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_262),
.C(n_243),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_263),
.C(n_266),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_280),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_299),
.C(n_281),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_264),
.C(n_272),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_290),
.C(n_281),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_300),
.A2(n_301),
.B(n_305),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_282),
.A2(n_265),
.B(n_251),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_283),
.A2(n_277),
.B1(n_278),
.B2(n_251),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_294),
.B1(n_293),
.B2(n_198),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_198),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_307),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_311),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_175),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_304),
.B(n_231),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.Y(n_321)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_301),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_297),
.C(n_298),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_296),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_299),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_319),
.B(n_322),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_303),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_309),
.B(n_306),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_308),
.Y(n_324)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_321),
.B(n_317),
.C(n_318),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_320),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_317),
.B(n_302),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_328),
.B(n_327),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_329),
.C(n_231),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_183),
.Y(n_332)
);


endmodule