module fake_aes_8222_n_1600 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1600);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1600;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1571;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_1594;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1527;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_1528;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1598;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_1536;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_1597;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1573;
wire n_1580;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_1595;
wire n_610;
wire n_771;
wire n_1561;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1525;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_1569;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1547;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1582;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_1551;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1522;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_994;
wire n_930;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1590;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_1533;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_1563;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1542;
wire n_1311;
wire n_1558;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_1557;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_1564;
wire n_1521;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_1539;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_1543;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_1581;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1537;
wire n_634;
wire n_1271;
wire n_1520;
wire n_696;
wire n_1203;
wire n_1546;
wire n_1524;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_1540;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_1593;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1562;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1541;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_1553;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1432;
wire n_1315;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1529;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1577;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_1583;
wire n_606;
wire n_1585;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_1586;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1566;
wire n_1236;
wire n_791;
wire n_707;
wire n_1599;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1559;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_1530;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_1554;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1572;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_1579;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_1575;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_1526;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_1576;
wire n_832;
wire n_996;
wire n_1578;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1517;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1565;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1552;
wire n_1170;
wire n_1523;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_1550;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1587;
wire n_1489;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1592;
wire n_1168;
wire n_1574;
wire n_458;
wire n_1084;
wire n_618;
wire n_1596;
wire n_470;
wire n_1085;
wire n_1538;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1555;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_1570;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_1544;
wire n_743;
wire n_757;
wire n_1568;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1545;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_1534;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_1518;
wire n_945;
wire n_554;
wire n_726;
wire n_1519;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_1589;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_1560;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_1532;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1291;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1535;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1567;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1591;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1549;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_1531;
wire n_371;
wire n_1548;
wire n_1584;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_1588;
wire n_480;
wire n_453;
wire n_833;
wire n_1556;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1442;
INVx2_ASAP7_75t_L g347 ( .A(n_101), .Y(n_347) );
CKINVDCx5p33_ASAP7_75t_R g348 ( .A(n_130), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_196), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_87), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_234), .B(n_161), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_77), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_319), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_310), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_276), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_38), .Y(n_356) );
NOR2xp67_ASAP7_75t_L g357 ( .A(n_15), .B(n_126), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_339), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_88), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_244), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_162), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_141), .Y(n_362) );
BUFx5_ASAP7_75t_L g363 ( .A(n_113), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_100), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_118), .Y(n_365) );
CKINVDCx5p33_ASAP7_75t_R g366 ( .A(n_4), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_246), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_166), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_201), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_284), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_336), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_249), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_148), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_262), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_150), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_82), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_82), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_329), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_184), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_254), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_156), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_90), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_235), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_321), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_306), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_239), .Y(n_386) );
CKINVDCx20_ASAP7_75t_R g387 ( .A(n_96), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_241), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_39), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_193), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_183), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_314), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_189), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_130), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_221), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_119), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_25), .Y(n_397) );
CKINVDCx5p33_ASAP7_75t_R g398 ( .A(n_222), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_121), .Y(n_399) );
NOR2xp67_ASAP7_75t_L g400 ( .A(n_121), .B(n_93), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_190), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_281), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_226), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g404 ( .A(n_111), .Y(n_404) );
BUFx3_ASAP7_75t_L g405 ( .A(n_265), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_73), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_182), .Y(n_407) );
CKINVDCx5p33_ASAP7_75t_R g408 ( .A(n_128), .Y(n_408) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_143), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_75), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_167), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_258), .Y(n_412) );
BUFx3_ASAP7_75t_L g413 ( .A(n_188), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_106), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_299), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_259), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_297), .Y(n_417) );
INVxp67_ASAP7_75t_SL g418 ( .A(n_44), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_126), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_287), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_194), .Y(n_421) );
CKINVDCx5p33_ASAP7_75t_R g422 ( .A(n_61), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_334), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_136), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_0), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_209), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_59), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_275), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_158), .Y(n_429) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_267), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_170), .Y(n_431) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_253), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_342), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_119), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_169), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_294), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_94), .Y(n_437) );
INVx3_ASAP7_75t_L g438 ( .A(n_325), .Y(n_438) );
NOR2xp67_ASAP7_75t_L g439 ( .A(n_315), .B(n_327), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_134), .Y(n_440) );
INVxp67_ASAP7_75t_L g441 ( .A(n_142), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_174), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g443 ( .A(n_279), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_61), .Y(n_444) );
INVxp33_ASAP7_75t_L g445 ( .A(n_269), .Y(n_445) );
BUFx2_ASAP7_75t_L g446 ( .A(n_318), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_125), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_263), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_128), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_144), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_22), .Y(n_451) );
BUFx3_ASAP7_75t_L g452 ( .A(n_290), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_286), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_323), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_213), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_317), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_331), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_346), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_125), .Y(n_459) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_65), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_309), .Y(n_461) );
INVxp67_ASAP7_75t_L g462 ( .A(n_187), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_90), .Y(n_463) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_6), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_197), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_177), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_289), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_192), .Y(n_468) );
INVxp67_ASAP7_75t_SL g469 ( .A(n_165), .Y(n_469) );
CKINVDCx14_ASAP7_75t_R g470 ( .A(n_178), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_153), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_231), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_322), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_312), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_40), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_114), .Y(n_476) );
NOR2xp67_ASAP7_75t_L g477 ( .A(n_77), .B(n_145), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_4), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_207), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_146), .Y(n_480) );
CKINVDCx5p33_ASAP7_75t_R g481 ( .A(n_271), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_36), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_62), .Y(n_483) );
INVxp67_ASAP7_75t_SL g484 ( .A(n_320), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g485 ( .A(n_277), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_123), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_203), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_343), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_307), .Y(n_489) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_288), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_311), .Y(n_491) );
INVxp67_ASAP7_75t_SL g492 ( .A(n_120), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_204), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_27), .Y(n_494) );
HB1xp67_ASAP7_75t_SL g495 ( .A(n_29), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_224), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_304), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_313), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_7), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_283), .Y(n_500) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_316), .Y(n_501) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_131), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_78), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_21), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_171), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_285), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_139), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_232), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_1), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_46), .Y(n_510) );
CKINVDCx16_ASAP7_75t_R g511 ( .A(n_252), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_41), .Y(n_512) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_256), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_301), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_160), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_131), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_55), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_335), .Y(n_518) );
NOR2xp67_ASAP7_75t_L g519 ( .A(n_260), .B(n_15), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_37), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_238), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_75), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g523 ( .A(n_39), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_185), .Y(n_524) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_9), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_270), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_24), .Y(n_527) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_245), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_168), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_300), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_57), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_293), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_26), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_84), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_36), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_38), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_157), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_92), .Y(n_538) );
CKINVDCx5p33_ASAP7_75t_R g539 ( .A(n_110), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_261), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g541 ( .A(n_278), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_326), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_445), .B(n_0), .Y(n_543) );
INVx3_ASAP7_75t_L g544 ( .A(n_363), .Y(n_544) );
CKINVDCx11_ASAP7_75t_R g545 ( .A(n_356), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_449), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_438), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_438), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_368), .B(n_1), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_438), .Y(n_550) );
NOR2xp33_ASAP7_75t_SL g551 ( .A(n_511), .B(n_137), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_414), .Y(n_552) );
INVx5_ASAP7_75t_L g553 ( .A(n_455), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_363), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_404), .A2(n_5), .B1(n_2), .B2(n_3), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_362), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_455), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_455), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_446), .B(n_2), .Y(n_559) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_455), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_501), .Y(n_563) );
INVx4_ASAP7_75t_L g564 ( .A(n_405), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_501), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_539), .A2(n_6), .B1(n_3), .B2(n_5), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_363), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_495), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_568) );
INVx3_ASAP7_75t_L g569 ( .A(n_363), .Y(n_569) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_528), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_363), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_528), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
NOR2xp33_ASAP7_75t_SL g574 ( .A(n_361), .B(n_345), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_350), .B(n_8), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_363), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_528), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_352), .B(n_10), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_363), .Y(n_579) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_349), .A2(n_140), .B(n_138), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_347), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_349), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_419), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_414), .Y(n_584) );
AND2x2_ASAP7_75t_SL g585 ( .A(n_353), .B(n_344), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_552), .B(n_445), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_552), .B(n_539), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_546), .B(n_433), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_544), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_560), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_543), .B(n_361), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_544), .Y(n_592) );
OR2x6_ASAP7_75t_L g593 ( .A(n_568), .B(n_357), .Y(n_593) );
AND2x6_ASAP7_75t_L g594 ( .A(n_543), .B(n_405), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_544), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_544), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_569), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_547), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_543), .B(n_383), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_569), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_564), .B(n_541), .Y(n_602) );
AND3x2_ASAP7_75t_L g603 ( .A(n_546), .B(n_509), .C(n_460), .Y(n_603) );
INVx4_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_576), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_576), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_576), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_576), .Y(n_608) );
INVx6_ASAP7_75t_L g609 ( .A(n_564), .Y(n_609) );
INVx3_ASAP7_75t_L g610 ( .A(n_547), .Y(n_610) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_585), .B(n_541), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_564), .B(n_542), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_564), .B(n_542), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_554), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_560), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_583), .B(n_441), .Y(n_616) );
INVx2_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_584), .B(n_470), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_585), .B(n_456), .Y(n_619) );
BUFx3_ASAP7_75t_L g620 ( .A(n_584), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_551), .B(n_462), .Y(n_621) );
NAND2xp33_ASAP7_75t_L g622 ( .A(n_547), .B(n_358), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_548), .B(n_535), .Y(n_623) );
OR2x6_ASAP7_75t_L g624 ( .A(n_568), .B(n_400), .Y(n_624) );
NAND2xp33_ASAP7_75t_L g625 ( .A(n_548), .B(n_360), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
BUFx2_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_627), .B(n_556), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_623), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_620), .Y(n_630) );
NOR2xp33_ASAP7_75t_L g631 ( .A(n_586), .B(n_559), .Y(n_631) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_620), .Y(n_632) );
OAI22xp5_ASAP7_75t_SL g633 ( .A1(n_593), .A2(n_377), .B1(n_387), .B2(n_356), .Y(n_633) );
CKINVDCx6p67_ASAP7_75t_R g634 ( .A(n_593), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_627), .Y(n_635) );
INVxp67_ASAP7_75t_L g636 ( .A(n_591), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_593), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_600), .Y(n_638) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_616), .A2(n_555), .B1(n_575), .B2(n_578), .C(n_559), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_587), .B(n_549), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_588), .B(n_584), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_594), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_619), .B(n_575), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_594), .B(n_578), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_623), .Y(n_645) );
NAND2x1p5_ASAP7_75t_L g646 ( .A(n_621), .B(n_623), .Y(n_646) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_620), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_593), .B(n_551), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_623), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_593), .B(n_348), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_594), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_624), .B(n_555), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g653 ( .A(n_611), .B(n_574), .C(n_566), .Y(n_653) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_614), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_599), .Y(n_655) );
INVx4_ASAP7_75t_L g656 ( .A(n_594), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_594), .B(n_548), .Y(n_657) );
INVx5_ASAP7_75t_L g658 ( .A(n_594), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_594), .A2(n_567), .B1(n_579), .B2(n_571), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_614), .A2(n_581), .B1(n_492), .B2(n_478), .C(n_418), .Y(n_660) );
AOI22x1_ASAP7_75t_SL g661 ( .A1(n_624), .A2(n_387), .B1(n_399), .B2(n_377), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
AND2x6_ASAP7_75t_SL g663 ( .A(n_624), .B(n_545), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_602), .B(n_581), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_599), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_624), .A2(n_571), .B1(n_579), .B2(n_582), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_612), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_610), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_603), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_613), .B(n_393), .Y(n_670) );
INVxp67_ASAP7_75t_L g671 ( .A(n_618), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g672 ( .A1(n_624), .A2(n_582), .B(n_359), .C(n_382), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_622), .A2(n_362), .B1(n_409), .B2(n_379), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_610), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g675 ( .A(n_610), .B(n_550), .Y(n_675) );
NAND2x1p5_ASAP7_75t_L g676 ( .A(n_610), .B(n_566), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_601), .B(n_604), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_626), .A2(n_409), .B1(n_420), .B2(n_379), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_601), .B(n_550), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_626), .A2(n_582), .B1(n_364), .B2(n_396), .Y(n_680) );
NAND3xp33_ASAP7_75t_SL g681 ( .A(n_592), .B(n_366), .C(n_365), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_592), .Y(n_682) );
NOR2xp33_ASAP7_75t_SL g683 ( .A(n_601), .B(n_420), .Y(n_683) );
INVx2_ASAP7_75t_SL g684 ( .A(n_609), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_601), .B(n_354), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_617), .A2(n_389), .B1(n_406), .B2(n_397), .Y(n_686) );
AOI22xp33_ASAP7_75t_SL g687 ( .A1(n_625), .A2(n_399), .B1(n_512), .B2(n_440), .Y(n_687) );
INVx2_ASAP7_75t_L g688 ( .A(n_609), .Y(n_688) );
BUFx4_ASAP7_75t_L g689 ( .A(n_596), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_617), .A2(n_410), .B1(n_427), .B2(n_425), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_604), .B(n_370), .Y(n_691) );
INVx2_ASAP7_75t_SL g692 ( .A(n_609), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_604), .B(n_371), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_596), .B(n_374), .Y(n_694) );
INVxp67_ASAP7_75t_L g695 ( .A(n_598), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_598), .B(n_386), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_605), .B(n_388), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_605), .B(n_390), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_606), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_606), .B(n_398), .Y(n_700) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_607), .B(n_401), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_607), .A2(n_461), .B1(n_471), .B2(n_458), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_589), .B(n_402), .Y(n_703) );
AND2x4_ASAP7_75t_L g704 ( .A(n_589), .B(n_458), .Y(n_704) );
INVx2_ASAP7_75t_L g705 ( .A(n_595), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_595), .B(n_416), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_597), .B(n_426), .Y(n_707) );
AND2x2_ASAP7_75t_SL g708 ( .A(n_608), .B(n_580), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_615), .B(n_432), .Y(n_709) );
BUFx3_ASAP7_75t_L g710 ( .A(n_590), .Y(n_710) );
BUFx3_ASAP7_75t_L g711 ( .A(n_590), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_635), .B(n_461), .Y(n_712) );
BUFx12f_ASAP7_75t_L g713 ( .A(n_663), .Y(n_713) );
AND2x6_ASAP7_75t_L g714 ( .A(n_651), .B(n_413), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g715 ( .A1(n_677), .A2(n_580), .B(n_351), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_631), .B(n_376), .Y(n_716) );
NAND3xp33_ASAP7_75t_L g717 ( .A(n_639), .B(n_408), .C(n_394), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_629), .Y(n_718) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_632), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_636), .B(n_422), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_678), .B(n_440), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_645), .Y(n_722) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_632), .Y(n_723) );
NOR2xp33_ASAP7_75t_R g724 ( .A(n_683), .B(n_471), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_654), .A2(n_506), .B1(n_485), .B2(n_512), .Y(n_725) );
OAI21xp33_ASAP7_75t_SL g726 ( .A1(n_654), .A2(n_437), .B(n_434), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g727 ( .A1(n_643), .A2(n_535), .B(n_463), .C(n_475), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_636), .B(n_451), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_638), .B(n_628), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_679), .A2(n_580), .B(n_430), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_649), .Y(n_731) );
BUFx6f_ASAP7_75t_L g732 ( .A(n_632), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_702), .B(n_538), .C(n_502), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_643), .B(n_499), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_656), .B(n_485), .Y(n_735) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_708), .A2(n_695), .B(n_667), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_648), .A2(n_506), .B1(n_476), .B2(n_482), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_695), .A2(n_580), .B(n_469), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_650), .B(n_504), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_671), .B(n_516), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_671), .B(n_520), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_640), .B(n_522), .Y(n_742) );
BUFx12f_ASAP7_75t_L g743 ( .A(n_669), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_682), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_704), .A2(n_483), .B1(n_494), .B2(n_459), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_653), .A2(n_523), .B1(n_510), .B2(n_517), .Y(n_746) );
OAI22x1_ASAP7_75t_L g747 ( .A1(n_673), .A2(n_527), .B1(n_531), .B2(n_503), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_634), .B(n_534), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_644), .A2(n_580), .B(n_484), .Y(n_749) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_658), .B(n_435), .Y(n_750) );
INVx2_ASAP7_75t_L g751 ( .A(n_647), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_704), .B(n_347), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g753 ( .A1(n_708), .A2(n_367), .B(n_355), .Y(n_753) );
NOR2xp67_ASAP7_75t_L g754 ( .A(n_681), .B(n_10), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_667), .B(n_444), .Y(n_755) );
AOI21xp5_ASAP7_75t_L g756 ( .A1(n_699), .A2(n_375), .B(n_373), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_658), .B(n_642), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_657), .A2(n_380), .B(n_378), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_675), .Y(n_759) );
OAI22xp5_ASAP7_75t_SL g760 ( .A1(n_633), .A2(n_444), .B1(n_486), .B2(n_447), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_676), .A2(n_385), .B1(n_392), .B2(n_381), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_676), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g763 ( .A1(n_672), .A2(n_486), .B(n_536), .C(n_447), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_637), .B(n_536), .Y(n_764) );
OAI21x1_ASAP7_75t_L g765 ( .A1(n_646), .A2(n_615), .B(n_372), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_666), .B(n_443), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_666), .B(n_450), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_652), .B(n_454), .Y(n_768) );
AND2x6_ASAP7_75t_L g769 ( .A(n_658), .B(n_413), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_659), .A2(n_525), .B1(n_533), .B2(n_464), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g771 ( .A(n_696), .B(n_466), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_693), .A2(n_412), .B(n_411), .Y(n_772) );
A2O1A1Ixp33_ASAP7_75t_L g773 ( .A1(n_664), .A2(n_519), .B(n_477), .C(n_417), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_664), .B(n_479), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_685), .A2(n_421), .B(n_415), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_681), .A2(n_525), .B1(n_533), .B2(n_464), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_659), .B(n_481), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g778 ( .A(n_691), .B(n_490), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_641), .A2(n_428), .B(n_423), .Y(n_779) );
OR2x6_ASAP7_75t_SL g780 ( .A(n_689), .B(n_500), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_670), .B(n_505), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_660), .A2(n_431), .B1(n_436), .B2(n_429), .Y(n_782) );
OAI22xp5_ASAP7_75t_L g783 ( .A1(n_680), .A2(n_525), .B1(n_533), .B2(n_464), .Y(n_783) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_647), .B(n_507), .Y(n_784) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_694), .A2(n_448), .B(n_442), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_686), .B(n_690), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_697), .A2(n_457), .B(n_453), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g788 ( .A1(n_687), .A2(n_464), .B1(n_533), .B2(n_525), .C(n_468), .Y(n_788) );
NAND2xp33_ASAP7_75t_L g789 ( .A(n_647), .B(n_508), .Y(n_789) );
AOI21xp5_ASAP7_75t_L g790 ( .A1(n_698), .A2(n_473), .B(n_472), .Y(n_790) );
OR2x2_ASAP7_75t_L g791 ( .A(n_687), .B(n_11), .Y(n_791) );
OR2x6_ASAP7_75t_L g792 ( .A(n_661), .B(n_439), .Y(n_792) );
NAND2x1_ASAP7_75t_L g793 ( .A(n_647), .B(n_369), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_703), .A2(n_480), .B(n_474), .Y(n_794) );
NAND2x1p5_ASAP7_75t_L g795 ( .A(n_700), .B(n_452), .Y(n_795) );
NOR2xp33_ASAP7_75t_L g796 ( .A(n_701), .B(n_513), .Y(n_796) );
NAND2xp5_ASAP7_75t_SL g797 ( .A(n_706), .B(n_487), .Y(n_797) );
AOI21xp5_ASAP7_75t_L g798 ( .A1(n_707), .A2(n_489), .B(n_488), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_688), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_686), .B(n_491), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_705), .A2(n_496), .B(n_493), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g802 ( .A1(n_655), .A2(n_498), .B(n_497), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_646), .B(n_514), .Y(n_803) );
NOR2xp33_ASAP7_75t_SL g804 ( .A(n_630), .B(n_452), .Y(n_804) );
AO21x1_ASAP7_75t_L g805 ( .A1(n_665), .A2(n_521), .B(n_518), .Y(n_805) );
AOI21xp5_ASAP7_75t_L g806 ( .A1(n_709), .A2(n_526), .B(n_524), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_680), .A2(n_532), .B1(n_537), .B2(n_530), .Y(n_807) );
A2O1A1Ixp33_ASAP7_75t_L g808 ( .A1(n_668), .A2(n_540), .B(n_391), .C(n_395), .Y(n_808) );
INVx8_ASAP7_75t_L g809 ( .A(n_690), .Y(n_809) );
BUFx3_ASAP7_75t_L g810 ( .A(n_662), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g811 ( .A1(n_674), .A2(n_391), .B(n_384), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_684), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_692), .B(n_11), .Y(n_813) );
O2A1O1Ixp33_ASAP7_75t_L g814 ( .A1(n_710), .A2(n_407), .B(n_424), .C(n_403), .Y(n_814) );
OAI22xp5_ASAP7_75t_L g815 ( .A1(n_711), .A2(n_424), .B1(n_465), .B2(n_407), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_636), .B(n_12), .Y(n_816) );
INVx6_ASAP7_75t_L g817 ( .A(n_628), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_678), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_629), .Y(n_819) );
AOI221xp5_ASAP7_75t_L g820 ( .A1(n_639), .A2(n_515), .B1(n_529), .B2(n_467), .C(n_465), .Y(n_820) );
OAI21x1_ASAP7_75t_L g821 ( .A1(n_657), .A2(n_615), .B(n_515), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_677), .A2(n_529), .B(n_467), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g823 ( .A(n_636), .B(n_13), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_629), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_631), .B(n_13), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_648), .A2(n_557), .B1(n_561), .B2(n_558), .Y(n_826) );
BUFx6f_ASAP7_75t_L g827 ( .A(n_632), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_648), .A2(n_558), .B1(n_562), .B2(n_561), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_635), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_631), .B(n_14), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_635), .B(n_14), .Y(n_831) );
OAI21xp5_ASAP7_75t_L g832 ( .A1(n_708), .A2(n_563), .B(n_562), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_648), .A2(n_565), .B1(n_573), .B2(n_563), .Y(n_833) );
INVx2_ASAP7_75t_L g834 ( .A(n_632), .Y(n_834) );
BUFx3_ASAP7_75t_L g835 ( .A(n_635), .Y(n_835) );
A2O1A1Ixp33_ASAP7_75t_L g836 ( .A1(n_631), .A2(n_565), .B(n_573), .C(n_563), .Y(n_836) );
NOR2xp67_ASAP7_75t_SL g837 ( .A(n_658), .B(n_553), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_631), .B(n_16), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_631), .B(n_16), .Y(n_839) );
BUFx2_ASAP7_75t_SL g840 ( .A(n_635), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_629), .Y(n_841) );
AO32x2_ASAP7_75t_L g842 ( .A1(n_638), .A2(n_572), .A3(n_570), .B1(n_560), .B2(n_565), .Y(n_842) );
OAI22xp5_ASAP7_75t_L g843 ( .A1(n_809), .A2(n_573), .B1(n_577), .B2(n_553), .Y(n_843) );
AO31x2_ASAP7_75t_L g844 ( .A1(n_805), .A2(n_577), .A3(n_560), .B(n_572), .Y(n_844) );
INVx2_ASAP7_75t_SL g845 ( .A(n_835), .Y(n_845) );
OAI21x1_ASAP7_75t_L g846 ( .A1(n_821), .A2(n_577), .B(n_570), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_729), .B(n_17), .Y(n_847) );
OAI21x1_ASAP7_75t_L g848 ( .A1(n_765), .A2(n_570), .B(n_560), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_762), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_786), .B(n_742), .Y(n_850) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_780), .Y(n_851) );
O2A1O1Ixp33_ASAP7_75t_L g852 ( .A1(n_727), .A2(n_19), .B(n_17), .C(n_18), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_715), .A2(n_590), .B(n_553), .Y(n_853) );
NAND3xp33_ASAP7_75t_L g854 ( .A(n_776), .B(n_553), .C(n_560), .Y(n_854) );
OA21x2_ASAP7_75t_L g855 ( .A1(n_738), .A2(n_572), .B(n_570), .Y(n_855) );
AO32x2_ASAP7_75t_L g856 ( .A1(n_783), .A2(n_570), .A3(n_572), .B1(n_20), .B2(n_21), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_726), .B(n_18), .Y(n_857) );
INVx2_ASAP7_75t_SL g858 ( .A(n_817), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_809), .B(n_19), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_829), .B(n_20), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_744), .Y(n_861) );
OAI21xp5_ASAP7_75t_L g862 ( .A1(n_749), .A2(n_572), .B(n_570), .Y(n_862) );
BUFx4_ASAP7_75t_SL g863 ( .A(n_791), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_809), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_730), .A2(n_590), .B(n_149), .Y(n_865) );
OAI21x1_ASAP7_75t_L g866 ( .A1(n_832), .A2(n_151), .B(n_147), .Y(n_866) );
INVx3_ASAP7_75t_R g867 ( .A(n_743), .Y(n_867) );
INVxp67_ASAP7_75t_SL g868 ( .A(n_725), .Y(n_868) );
BUFx3_ASAP7_75t_L g869 ( .A(n_817), .Y(n_869) );
OR2x2_ASAP7_75t_L g870 ( .A(n_721), .B(n_23), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_799), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_840), .B(n_25), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_736), .A2(n_28), .B1(n_26), .B2(n_27), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_753), .A2(n_154), .B(n_152), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g875 ( .A1(n_818), .A2(n_30), .B1(n_28), .B2(n_29), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g876 ( .A1(n_772), .A2(n_159), .B(n_155), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_825), .A2(n_32), .B1(n_30), .B2(n_31), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_752), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_758), .A2(n_164), .B(n_163), .Y(n_879) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_830), .A2(n_33), .B1(n_31), .B2(n_32), .Y(n_880) );
AND2x6_ASAP7_75t_L g881 ( .A(n_718), .B(n_33), .Y(n_881) );
NAND2x1p5_ASAP7_75t_L g882 ( .A(n_712), .B(n_34), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_816), .B(n_34), .Y(n_883) );
INVx2_ASAP7_75t_L g884 ( .A(n_722), .Y(n_884) );
BUFx6f_ASAP7_75t_L g885 ( .A(n_719), .Y(n_885) );
AOI21xp5_ASAP7_75t_L g886 ( .A1(n_774), .A2(n_173), .B(n_172), .Y(n_886) );
AND2x4_ASAP7_75t_L g887 ( .A(n_831), .B(n_35), .Y(n_887) );
INVx2_ASAP7_75t_SL g888 ( .A(n_724), .Y(n_888) );
AOI211x1_ASAP7_75t_L g889 ( .A1(n_717), .A2(n_40), .B(n_35), .C(n_37), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g890 ( .A1(n_737), .A2(n_43), .B1(n_41), .B2(n_42), .Y(n_890) );
OAI21x1_ASAP7_75t_L g891 ( .A1(n_793), .A2(n_176), .B(n_175), .Y(n_891) );
AND2x4_ASAP7_75t_L g892 ( .A(n_731), .B(n_42), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g893 ( .A(n_823), .B(n_43), .Y(n_893) );
BUFx2_ASAP7_75t_L g894 ( .A(n_769), .Y(n_894) );
INVx3_ASAP7_75t_L g895 ( .A(n_713), .Y(n_895) );
BUFx3_ASAP7_75t_L g896 ( .A(n_812), .Y(n_896) );
INVxp67_ASAP7_75t_L g897 ( .A(n_740), .Y(n_897) );
AO32x2_ASAP7_75t_L g898 ( .A1(n_770), .A2(n_44), .A3(n_45), .B1(n_46), .B2(n_47), .Y(n_898) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_797), .A2(n_180), .B(n_179), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g900 ( .A1(n_806), .A2(n_186), .B(n_181), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_755), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_733), .B(n_45), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_739), .B(n_47), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_741), .Y(n_904) );
INVx2_ASAP7_75t_SL g905 ( .A(n_795), .Y(n_905) );
AOI21xp5_ASAP7_75t_L g906 ( .A1(n_779), .A2(n_195), .B(n_191), .Y(n_906) );
NAND2xp5_ASAP7_75t_SL g907 ( .A(n_720), .B(n_48), .Y(n_907) );
INVx1_ASAP7_75t_SL g908 ( .A(n_728), .Y(n_908) );
AOI21xp33_ASAP7_75t_L g909 ( .A1(n_768), .A2(n_48), .B(n_49), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_745), .B(n_49), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_819), .Y(n_911) );
AND2x4_ASAP7_75t_L g912 ( .A(n_824), .B(n_50), .Y(n_912) );
AND2x4_ASAP7_75t_L g913 ( .A(n_841), .B(n_50), .Y(n_913) );
AOI21xp5_ASAP7_75t_L g914 ( .A1(n_778), .A2(n_199), .B(n_198), .Y(n_914) );
AO31x2_ASAP7_75t_L g915 ( .A1(n_773), .A2(n_51), .A3(n_52), .B(n_53), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_761), .B(n_51), .Y(n_916) );
OAI21xp33_ASAP7_75t_L g917 ( .A1(n_716), .A2(n_52), .B(n_53), .Y(n_917) );
OAI21xp5_ASAP7_75t_L g918 ( .A1(n_775), .A2(n_202), .B(n_200), .Y(n_918) );
AO21x2_ASAP7_75t_L g919 ( .A1(n_836), .A2(n_206), .B(n_205), .Y(n_919) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_735), .B(n_54), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g921 ( .A1(n_838), .A2(n_210), .B(n_208), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_760), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_922) );
NAND3xp33_ASAP7_75t_SL g923 ( .A(n_788), .B(n_56), .C(n_57), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_822), .A2(n_212), .B(n_211), .Y(n_924) );
BUFx6f_ASAP7_75t_L g925 ( .A(n_719), .Y(n_925) );
OAI21xp5_ASAP7_75t_L g926 ( .A1(n_756), .A2(n_215), .B(n_214), .Y(n_926) );
AOI21xp5_ASAP7_75t_L g927 ( .A1(n_839), .A2(n_217), .B(n_216), .Y(n_927) );
AOI21xp5_ASAP7_75t_L g928 ( .A1(n_785), .A2(n_219), .B(n_218), .Y(n_928) );
BUFx4f_ASAP7_75t_L g929 ( .A(n_792), .Y(n_929) );
AOI21xp5_ASAP7_75t_L g930 ( .A1(n_787), .A2(n_223), .B(n_220), .Y(n_930) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_792), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_746), .B(n_58), .Y(n_932) );
AO221x2_ASAP7_75t_L g933 ( .A1(n_747), .A2(n_58), .B1(n_59), .B2(n_60), .C(n_62), .Y(n_933) );
INVx5_ASAP7_75t_L g934 ( .A(n_769), .Y(n_934) );
OAI21xp33_ASAP7_75t_L g935 ( .A1(n_734), .A2(n_60), .B(n_63), .Y(n_935) );
NAND3xp33_ASAP7_75t_L g936 ( .A(n_820), .B(n_63), .C(n_64), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_808), .A2(n_64), .A3(n_65), .B(n_66), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_800), .Y(n_938) );
AOI21xp5_ASAP7_75t_L g939 ( .A1(n_790), .A2(n_227), .B(n_225), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_748), .B(n_66), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_813), .Y(n_941) );
A2O1A1Ixp33_ASAP7_75t_L g942 ( .A1(n_763), .A2(n_67), .B(n_68), .C(n_69), .Y(n_942) );
BUFx10_ASAP7_75t_L g943 ( .A(n_764), .Y(n_943) );
INVxp67_ASAP7_75t_L g944 ( .A(n_803), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_782), .B(n_67), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_766), .A2(n_68), .B1(n_69), .B2(n_70), .Y(n_946) );
AOI21xp5_ASAP7_75t_L g947 ( .A1(n_794), .A2(n_229), .B(n_228), .Y(n_947) );
O2A1O1Ixp33_ASAP7_75t_SL g948 ( .A1(n_757), .A2(n_257), .B(n_341), .C(n_340), .Y(n_948) );
OAI21x1_ASAP7_75t_SL g949 ( .A1(n_802), .A2(n_71), .B(n_72), .Y(n_949) );
OAI21xp5_ASAP7_75t_L g950 ( .A1(n_798), .A2(n_233), .B(n_230), .Y(n_950) );
BUFx8_ASAP7_75t_L g951 ( .A(n_759), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_751), .Y(n_952) );
INVx2_ASAP7_75t_SL g953 ( .A(n_784), .Y(n_953) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_807), .B(n_73), .Y(n_954) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_777), .A2(n_237), .B(n_236), .Y(n_955) );
OAI22x1_ASAP7_75t_L g956 ( .A1(n_754), .A2(n_74), .B1(n_76), .B2(n_78), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_811), .Y(n_957) );
OAI21xp5_ASAP7_75t_L g958 ( .A1(n_801), .A2(n_242), .B(n_240), .Y(n_958) );
OAI22xp5_ASAP7_75t_L g959 ( .A1(n_767), .A2(n_74), .B1(n_76), .B2(n_79), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_815), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_781), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_961) );
BUFx2_ASAP7_75t_L g962 ( .A(n_769), .Y(n_962) );
AOI21xp5_ASAP7_75t_L g963 ( .A1(n_834), .A2(n_272), .B(n_338), .Y(n_963) );
INVx5_ASAP7_75t_L g964 ( .A(n_769), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_771), .B(n_80), .Y(n_965) );
OAI21x1_ASAP7_75t_L g966 ( .A1(n_826), .A2(n_268), .B(n_337), .Y(n_966) );
BUFx2_ASAP7_75t_L g967 ( .A(n_810), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_828), .A2(n_266), .B(n_333), .Y(n_968) );
NAND2xp5_ASAP7_75t_SL g969 ( .A(n_804), .B(n_83), .Y(n_969) );
BUFx10_ASAP7_75t_L g970 ( .A(n_796), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g971 ( .A1(n_833), .A2(n_85), .B1(n_86), .B2(n_87), .Y(n_971) );
OAI21xp5_ASAP7_75t_L g972 ( .A1(n_814), .A2(n_274), .B(n_332), .Y(n_972) );
OAI21xp5_ASAP7_75t_L g973 ( .A1(n_750), .A2(n_273), .B(n_330), .Y(n_973) );
OAI22x1_ASAP7_75t_L g974 ( .A1(n_842), .A2(n_85), .B1(n_86), .B2(n_88), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_842), .Y(n_975) );
AOI21xp33_ASAP7_75t_L g976 ( .A1(n_789), .A2(n_89), .B(n_91), .Y(n_976) );
AO31x2_ASAP7_75t_L g977 ( .A1(n_842), .A2(n_89), .A3(n_91), .B(n_92), .Y(n_977) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_723), .A2(n_280), .B(n_328), .Y(n_978) );
AND2x6_ASAP7_75t_L g979 ( .A(n_723), .B(n_93), .Y(n_979) );
INVx2_ASAP7_75t_L g980 ( .A(n_732), .Y(n_980) );
INVx1_ASAP7_75t_L g981 ( .A(n_732), .Y(n_981) );
AO32x2_ASAP7_75t_L g982 ( .A1(n_714), .A2(n_94), .A3(n_95), .B1(n_96), .B2(n_97), .Y(n_982) );
OA21x2_ASAP7_75t_L g983 ( .A1(n_714), .A2(n_827), .B(n_837), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_714), .A2(n_95), .B1(n_97), .B2(n_98), .Y(n_984) );
BUFx12f_ASAP7_75t_L g985 ( .A(n_827), .Y(n_985) );
OAI21x1_ASAP7_75t_L g986 ( .A1(n_714), .A2(n_282), .B(n_324), .Y(n_986) );
AND2x2_ASAP7_75t_L g987 ( .A(n_729), .B(n_98), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_762), .Y(n_988) );
INVx1_ASAP7_75t_L g989 ( .A(n_762), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_817), .B(n_99), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_729), .B(n_99), .Y(n_991) );
BUFx6f_ASAP7_75t_L g992 ( .A(n_719), .Y(n_992) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_809), .A2(n_100), .B1(n_101), .B2(n_102), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_762), .B(n_102), .Y(n_994) );
INVx1_ASAP7_75t_L g995 ( .A(n_762), .Y(n_995) );
BUFx6f_ASAP7_75t_L g996 ( .A(n_719), .Y(n_996) );
AND2x4_ASAP7_75t_L g997 ( .A(n_762), .B(n_103), .Y(n_997) );
AOI21xp33_ASAP7_75t_L g998 ( .A1(n_729), .A2(n_103), .B(n_104), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_809), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_999) );
A2O1A1Ixp33_ASAP7_75t_L g1000 ( .A1(n_753), .A2(n_105), .B(n_107), .C(n_108), .Y(n_1000) );
A2O1A1Ixp33_ASAP7_75t_L g1001 ( .A1(n_753), .A2(n_107), .B(n_108), .C(n_109), .Y(n_1001) );
INVxp67_ASAP7_75t_SL g1002 ( .A(n_725), .Y(n_1002) );
AO31x2_ASAP7_75t_L g1003 ( .A1(n_805), .A2(n_110), .A3(n_111), .B(n_112), .Y(n_1003) );
BUFx2_ASAP7_75t_L g1004 ( .A(n_724), .Y(n_1004) );
AOI221xp5_ASAP7_75t_SL g1005 ( .A1(n_788), .A2(n_112), .B1(n_113), .B2(n_114), .C(n_115), .Y(n_1005) );
AOI21xp33_ASAP7_75t_L g1006 ( .A1(n_850), .A2(n_115), .B(n_116), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_868), .B(n_116), .Y(n_1007) );
NAND2x1p5_ASAP7_75t_L g1008 ( .A(n_869), .B(n_117), .Y(n_1008) );
OAI21x1_ASAP7_75t_SL g1009 ( .A1(n_949), .A2(n_117), .B(n_118), .Y(n_1009) );
INVx2_ASAP7_75t_L g1010 ( .A(n_884), .Y(n_1010) );
INVx5_ASAP7_75t_L g1011 ( .A(n_979), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1002), .B(n_901), .Y(n_1012) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_944), .B(n_908), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_867), .Y(n_1014) );
BUFx10_ASAP7_75t_L g1015 ( .A(n_994), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_878), .B(n_120), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_897), .B(n_122), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_861), .B(n_122), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1019 ( .A(n_888), .B(n_123), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_911), .Y(n_1020) );
AO21x2_ASAP7_75t_L g1021 ( .A1(n_975), .A2(n_846), .B(n_972), .Y(n_1021) );
OR2x2_ASAP7_75t_L g1022 ( .A(n_870), .B(n_124), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_957), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_892), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_851), .Y(n_1025) );
INVx2_ASAP7_75t_L g1026 ( .A(n_871), .Y(n_1026) );
NAND2x1p5_ASAP7_75t_L g1027 ( .A(n_845), .B(n_124), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_849), .Y(n_1028) );
INVx2_ASAP7_75t_L g1029 ( .A(n_988), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_938), .Y(n_1030) );
AO31x2_ASAP7_75t_L g1031 ( .A1(n_974), .A2(n_127), .A3(n_129), .B(n_132), .Y(n_1031) );
BUFx6f_ASAP7_75t_L g1032 ( .A(n_985), .Y(n_1032) );
INVxp67_ASAP7_75t_SL g1033 ( .A(n_892), .Y(n_1033) );
AOI21xp33_ASAP7_75t_SL g1034 ( .A1(n_895), .A2(n_127), .B(n_129), .Y(n_1034) );
OA21x2_ASAP7_75t_L g1035 ( .A1(n_866), .A2(n_291), .B(n_308), .Y(n_1035) );
INVx2_ASAP7_75t_L g1036 ( .A(n_989), .Y(n_1036) );
AO31x2_ASAP7_75t_L g1037 ( .A1(n_873), .A2(n_132), .A3(n_133), .B(n_134), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_1004), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_904), .A2(n_133), .B1(n_135), .B2(n_243), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_987), .B(n_135), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_912), .Y(n_1041) );
INVx2_ASAP7_75t_L g1042 ( .A(n_995), .Y(n_1042) );
AO31x2_ASAP7_75t_L g1043 ( .A1(n_843), .A2(n_247), .A3(n_248), .B(n_250), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_860), .B(n_251), .Y(n_1044) );
NAND2x1p5_ASAP7_75t_L g1045 ( .A(n_934), .B(n_964), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_856), .Y(n_1046) );
OA21x2_ASAP7_75t_L g1047 ( .A1(n_966), .A2(n_255), .B(n_264), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_912), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_858), .B(n_292), .Y(n_1049) );
NOR2xp33_ASAP7_75t_L g1050 ( .A(n_943), .B(n_295), .Y(n_1050) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_863), .Y(n_1051) );
OA21x2_ASAP7_75t_L g1052 ( .A1(n_968), .A2(n_296), .B(n_298), .Y(n_1052) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_979), .Y(n_1053) );
NAND2x1p5_ASAP7_75t_L g1054 ( .A(n_934), .B(n_302), .Y(n_1054) );
NAND2x1p5_ASAP7_75t_L g1055 ( .A(n_934), .B(n_964), .Y(n_1055) );
OR2x2_ASAP7_75t_L g1056 ( .A(n_967), .B(n_303), .Y(n_1056) );
INVx2_ASAP7_75t_L g1057 ( .A(n_856), .Y(n_1057) );
NOR2xp67_ASAP7_75t_SL g1058 ( .A(n_964), .B(n_305), .Y(n_1058) );
OAI21x1_ASAP7_75t_L g1059 ( .A1(n_986), .A2(n_891), .B(n_924), .Y(n_1059) );
AOI21xp5_ASAP7_75t_L g1060 ( .A1(n_941), .A2(n_874), .B(n_883), .Y(n_1060) );
AOI21xp5_ASAP7_75t_L g1061 ( .A1(n_893), .A2(n_955), .B(n_886), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_903), .B(n_945), .Y(n_1062) );
AND2x2_ASAP7_75t_L g1063 ( .A(n_860), .B(n_994), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_856), .Y(n_1064) );
AO31x2_ASAP7_75t_L g1065 ( .A1(n_1000), .A2(n_1001), .A3(n_942), .B(n_960), .Y(n_1065) );
INVx2_ASAP7_75t_L g1066 ( .A(n_952), .Y(n_1066) );
OAI21xp5_ASAP7_75t_L g1067 ( .A1(n_936), .A2(n_847), .B(n_991), .Y(n_1067) );
AO31x2_ASAP7_75t_L g1068 ( .A1(n_864), .A2(n_993), .A3(n_959), .B(n_946), .Y(n_1068) );
INVx1_ASAP7_75t_L g1069 ( .A(n_913), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_910), .B(n_887), .Y(n_1070) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_887), .B(n_940), .Y(n_1071) );
AND2x4_ASAP7_75t_L g1072 ( .A(n_872), .B(n_953), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_913), .Y(n_1073) );
AND2x4_ASAP7_75t_L g1074 ( .A(n_896), .B(n_997), .Y(n_1074) );
INVx1_ASAP7_75t_L g1075 ( .A(n_881), .Y(n_1075) );
OAI21xp5_ASAP7_75t_L g1076 ( .A1(n_923), .A2(n_916), .B(n_965), .Y(n_1076) );
AOI22xp5_ASAP7_75t_L g1077 ( .A1(n_920), .A2(n_990), .B1(n_902), .B2(n_859), .Y(n_1077) );
NAND2xp5_ASAP7_75t_SL g1078 ( .A(n_882), .B(n_885), .Y(n_1078) );
AO31x2_ASAP7_75t_L g1079 ( .A1(n_921), .A2(n_927), .A3(n_956), .B(n_877), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_881), .Y(n_1080) );
OA21x2_ASAP7_75t_L g1081 ( .A1(n_1005), .A2(n_918), .B(n_950), .Y(n_1081) );
INVxp33_ASAP7_75t_L g1082 ( .A(n_929), .Y(n_1082) );
OA21x2_ASAP7_75t_L g1083 ( .A1(n_958), .A2(n_926), .B(n_935), .Y(n_1083) );
INVx3_ASAP7_75t_L g1084 ( .A(n_885), .Y(n_1084) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_933), .B(n_922), .Y(n_1085) );
NOR2xp33_ASAP7_75t_L g1086 ( .A(n_970), .B(n_931), .Y(n_1086) );
OA21x2_ASAP7_75t_L g1087 ( .A1(n_917), .A2(n_879), .B(n_973), .Y(n_1087) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_979), .Y(n_1088) );
OA21x2_ASAP7_75t_L g1089 ( .A1(n_906), .A2(n_876), .B(n_900), .Y(n_1089) );
INVx1_ASAP7_75t_L g1090 ( .A(n_857), .Y(n_1090) );
INVx3_ASAP7_75t_L g1091 ( .A(n_925), .Y(n_1091) );
OAI21x1_ASAP7_75t_SL g1092 ( .A1(n_983), .A2(n_890), .B(n_905), .Y(n_1092) );
OAI21x1_ASAP7_75t_L g1093 ( .A1(n_980), .A2(n_981), .B(n_978), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_954), .B(n_907), .Y(n_1094) );
AO31x2_ASAP7_75t_L g1095 ( .A1(n_880), .A2(n_971), .A3(n_963), .B(n_930), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1096 ( .A(n_875), .B(n_932), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_951), .B(n_909), .Y(n_1097) );
A2O1A1Ixp33_ASAP7_75t_L g1098 ( .A1(n_852), .A2(n_961), .B(n_998), .C(n_939), .Y(n_1098) );
OR2x2_ASAP7_75t_L g1099 ( .A(n_933), .B(n_915), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1100 ( .A(n_951), .B(n_999), .Y(n_1100) );
A2O1A1Ixp33_ASAP7_75t_L g1101 ( .A1(n_928), .A2(n_976), .B(n_947), .C(n_914), .Y(n_1101) );
OA21x2_ASAP7_75t_L g1102 ( .A1(n_854), .A2(n_899), .B(n_984), .Y(n_1102) );
OR2x2_ASAP7_75t_L g1103 ( .A(n_915), .B(n_1003), .Y(n_1103) );
AND2x4_ASAP7_75t_L g1104 ( .A(n_894), .B(n_962), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1003), .Y(n_1105) );
OR2x2_ASAP7_75t_L g1106 ( .A(n_915), .B(n_1003), .Y(n_1106) );
AO31x2_ASAP7_75t_L g1107 ( .A1(n_844), .A2(n_977), .A3(n_889), .B(n_937), .Y(n_1107) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_969), .A2(n_919), .B1(n_996), .B2(n_992), .Y(n_1108) );
NOR2x1_ASAP7_75t_SL g1109 ( .A(n_996), .B(n_982), .Y(n_1109) );
OA21x2_ASAP7_75t_L g1110 ( .A1(n_844), .A2(n_977), .B(n_982), .Y(n_1110) );
AO31x2_ASAP7_75t_L g1111 ( .A1(n_977), .A2(n_937), .A3(n_982), .B(n_898), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_898), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_898), .Y(n_1113) );
OA21x2_ASAP7_75t_L g1114 ( .A1(n_948), .A2(n_862), .B(n_975), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_870), .B(n_725), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_861), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_868), .A2(n_809), .B1(n_633), .B2(n_818), .Y(n_1117) );
AOI21xp5_ASAP7_75t_L g1118 ( .A1(n_862), .A2(n_738), .B(n_853), .Y(n_1118) );
BUFx6f_ASAP7_75t_L g1119 ( .A(n_985), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_861), .Y(n_1120) );
INVx1_ASAP7_75t_L g1121 ( .A(n_861), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_849), .B(n_762), .Y(n_1122) );
OA21x2_ASAP7_75t_L g1123 ( .A1(n_862), .A2(n_975), .B(n_846), .Y(n_1123) );
OAI21x1_ASAP7_75t_L g1124 ( .A1(n_848), .A2(n_846), .B(n_862), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_868), .B(n_627), .Y(n_1125) );
NAND2x1p5_ASAP7_75t_L g1126 ( .A(n_869), .B(n_845), .Y(n_1126) );
OAI21x1_ASAP7_75t_SL g1127 ( .A1(n_949), .A2(n_972), .B(n_736), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_851), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_861), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_870), .B(n_725), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_861), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_869), .Y(n_1132) );
NOR2x1_ASAP7_75t_R g1133 ( .A(n_851), .B(n_545), .Y(n_1133) );
CKINVDCx5p33_ASAP7_75t_R g1134 ( .A(n_851), .Y(n_1134) );
A2O1A1Ixp33_ASAP7_75t_L g1135 ( .A1(n_850), .A2(n_903), .B(n_965), .C(n_852), .Y(n_1135) );
INVx3_ASAP7_75t_L g1136 ( .A(n_985), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_861), .Y(n_1137) );
INVx4_ASAP7_75t_SL g1138 ( .A(n_979), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_861), .Y(n_1139) );
INVx2_ASAP7_75t_L g1140 ( .A(n_884), .Y(n_1140) );
AOI21x1_ASAP7_75t_L g1141 ( .A1(n_975), .A2(n_855), .B(n_862), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1142 ( .A(n_868), .B(n_631), .Y(n_1142) );
AOI21xp33_ASAP7_75t_SL g1143 ( .A1(n_851), .A2(n_725), .B(n_678), .Y(n_1143) );
AOI21xp5_ASAP7_75t_L g1144 ( .A1(n_862), .A2(n_738), .B(n_853), .Y(n_1144) );
AOI21xp5_ASAP7_75t_L g1145 ( .A1(n_862), .A2(n_738), .B(n_853), .Y(n_1145) );
OAI21x1_ASAP7_75t_L g1146 ( .A1(n_848), .A2(n_846), .B(n_862), .Y(n_1146) );
AO21x2_ASAP7_75t_L g1147 ( .A1(n_862), .A2(n_975), .B(n_865), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_861), .Y(n_1148) );
AO31x2_ASAP7_75t_L g1149 ( .A1(n_975), .A2(n_974), .A3(n_805), .B(n_865), .Y(n_1149) );
AOI21xp5_ASAP7_75t_L g1150 ( .A1(n_862), .A2(n_738), .B(n_853), .Y(n_1150) );
OA21x2_ASAP7_75t_L g1151 ( .A1(n_862), .A2(n_975), .B(n_846), .Y(n_1151) );
NAND2xp5_ASAP7_75t_SL g1152 ( .A(n_1004), .B(n_724), .Y(n_1152) );
OAI21x1_ASAP7_75t_L g1153 ( .A1(n_848), .A2(n_846), .B(n_862), .Y(n_1153) );
BUFx2_ASAP7_75t_L g1154 ( .A(n_869), .Y(n_1154) );
OA21x2_ASAP7_75t_L g1155 ( .A1(n_862), .A2(n_975), .B(n_846), .Y(n_1155) );
OAI22xp5_ASAP7_75t_L g1156 ( .A1(n_868), .A2(n_809), .B1(n_704), .B2(n_737), .Y(n_1156) );
INVx1_ASAP7_75t_SL g1157 ( .A(n_1032), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1023), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1125), .B(n_1142), .Y(n_1159) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1116), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1116), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1120), .Y(n_1162) );
AO21x2_ASAP7_75t_L g1163 ( .A1(n_1127), .A2(n_1144), .B(n_1118), .Y(n_1163) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1141), .Y(n_1164) );
AO21x2_ASAP7_75t_L g1165 ( .A1(n_1145), .A2(n_1150), .B(n_1105), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1120), .Y(n_1166) );
OR2x6_ASAP7_75t_L g1167 ( .A(n_1053), .B(n_1088), .Y(n_1167) );
INVx2_ASAP7_75t_L g1168 ( .A(n_1123), .Y(n_1168) );
INVx2_ASAP7_75t_L g1169 ( .A(n_1151), .Y(n_1169) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1121), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1022), .B(n_1115), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1121), .Y(n_1172) );
OAI21xp5_ASAP7_75t_L g1173 ( .A1(n_1135), .A2(n_1098), .B(n_1076), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1151), .Y(n_1174) );
HB1xp67_ASAP7_75t_L g1175 ( .A(n_1011), .Y(n_1175) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1155), .Y(n_1176) );
INVx4_ASAP7_75t_L g1177 ( .A(n_1138), .Y(n_1177) );
INVx1_ASAP7_75t_L g1178 ( .A(n_1129), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1129), .Y(n_1179) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_1032), .Y(n_1180) );
OA21x2_ASAP7_75t_L g1181 ( .A1(n_1124), .A2(n_1153), .B(n_1146), .Y(n_1181) );
OR2x6_ASAP7_75t_L g1182 ( .A(n_1075), .B(n_1080), .Y(n_1182) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1010), .B(n_1140), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1131), .Y(n_1184) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_1011), .Y(n_1185) );
INVx3_ASAP7_75t_L g1186 ( .A(n_1011), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1130), .B(n_1013), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_1032), .Y(n_1188) );
HB1xp67_ASAP7_75t_L g1189 ( .A(n_1033), .Y(n_1189) );
INVx2_ASAP7_75t_SL g1190 ( .A(n_1119), .Y(n_1190) );
INVx3_ASAP7_75t_L g1191 ( .A(n_1045), .Y(n_1191) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1070), .B(n_1063), .Y(n_1192) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1055), .Y(n_1193) );
AND2x4_ASAP7_75t_L g1194 ( .A(n_1030), .B(n_1104), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1195 ( .A(n_1028), .B(n_1029), .Y(n_1195) );
BUFx2_ASAP7_75t_L g1196 ( .A(n_1119), .Y(n_1196) );
INVx3_ASAP7_75t_L g1197 ( .A(n_1084), .Y(n_1197) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1137), .Y(n_1198) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1137), .Y(n_1199) );
INVx1_ASAP7_75t_L g1200 ( .A(n_1139), .Y(n_1200) );
BUFx6f_ASAP7_75t_L g1201 ( .A(n_1084), .Y(n_1201) );
INVx1_ASAP7_75t_SL g1202 ( .A(n_1119), .Y(n_1202) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1030), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1204 ( .A(n_1136), .Y(n_1204) );
AO21x2_ASAP7_75t_L g1205 ( .A1(n_1092), .A2(n_1021), .B(n_1147), .Y(n_1205) );
AND2x4_ASAP7_75t_L g1206 ( .A(n_1104), .B(n_1139), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1148), .Y(n_1207) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1148), .Y(n_1208) );
AO31x2_ASAP7_75t_L g1209 ( .A1(n_1109), .A2(n_1046), .A3(n_1057), .B(n_1064), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1020), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1211 ( .A(n_1117), .B(n_1012), .Y(n_1211) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1036), .Y(n_1212) );
INVx1_ASAP7_75t_SL g1213 ( .A(n_1136), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1042), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1215 ( .A(n_1071), .B(n_1074), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1026), .Y(n_1216) );
OA21x2_ASAP7_75t_L g1217 ( .A1(n_1103), .A2(n_1106), .B(n_1112), .Y(n_1217) );
BUFx2_ASAP7_75t_L g1218 ( .A(n_1074), .Y(n_1218) );
OAI211xp5_ASAP7_75t_L g1219 ( .A1(n_1143), .A2(n_1077), .B(n_1034), .C(n_1100), .Y(n_1219) );
NOR2xp33_ASAP7_75t_R g1220 ( .A(n_1014), .B(n_1051), .Y(n_1220) );
OAI22xp5_ASAP7_75t_L g1221 ( .A1(n_1156), .A2(n_1096), .B1(n_1062), .B2(n_1099), .Y(n_1221) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1018), .Y(n_1222) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1016), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1066), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1122), .B(n_1056), .Y(n_1225) );
AO21x1_ASAP7_75t_SL g1226 ( .A1(n_1024), .A2(n_1069), .B(n_1048), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1122), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1090), .B(n_1085), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1113), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1027), .Y(n_1230) );
INVx3_ASAP7_75t_L g1231 ( .A(n_1091), .Y(n_1231) );
OAI211xp5_ASAP7_75t_L g1232 ( .A1(n_1097), .A2(n_1019), .B(n_1152), .C(n_1006), .Y(n_1232) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1017), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1041), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1007), .B(n_1072), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1073), .Y(n_1236) );
OA21x2_ASAP7_75t_L g1237 ( .A1(n_1059), .A2(n_1060), .B(n_1061), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1049), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1008), .Y(n_1239) );
INVx3_ASAP7_75t_L g1240 ( .A(n_1091), .Y(n_1240) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1107), .B(n_1065), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1107), .B(n_1065), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1037), .Y(n_1243) );
INVx5_ASAP7_75t_L g1244 ( .A(n_1015), .Y(n_1244) );
INVx1_ASAP7_75t_L g1245 ( .A(n_1037), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1037), .Y(n_1246) );
AOI21x1_ASAP7_75t_L g1247 ( .A1(n_1083), .A2(n_1114), .B(n_1110), .Y(n_1247) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1040), .B(n_1154), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1107), .B(n_1065), .Y(n_1249) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1031), .Y(n_1250) );
INVx2_ASAP7_75t_SL g1251 ( .A(n_1015), .Y(n_1251) );
INVx1_ASAP7_75t_L g1252 ( .A(n_1031), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1044), .Y(n_1253) );
AO21x2_ASAP7_75t_L g1254 ( .A1(n_1109), .A2(n_1009), .B(n_1108), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1132), .B(n_1126), .Y(n_1255) );
OAI21xp5_ASAP7_75t_L g1256 ( .A1(n_1067), .A2(n_1094), .B(n_1101), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1039), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1111), .B(n_1110), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1111), .B(n_1068), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1111), .B(n_1068), .Y(n_1260) );
OR2x6_ASAP7_75t_L g1261 ( .A(n_1054), .B(n_1078), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1068), .B(n_1149), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1149), .B(n_1079), .Y(n_1263) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1050), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1149), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1086), .B(n_1082), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1079), .B(n_1081), .Y(n_1267) );
INVx2_ASAP7_75t_L g1268 ( .A(n_1093), .Y(n_1268) );
INVx3_ASAP7_75t_L g1269 ( .A(n_1079), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1270 ( .A(n_1043), .B(n_1095), .Y(n_1270) );
OR2x2_ASAP7_75t_L g1271 ( .A(n_1128), .B(n_1134), .Y(n_1271) );
INVx3_ASAP7_75t_L g1272 ( .A(n_1095), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1043), .B(n_1095), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1038), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1275 ( .A(n_1083), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1087), .B(n_1089), .Y(n_1276) );
AOI21x1_ASAP7_75t_L g1277 ( .A1(n_1047), .A2(n_1052), .B(n_1087), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1058), .Y(n_1278) );
BUFx3_ASAP7_75t_L g1279 ( .A(n_1025), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1280 ( .A(n_1089), .B(n_1102), .Y(n_1280) );
OR2x2_ASAP7_75t_SL g1281 ( .A(n_1189), .B(n_1035), .Y(n_1281) );
BUFx12f_ASAP7_75t_L g1282 ( .A(n_1196), .Y(n_1282) );
INVx2_ASAP7_75t_SL g1283 ( .A(n_1244), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1158), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1159), .B(n_1133), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1187), .B(n_1102), .Y(n_1286) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1195), .Y(n_1287) );
INVx3_ASAP7_75t_L g1288 ( .A(n_1186), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1259), .B(n_1035), .Y(n_1289) );
INVx2_ASAP7_75t_SL g1290 ( .A(n_1244), .Y(n_1290) );
INVxp67_ASAP7_75t_L g1291 ( .A(n_1188), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1183), .B(n_1228), .Y(n_1292) );
BUFx2_ASAP7_75t_L g1293 ( .A(n_1189), .Y(n_1293) );
INVx3_ASAP7_75t_L g1294 ( .A(n_1186), .Y(n_1294) );
AOI22xp33_ASAP7_75t_SL g1295 ( .A1(n_1221), .A2(n_1219), .B1(n_1194), .B2(n_1206), .Y(n_1295) );
OR2x2_ASAP7_75t_L g1296 ( .A(n_1260), .B(n_1203), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1183), .Y(n_1297) );
NOR2x1_ASAP7_75t_L g1298 ( .A(n_1177), .B(n_1180), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1241), .B(n_1242), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1241), .B(n_1242), .Y(n_1300) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1160), .Y(n_1301) );
INVx3_ASAP7_75t_L g1302 ( .A(n_1186), .Y(n_1302) );
INVx2_ASAP7_75t_SL g1303 ( .A(n_1244), .Y(n_1303) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1161), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1228), .B(n_1171), .Y(n_1305) );
HB1xp67_ASAP7_75t_L g1306 ( .A(n_1206), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1249), .B(n_1262), .Y(n_1307) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1249), .B(n_1262), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1243), .B(n_1245), .Y(n_1309) );
OR2x2_ASAP7_75t_L g1310 ( .A(n_1246), .B(n_1211), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1210), .B(n_1212), .Y(n_1311) );
NAND3xp33_ASAP7_75t_L g1312 ( .A(n_1173), .B(n_1232), .C(n_1256), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1162), .Y(n_1313) );
INVx2_ASAP7_75t_SL g1314 ( .A(n_1244), .Y(n_1314) );
AND2x4_ASAP7_75t_SL g1315 ( .A(n_1177), .B(n_1191), .Y(n_1315) );
BUFx2_ASAP7_75t_L g1316 ( .A(n_1167), .Y(n_1316) );
AND2x4_ASAP7_75t_SL g1317 ( .A(n_1177), .B(n_1191), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1166), .Y(n_1318) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1170), .B(n_1172), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1178), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1179), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g1322 ( .A1(n_1257), .A2(n_1235), .B1(n_1264), .B2(n_1194), .Y(n_1322) );
OR2x2_ASAP7_75t_SL g1323 ( .A(n_1175), .B(n_1185), .Y(n_1323) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1184), .Y(n_1324) );
INVxp67_ASAP7_75t_SL g1325 ( .A(n_1194), .Y(n_1325) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1198), .Y(n_1326) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1258), .B(n_1199), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1200), .Y(n_1328) );
HB1xp67_ASAP7_75t_L g1329 ( .A(n_1214), .Y(n_1329) );
OR2x2_ASAP7_75t_L g1330 ( .A(n_1207), .B(n_1208), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1216), .Y(n_1331) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_1167), .Y(n_1332) );
AND2x2_ASAP7_75t_L g1333 ( .A(n_1263), .B(n_1270), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1224), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1234), .Y(n_1335) );
NOR2xp67_ASAP7_75t_L g1336 ( .A(n_1188), .B(n_1190), .Y(n_1336) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_1253), .A2(n_1233), .B1(n_1222), .B2(n_1192), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1273), .B(n_1267), .Y(n_1338) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1168), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1340 ( .A(n_1217), .B(n_1265), .Y(n_1340) );
BUFx2_ASAP7_75t_L g1341 ( .A(n_1167), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1236), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1217), .B(n_1272), .Y(n_1343) );
BUFx3_ASAP7_75t_L g1344 ( .A(n_1180), .Y(n_1344) );
BUFx2_ASAP7_75t_L g1345 ( .A(n_1175), .Y(n_1345) );
AND2x4_ASAP7_75t_L g1346 ( .A(n_1182), .B(n_1269), .Y(n_1346) );
AND2x4_ASAP7_75t_L g1347 ( .A(n_1182), .B(n_1269), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1215), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1227), .Y(n_1349) );
INVx1_ASAP7_75t_SL g1350 ( .A(n_1157), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1238), .Y(n_1351) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1185), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1230), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1209), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1209), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1209), .Y(n_1356) );
INVx4_ASAP7_75t_L g1357 ( .A(n_1261), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1272), .B(n_1250), .Y(n_1358) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1252), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1360 ( .A(n_1223), .B(n_1225), .Y(n_1360) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1229), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1269), .B(n_1165), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1363 ( .A(n_1218), .B(n_1248), .Y(n_1363) );
INVx1_ASAP7_75t_L g1364 ( .A(n_1229), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1165), .B(n_1163), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1163), .B(n_1280), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1299), .B(n_1280), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1329), .Y(n_1368) );
CKINVDCx20_ASAP7_75t_R g1369 ( .A(n_1282), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1297), .B(n_1239), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1300), .B(n_1276), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1351), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1319), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1345), .Y(n_1374) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1319), .Y(n_1375) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1339), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1377 ( .A(n_1300), .B(n_1276), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1307), .B(n_1164), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1308), .B(n_1169), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1330), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1287), .B(n_1190), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1292), .B(n_1202), .Y(n_1382) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1330), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1301), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1348), .B(n_1213), .Y(n_1385) );
AND2x4_ASAP7_75t_SL g1386 ( .A(n_1357), .B(n_1193), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1308), .B(n_1174), .Y(n_1387) );
OR2x2_ASAP7_75t_L g1388 ( .A(n_1296), .B(n_1275), .Y(n_1388) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1304), .Y(n_1389) );
INVx4_ASAP7_75t_L g1390 ( .A(n_1357), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1305), .B(n_1204), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1392 ( .A(n_1337), .B(n_1182), .Y(n_1392) );
AND2x4_ASAP7_75t_L g1393 ( .A(n_1346), .B(n_1254), .Y(n_1393) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_1346), .B(n_1254), .Y(n_1394) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1293), .B(n_1333), .Y(n_1395) );
NOR2xp33_ASAP7_75t_L g1396 ( .A(n_1285), .B(n_1266), .Y(n_1396) );
INVxp67_ASAP7_75t_L g1397 ( .A(n_1345), .Y(n_1397) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_1333), .B(n_1176), .Y(n_1398) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1359), .Y(n_1399) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1313), .Y(n_1400) );
OR2x2_ASAP7_75t_L g1401 ( .A(n_1310), .B(n_1205), .Y(n_1401) );
BUFx2_ASAP7_75t_L g1402 ( .A(n_1323), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1338), .B(n_1247), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1327), .B(n_1237), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_1331), .B(n_1274), .Y(n_1405) );
BUFx2_ASAP7_75t_L g1406 ( .A(n_1323), .Y(n_1406) );
INVx1_ASAP7_75t_L g1407 ( .A(n_1318), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1366), .B(n_1237), .Y(n_1408) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1320), .Y(n_1409) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1321), .Y(n_1410) );
INVx1_ASAP7_75t_SL g1411 ( .A(n_1282), .Y(n_1411) );
OAI21xp5_ASAP7_75t_L g1412 ( .A1(n_1312), .A2(n_1251), .B(n_1278), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1324), .Y(n_1413) );
BUFx2_ASAP7_75t_SL g1414 ( .A(n_1283), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1415 ( .A(n_1340), .B(n_1268), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g1416 ( .A1(n_1322), .A2(n_1251), .B1(n_1279), .B2(n_1191), .C(n_1193), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1340), .B(n_1181), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g1418 ( .A1(n_1295), .A2(n_1261), .B1(n_1226), .B2(n_1240), .Y(n_1418) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1334), .B(n_1240), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1358), .B(n_1343), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1421 ( .A(n_1360), .B(n_1240), .Y(n_1421) );
INVx2_ASAP7_75t_SL g1422 ( .A(n_1352), .Y(n_1422) );
INVxp67_ASAP7_75t_SL g1423 ( .A(n_1352), .Y(n_1423) );
INVx2_ASAP7_75t_SL g1424 ( .A(n_1283), .Y(n_1424) );
BUFx2_ASAP7_75t_L g1425 ( .A(n_1316), .Y(n_1425) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1359), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1420), .B(n_1362), .Y(n_1427) );
HB1xp67_ASAP7_75t_L g1428 ( .A(n_1422), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1371), .B(n_1365), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1430 ( .A(n_1371), .B(n_1289), .Y(n_1430) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1373), .B(n_1326), .Y(n_1431) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1399), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1377), .B(n_1289), .Y(n_1433) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1377), .B(n_1354), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1426), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1367), .B(n_1354), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_1375), .B(n_1328), .Y(n_1437) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1368), .Y(n_1438) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1380), .B(n_1335), .Y(n_1439) );
OAI21xp33_ASAP7_75t_SL g1440 ( .A1(n_1424), .A2(n_1357), .B(n_1303), .Y(n_1440) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1384), .Y(n_1441) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1376), .Y(n_1442) );
AND2x4_ASAP7_75t_L g1443 ( .A(n_1393), .B(n_1347), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1444 ( .A(n_1367), .B(n_1355), .Y(n_1444) );
AND2x4_ASAP7_75t_L g1445 ( .A(n_1393), .B(n_1347), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1389), .Y(n_1446) );
BUFx2_ASAP7_75t_L g1447 ( .A(n_1424), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_1403), .B(n_1355), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1403), .B(n_1356), .Y(n_1449) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1400), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1451 ( .A(n_1395), .B(n_1286), .Y(n_1451) );
NOR2x1_ASAP7_75t_L g1452 ( .A(n_1369), .B(n_1298), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_1395), .B(n_1361), .Y(n_1453) );
INVx1_ASAP7_75t_SL g1454 ( .A(n_1369), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1407), .Y(n_1455) );
OR2x2_ASAP7_75t_L g1456 ( .A(n_1398), .B(n_1361), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1457 ( .A1(n_1418), .A2(n_1325), .B1(n_1316), .B2(n_1332), .Y(n_1457) );
NAND2xp5_ASAP7_75t_L g1458 ( .A(n_1383), .B(n_1342), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1409), .Y(n_1459) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1410), .Y(n_1460) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1372), .B(n_1349), .Y(n_1461) );
INVx1_ASAP7_75t_L g1462 ( .A(n_1413), .Y(n_1462) );
INVx2_ASAP7_75t_SL g1463 ( .A(n_1422), .Y(n_1463) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1405), .B(n_1364), .Y(n_1464) );
INVx1_ASAP7_75t_SL g1465 ( .A(n_1411), .Y(n_1465) );
INVx1_ASAP7_75t_SL g1466 ( .A(n_1414), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1370), .Y(n_1467) );
OR2x2_ASAP7_75t_L g1468 ( .A(n_1398), .B(n_1364), .Y(n_1468) );
NAND2xp5_ASAP7_75t_L g1469 ( .A(n_1378), .B(n_1284), .Y(n_1469) );
INVx2_ASAP7_75t_SL g1470 ( .A(n_1386), .Y(n_1470) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1415), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g1472 ( .A(n_1374), .Y(n_1472) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1415), .Y(n_1473) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1388), .B(n_1309), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1378), .Y(n_1475) );
HB1xp67_ASAP7_75t_L g1476 ( .A(n_1397), .Y(n_1476) );
AND2x2_ASAP7_75t_L g1477 ( .A(n_1427), .B(n_1408), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1467), .B(n_1417), .Y(n_1478) );
INVx2_ASAP7_75t_L g1479 ( .A(n_1442), .Y(n_1479) );
XNOR2x2_ASAP7_75t_L g1480 ( .A(n_1452), .B(n_1466), .Y(n_1480) );
BUFx2_ASAP7_75t_L g1481 ( .A(n_1440), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1482 ( .A(n_1427), .B(n_1408), .Y(n_1482) );
INVx1_ASAP7_75t_SL g1483 ( .A(n_1454), .Y(n_1483) );
NAND2xp5_ASAP7_75t_SL g1484 ( .A(n_1470), .B(n_1402), .Y(n_1484) );
AND2x4_ASAP7_75t_L g1485 ( .A(n_1443), .B(n_1393), .Y(n_1485) );
NOR2x1_ASAP7_75t_L g1486 ( .A(n_1447), .B(n_1414), .Y(n_1486) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1429), .B(n_1404), .Y(n_1487) );
NOR2xp33_ASAP7_75t_L g1488 ( .A(n_1465), .B(n_1396), .Y(n_1488) );
INVxp67_ASAP7_75t_L g1489 ( .A(n_1447), .Y(n_1489) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_1451), .B(n_1388), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1429), .B(n_1404), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1430), .B(n_1379), .Y(n_1492) );
INVx3_ASAP7_75t_L g1493 ( .A(n_1443), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1494 ( .A(n_1430), .B(n_1379), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1432), .Y(n_1495) );
AOI21x1_ASAP7_75t_L g1496 ( .A1(n_1457), .A2(n_1277), .B(n_1406), .Y(n_1496) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1435), .Y(n_1497) );
O2A1O1Ixp5_ASAP7_75t_SL g1498 ( .A1(n_1438), .A2(n_1353), .B(n_1412), .C(n_1294), .Y(n_1498) );
INVxp67_ASAP7_75t_SL g1499 ( .A(n_1428), .Y(n_1499) );
INVx1_ASAP7_75t_SL g1500 ( .A(n_1470), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1441), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1433), .B(n_1387), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1441), .Y(n_1503) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1451), .B(n_1401), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1433), .B(n_1387), .Y(n_1505) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1446), .Y(n_1506) );
INVx1_ASAP7_75t_SL g1507 ( .A(n_1456), .Y(n_1507) );
INVx2_ASAP7_75t_L g1508 ( .A(n_1479), .Y(n_1508) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1490), .Y(n_1509) );
OAI21xp5_ASAP7_75t_SL g1510 ( .A1(n_1481), .A2(n_1317), .B(n_1315), .Y(n_1510) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1490), .Y(n_1511) );
INVx2_ASAP7_75t_L g1512 ( .A(n_1479), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1507), .B(n_1448), .Y(n_1513) );
INVx1_ASAP7_75t_L g1514 ( .A(n_1501), .Y(n_1514) );
OAI22xp5_ASAP7_75t_L g1515 ( .A1(n_1481), .A2(n_1402), .B1(n_1406), .B2(n_1474), .Y(n_1515) );
INVx2_ASAP7_75t_L g1516 ( .A(n_1479), .Y(n_1516) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1504), .B(n_1471), .Y(n_1517) );
OR2x2_ASAP7_75t_L g1518 ( .A(n_1504), .B(n_1471), .Y(n_1518) );
INVxp67_ASAP7_75t_L g1519 ( .A(n_1488), .Y(n_1519) );
XNOR2x2_ASAP7_75t_L g1520 ( .A(n_1480), .B(n_1416), .Y(n_1520) );
OA21x2_ASAP7_75t_L g1521 ( .A1(n_1484), .A2(n_1464), .B(n_1449), .Y(n_1521) );
INVxp67_ASAP7_75t_L g1522 ( .A(n_1499), .Y(n_1522) );
OAI21xp5_ASAP7_75t_L g1523 ( .A1(n_1486), .A2(n_1423), .B(n_1303), .Y(n_1523) );
NOR2xp33_ASAP7_75t_L g1524 ( .A(n_1483), .B(n_1472), .Y(n_1524) );
AND2x4_ASAP7_75t_L g1525 ( .A(n_1486), .B(n_1443), .Y(n_1525) );
HB1xp67_ASAP7_75t_L g1526 ( .A(n_1489), .Y(n_1526) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1501), .Y(n_1527) );
AOI22xp5_ASAP7_75t_L g1528 ( .A1(n_1500), .A2(n_1448), .B1(n_1449), .B2(n_1444), .Y(n_1528) );
AO22x2_ASAP7_75t_L g1529 ( .A1(n_1493), .A2(n_1463), .B1(n_1459), .B2(n_1455), .Y(n_1529) );
O2A1O1Ixp33_ASAP7_75t_L g1530 ( .A1(n_1478), .A2(n_1476), .B(n_1385), .C(n_1391), .Y(n_1530) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1503), .Y(n_1531) );
INVx1_ASAP7_75t_L g1532 ( .A(n_1503), .Y(n_1532) );
AOI21xp33_ASAP7_75t_L g1533 ( .A1(n_1506), .A2(n_1350), .B(n_1255), .Y(n_1533) );
AOI22xp5_ASAP7_75t_L g1534 ( .A1(n_1485), .A2(n_1434), .B1(n_1436), .B2(n_1444), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1514), .Y(n_1535) );
OAI22xp5_ASAP7_75t_L g1536 ( .A1(n_1510), .A2(n_1493), .B1(n_1485), .B2(n_1390), .Y(n_1536) );
AOI21xp33_ASAP7_75t_SL g1537 ( .A1(n_1510), .A2(n_1480), .B(n_1493), .Y(n_1537) );
OAI31xp33_ASAP7_75t_L g1538 ( .A1(n_1515), .A2(n_1493), .A3(n_1485), .B(n_1386), .Y(n_1538) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_1509), .B(n_1506), .Y(n_1539) );
OAI21xp33_ASAP7_75t_L g1540 ( .A1(n_1515), .A2(n_1496), .B(n_1482), .Y(n_1540) );
OAI21xp33_ASAP7_75t_L g1541 ( .A1(n_1529), .A2(n_1496), .B(n_1482), .Y(n_1541) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1527), .Y(n_1542) );
XOR2x2_ASAP7_75t_SL g1543 ( .A(n_1520), .B(n_1485), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1544 ( .A1(n_1524), .A2(n_1434), .B1(n_1436), .B2(n_1445), .Y(n_1544) );
NOR4xp25_ASAP7_75t_SL g1545 ( .A(n_1533), .B(n_1332), .C(n_1341), .D(n_1425), .Y(n_1545) );
NAND2xp33_ASAP7_75t_SL g1546 ( .A(n_1525), .B(n_1220), .Y(n_1546) );
OAI221xp5_ASAP7_75t_L g1547 ( .A1(n_1523), .A2(n_1463), .B1(n_1392), .B2(n_1453), .C(n_1458), .Y(n_1547) );
AOI222xp33_ASAP7_75t_L g1548 ( .A1(n_1519), .A2(n_1439), .B1(n_1431), .B2(n_1437), .C1(n_1462), .C2(n_1446), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1531), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1532), .Y(n_1550) );
AOI22xp5_ASAP7_75t_L g1551 ( .A1(n_1511), .A2(n_1445), .B1(n_1473), .B2(n_1475), .Y(n_1551) );
A2O1A1Ixp33_ASAP7_75t_L g1552 ( .A1(n_1530), .A2(n_1315), .B(n_1317), .C(n_1502), .Y(n_1552) );
AOI31xp33_ASAP7_75t_L g1553 ( .A1(n_1523), .A2(n_1314), .A3(n_1290), .B(n_1494), .Y(n_1553) );
INVx2_ASAP7_75t_L g1554 ( .A(n_1529), .Y(n_1554) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_1522), .B(n_1487), .Y(n_1555) );
AOI211xp5_ASAP7_75t_L g1556 ( .A1(n_1533), .A2(n_1220), .B(n_1445), .C(n_1279), .Y(n_1556) );
OAI22xp33_ASAP7_75t_L g1557 ( .A1(n_1521), .A2(n_1390), .B1(n_1474), .B2(n_1341), .Y(n_1557) );
OAI222xp33_ASAP7_75t_L g1558 ( .A1(n_1528), .A2(n_1505), .B1(n_1502), .B2(n_1492), .C1(n_1494), .C2(n_1390), .Y(n_1558) );
AOI21xp33_ASAP7_75t_L g1559 ( .A1(n_1521), .A2(n_1381), .B(n_1291), .Y(n_1559) );
AOI22xp33_ASAP7_75t_SL g1560 ( .A1(n_1525), .A2(n_1526), .B1(n_1505), .B2(n_1394), .Y(n_1560) );
AOI211x1_ASAP7_75t_SL g1561 ( .A1(n_1513), .A2(n_1382), .B(n_1461), .C(n_1363), .Y(n_1561) );
OAI21xp33_ASAP7_75t_L g1562 ( .A1(n_1534), .A2(n_1477), .B(n_1491), .Y(n_1562) );
OAI211xp5_ASAP7_75t_L g1563 ( .A1(n_1517), .A2(n_1425), .B(n_1421), .C(n_1453), .Y(n_1563) );
AOI21xp5_ASAP7_75t_L g1564 ( .A1(n_1518), .A2(n_1314), .B(n_1290), .Y(n_1564) );
AOI21xp5_ASAP7_75t_L g1565 ( .A1(n_1508), .A2(n_1469), .B(n_1468), .Y(n_1565) );
NOR2xp33_ASAP7_75t_SL g1566 ( .A(n_1512), .B(n_1344), .Y(n_1566) );
AND3x1_ASAP7_75t_L g1567 ( .A(n_1516), .B(n_1477), .C(n_1491), .Y(n_1567) );
OAI211xp5_ASAP7_75t_L g1568 ( .A1(n_1537), .A2(n_1540), .B(n_1546), .C(n_1538), .Y(n_1568) );
NAND4xp25_ASAP7_75t_L g1569 ( .A(n_1556), .B(n_1543), .C(n_1552), .D(n_1536), .Y(n_1569) );
NOR2x1_ASAP7_75t_L g1570 ( .A(n_1557), .B(n_1536), .Y(n_1570) );
AOI21xp33_ASAP7_75t_R g1571 ( .A1(n_1554), .A2(n_1541), .B(n_1539), .Y(n_1571) );
NAND4xp25_ASAP7_75t_L g1572 ( .A(n_1561), .B(n_1560), .C(n_1562), .D(n_1548), .Y(n_1572) );
AND2x4_ASAP7_75t_L g1573 ( .A(n_1567), .B(n_1564), .Y(n_1573) );
XNOR2x1_ASAP7_75t_L g1574 ( .A(n_1271), .B(n_1557), .Y(n_1574) );
NOR2xp33_ASAP7_75t_L g1575 ( .A(n_1558), .B(n_1555), .Y(n_1575) );
OAI211xp5_ASAP7_75t_L g1576 ( .A1(n_1545), .A2(n_1559), .B(n_1547), .C(n_1563), .Y(n_1576) );
AOI211x1_ASAP7_75t_L g1577 ( .A1(n_1553), .A2(n_1565), .B(n_1539), .C(n_1542), .Y(n_1577) );
NAND4xp25_ASAP7_75t_L g1578 ( .A(n_1569), .B(n_1577), .C(n_1568), .D(n_1570), .Y(n_1578) );
NOR3xp33_ASAP7_75t_L g1579 ( .A(n_1576), .B(n_1572), .C(n_1575), .Y(n_1579) );
NOR3xp33_ASAP7_75t_L g1580 ( .A(n_1573), .B(n_1193), .C(n_1549), .Y(n_1580) );
INVx2_ASAP7_75t_L g1581 ( .A(n_1574), .Y(n_1581) );
NOR2xp67_ASAP7_75t_L g1582 ( .A(n_1571), .B(n_1544), .Y(n_1582) );
NOR3xp33_ASAP7_75t_L g1583 ( .A(n_1568), .B(n_1550), .C(n_1535), .Y(n_1583) );
NAND4xp25_ASAP7_75t_L g1584 ( .A(n_1579), .B(n_1566), .C(n_1551), .D(n_1344), .Y(n_1584) );
NAND4xp25_ASAP7_75t_L g1585 ( .A(n_1578), .B(n_1336), .C(n_1311), .D(n_1394), .Y(n_1585) );
NAND4xp25_ASAP7_75t_L g1586 ( .A(n_1582), .B(n_1581), .C(n_1583), .D(n_1580), .Y(n_1586) );
INVx2_ASAP7_75t_SL g1587 ( .A(n_1581), .Y(n_1587) );
INVx3_ASAP7_75t_L g1588 ( .A(n_1587), .Y(n_1588) );
OR2x2_ASAP7_75t_L g1589 ( .A(n_1584), .B(n_1586), .Y(n_1589) );
HB1xp67_ASAP7_75t_L g1590 ( .A(n_1585), .Y(n_1590) );
OAI22xp5_ASAP7_75t_SL g1591 ( .A1(n_1589), .A2(n_1261), .B1(n_1281), .B2(n_1460), .Y(n_1591) );
NAND3xp33_ASAP7_75t_L g1592 ( .A(n_1588), .B(n_1498), .C(n_1201), .Y(n_1592) );
NAND2xp5_ASAP7_75t_L g1593 ( .A(n_1590), .B(n_1450), .Y(n_1593) );
O2A1O1Ixp33_ASAP7_75t_SL g1594 ( .A1(n_1593), .A2(n_1460), .B(n_1462), .C(n_1419), .Y(n_1594) );
XOR2xp5_ASAP7_75t_L g1595 ( .A(n_1591), .B(n_1306), .Y(n_1595) );
AOI21xp5_ASAP7_75t_L g1596 ( .A1(n_1592), .A2(n_1495), .B(n_1497), .Y(n_1596) );
AOI21xp5_ASAP7_75t_L g1597 ( .A1(n_1595), .A2(n_1594), .B(n_1596), .Y(n_1597) );
OR2x6_ASAP7_75t_L g1598 ( .A(n_1597), .B(n_1201), .Y(n_1598) );
OAI21xp5_ASAP7_75t_L g1599 ( .A1(n_1598), .A2(n_1288), .B(n_1302), .Y(n_1599) );
AOI21xp5_ASAP7_75t_L g1600 ( .A1(n_1599), .A2(n_1231), .B(n_1197), .Y(n_1600) );
endmodule