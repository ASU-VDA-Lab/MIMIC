module real_jpeg_27467_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_187;
wire n_75;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_0),
.A2(n_28),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_34),
.B1(n_44),
.B2(n_45),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_1),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_2),
.A2(n_62),
.B1(n_63),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_2),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_76),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_2),
.A2(n_44),
.B1(n_45),
.B2(n_76),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_2),
.A2(n_28),
.B1(n_33),
.B2(n_76),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_3),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g90 ( 
.A1(n_3),
.A2(n_59),
.B(n_63),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_89),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_61),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_45),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_45),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_78),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_3),
.A2(n_26),
.B1(n_199),
.B2(n_203),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_3),
.A2(n_62),
.B(n_215),
.Y(n_214)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_5),
.A2(n_62),
.B1(n_63),
.B2(n_84),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_5),
.A2(n_44),
.B1(n_45),
.B2(n_84),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_5),
.A2(n_28),
.B1(n_33),
.B2(n_84),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_6),
.A2(n_28),
.B1(n_33),
.B2(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_6),
.A2(n_51),
.B1(n_62),
.B2(n_63),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_8),
.A2(n_28),
.B1(n_33),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_8),
.Y(n_100)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_10),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_10),
.A2(n_43),
.B1(n_62),
.B2(n_63),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_10),
.A2(n_28),
.B1(n_33),
.B2(n_43),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_11),
.A2(n_28),
.B1(n_33),
.B2(n_48),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_11),
.A2(n_33),
.A3(n_45),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_12),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_62),
.B1(n_63),
.B2(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_12),
.A2(n_28),
.B1(n_33),
.B2(n_67),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_12),
.A2(n_44),
.B1(n_45),
.B2(n_67),
.Y(n_219)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_14),
.B(n_62),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_44),
.B1(n_45),
.B2(n_72),
.Y(n_74)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_14),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_28),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_15),
.A2(n_39),
.B1(n_44),
.B2(n_45),
.Y(n_111)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_17),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g135 ( 
.A1(n_17),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_17),
.A2(n_44),
.B1(n_45),
.B2(n_55),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_17),
.A2(n_28),
.B1(n_33),
.B2(n_55),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_123),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_103),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_22),
.B(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_79),
.C(n_97),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_23),
.B(n_97),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_52),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_24),
.B(n_53),
.C(n_68),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_25),
.B(n_40),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_26),
.A2(n_37),
.B1(n_38),
.B2(n_99),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_26),
.A2(n_35),
.B(n_99),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_26),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_26),
.A2(n_37),
.B1(n_193),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_26),
.A2(n_187),
.B1(n_188),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_27),
.A2(n_32),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_27),
.A2(n_36),
.B1(n_92),
.B2(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_27),
.A2(n_36),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_28),
.B(n_48),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_28),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_SL g188 ( 
.A(n_36),
.Y(n_188)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_42),
.A2(n_109),
.B1(n_112),
.B2(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g223 ( 
.A1(n_44),
.A2(n_62),
.A3(n_216),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_45),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_47),
.B1(n_50),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_46),
.A2(n_47),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_46),
.A2(n_47),
.B1(n_173),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_46),
.A2(n_47),
.B1(n_140),
.B2(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_47),
.B(n_89),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_68),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_61),
.B2(n_66),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_54),
.Y(n_86)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_65),
.B(n_89),
.C(n_90),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_58),
.A2(n_61),
.B1(n_66),
.B2(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_58),
.A2(n_61),
.B1(n_83),
.B2(n_137),
.Y(n_136)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_61),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_70)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_63),
.B(n_89),
.Y(n_216)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_75),
.B1(n_77),
.B2(n_78),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_69),
.A2(n_77),
.B1(n_78),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_69),
.A2(n_78),
.B1(n_135),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_74),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_70),
.A2(n_74),
.B1(n_95),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_70),
.A2(n_74),
.B1(n_155),
.B2(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_87),
.C(n_94),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_94),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_87),
.B(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_89),
.B(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_101),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_121),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_113),
.B2(n_114),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_109),
.A2(n_112),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx24_ASAP7_75t_SL g253 ( 
.A(n_115),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_118),
.CI(n_120),
.CON(n_115),
.SN(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_160),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_143),
.B(n_159),
.Y(n_125)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_141),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_141),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.C(n_131),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_131),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.C(n_138),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_146),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_151),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_147),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_150),
.Y(n_251)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_153),
.B(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_156),
.B(n_158),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_157),
.Y(n_229)
);

NOR3xp33_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.C(n_163),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_247),
.B(n_252),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_233),
.B(n_246),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_209),
.B(n_232),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_189),
.B(n_208),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_178),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_168),
.B(n_178),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_174),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_175),
.Y(n_195)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_172),
.Y(n_176)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_184),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_186),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_196),
.B(n_207),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_191),
.B(n_195),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_201),
.B(n_206),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_200),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_210),
.B(n_211),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_212),
.A2(n_222),
.B1(n_230),
.B2(n_231),
.Y(n_211)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_221),
.Y(n_212)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_217),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_217),
.B(n_221),
.C(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_228),
.Y(n_241)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_224),
.Y(n_227)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_234),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_242),
.C(n_244),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_244),
.B2(n_245),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);


endmodule