module fake_jpeg_2422_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_31),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_28),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_29),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_48),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_31),
.B1(n_33),
.B2(n_30),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_29),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_56),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_53),
.B1(n_43),
.B2(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_1),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_15),
.Y(n_67)
);

OAI22x1_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_13),
.B1(n_22),
.B2(n_20),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2x1_ASAP7_75t_SL g56 ( 
.A(n_47),
.B(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_3),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_5),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_67),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_68),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_55),
.B1(n_7),
.B2(n_8),
.Y(n_71)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_74),
.B1(n_76),
.B2(n_70),
.C(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_6),
.B(n_8),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_10),
.B(n_16),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g81 ( 
.A(n_75),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_77),
.B(n_9),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_83),
.B(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_71),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_79),
.C(n_80),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_88),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_90),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_86),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

OA21x2_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_85),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_18),
.Y(n_95)
);


endmodule