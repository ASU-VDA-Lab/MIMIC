module fake_jpeg_12986_n_193 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_193);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx24_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_10),
.Y(n_56)
);

INVx2_ASAP7_75t_R g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_84),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_89),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_68),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_77),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_57),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_98),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_57),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_63),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_55),
.C(n_53),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_75),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_78),
.B1(n_74),
.B2(n_79),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_104),
.A2(n_81),
.B1(n_79),
.B2(n_72),
.Y(n_108)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_107),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_120),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_104),
.A2(n_91),
.B1(n_81),
.B2(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_113),
.B1(n_70),
.B2(n_69),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_119),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_102),
.Y(n_112)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_73),
.B1(n_66),
.B2(n_67),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_71),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_122),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_102),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_124),
.Y(n_133)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_65),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_73),
.B1(n_67),
.B2(n_62),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_61),
.B1(n_65),
.B2(n_2),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_136),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_140),
.B1(n_142),
.B2(n_150),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g132 ( 
.A(n_117),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_143),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_129),
.B(n_146),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_139),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_61),
.B1(n_1),
.B2(n_2),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_0),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_4),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_151),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_5),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_163),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_8),
.B(n_9),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_160),
.B(n_155),
.Y(n_178)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_11),
.C(n_12),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_168),
.B1(n_50),
.B2(n_34),
.Y(n_175)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_157),
.B(n_161),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g158 ( 
.A(n_144),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_134),
.A2(n_16),
.B(n_17),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_23),
.B(n_25),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_149),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_166),
.Y(n_170)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_167),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_157),
.A2(n_140),
.B1(n_141),
.B2(n_35),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_174),
.B(n_175),
.Y(n_180)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_171),
.B(n_165),
.C(n_154),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_179),
.B(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_159),
.C(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_162),
.B(n_153),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_178),
.B1(n_174),
.B2(n_170),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_184),
.A2(n_183),
.B1(n_176),
.B2(n_169),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_184),
.C(n_180),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_185),
.A3(n_167),
.B1(n_172),
.B2(n_43),
.C1(n_45),
.C2(n_47),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_33),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_36),
.C(n_41),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_48),
.Y(n_193)
);


endmodule