module fake_jpeg_12772_n_91 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_10),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_32),
.Y(n_35)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_14),
.B1(n_17),
.B2(n_21),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_13),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_28),
.A2(n_13),
.B1(n_18),
.B2(n_32),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_41),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_11),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_26),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_23),
.B(n_16),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_53),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_23),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_52),
.B(n_15),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_39),
.B(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_51),
.A2(n_45),
.B1(n_44),
.B2(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_36),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_48),
.B1(n_53),
.B2(n_40),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_36),
.B1(n_43),
.B2(n_29),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_54),
.A2(n_36),
.B1(n_43),
.B2(n_25),
.Y(n_59)
);

AOI21x1_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_69),
.B(n_70),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_43),
.Y(n_65)
);

A2O1A1O1Ixp25_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_63),
.B(n_62),
.C(n_61),
.D(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_56),
.B(n_19),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_68),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_63),
.C(n_61),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_78),
.B(n_79),
.Y(n_83)
);

AO221x1_ASAP7_75t_L g80 ( 
.A1(n_72),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_81),
.B(n_82),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_74),
.B1(n_67),
.B2(n_71),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_82),
.A2(n_73),
.B(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_83),
.A2(n_71),
.B(n_75),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_SL g87 ( 
.A(n_84),
.B(n_77),
.C(n_5),
.Y(n_87)
);

AOI321xp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_3),
.A3(n_6),
.B1(n_7),
.B2(n_19),
.C(n_42),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_3),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_88),
.Y(n_91)
);


endmodule