module fake_netlist_6_1370_n_1674 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1674);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1674;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_90),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_94),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_29),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_26),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_69),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_135),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_30),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_46),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_38),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_70),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_20),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_125),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_73),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_103),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_17),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_129),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_82),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_23),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_124),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVxp33_ASAP7_75t_SL g200 ( 
.A(n_75),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_157),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_62),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_110),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_93),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_165),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_49),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_30),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_17),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_131),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_56),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_97),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_6),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_81),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_171),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_145),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_89),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_99),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_84),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_108),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_35),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_18),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_19),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_74),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_116),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_42),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_154),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_67),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_14),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_167),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_123),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_50),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_59),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_118),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_32),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_7),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_105),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_166),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_10),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_147),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_144),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_15),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_11),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_168),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_43),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_83),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_107),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_96),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_87),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g259 ( 
.A(n_55),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_138),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_160),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_35),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_52),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_153),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_61),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_79),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_53),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_100),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_128),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_152),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_15),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_146),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_28),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_41),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_25),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_27),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_106),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_161),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_112),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_3),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_95),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_20),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_139),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_134),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_130),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_40),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_162),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_114),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_49),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_1),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_53),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

CKINVDCx11_ASAP7_75t_R g296 ( 
.A(n_77),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_34),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_76),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_41),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_58),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_46),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_68),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_21),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_155),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_52),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_85),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_142),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_47),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_102),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_104),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_158),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_64),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_148),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_169),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_98),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_149),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_51),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_42),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_78),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_141),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_34),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_163),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_43),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_16),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_13),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_6),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_25),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_8),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_5),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_66),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_27),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_57),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g337 ( 
.A(n_38),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_156),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_121),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_18),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_64),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_120),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_92),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_37),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_202),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_297),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_259),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_221),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_213),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_259),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_225),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_259),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_259),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_205),
.B(n_0),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_259),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_223),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_211),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_259),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_208),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_208),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_236),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_256),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_259),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_259),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_229),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_192),
.B(n_1),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_231),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_176),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_298),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_331),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_192),
.B(n_2),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_221),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_221),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_331),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_234),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_296),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_240),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_277),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_199),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_277),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_214),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_173),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_215),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_179),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_200),
.B(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_183),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_217),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_243),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_309),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_241),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_216),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_219),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_218),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_250),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_263),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_244),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_266),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_273),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_243),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_284),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_224),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_276),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_284),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_247),
.Y(n_407)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_176),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_340),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_199),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_251),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_226),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_295),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_252),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_303),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_261),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_193),
.B(n_4),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_264),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_308),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_326),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_335),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_253),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_182),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_193),
.B(n_4),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_222),
.B(n_5),
.Y(n_426)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_182),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_187),
.Y(n_428)
);

OR2x2_ASAP7_75t_L g429 ( 
.A(n_340),
.B(n_8),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_227),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_291),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_346),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_383),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_373),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_360),
.B(n_291),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_385),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_389),
.Y(n_442)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_359),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_391),
.Y(n_445)
);

INVxp33_ASAP7_75t_L g446 ( 
.A(n_357),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_359),
.B(n_249),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_353),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_345),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_375),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_375),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_353),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_394),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_347),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_404),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_391),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_358),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_358),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_347),
.B(n_172),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_423),
.B(n_249),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_351),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_391),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_350),
.Y(n_464)
);

AND2x4_ASAP7_75t_L g465 ( 
.A(n_350),
.B(n_302),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_412),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_364),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_352),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_L g469 ( 
.A(n_346),
.B(n_187),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_356),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_355),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_430),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_377),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_363),
.B(n_302),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_431),
.B(n_316),
.Y(n_479)
);

CKINVDCx8_ASAP7_75t_R g480 ( 
.A(n_380),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_403),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_403),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_379),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g485 ( 
.A(n_365),
.B(n_367),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_406),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_381),
.B(n_316),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_365),
.B(n_175),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_406),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_409),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_409),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_367),
.Y(n_492)
);

OA21x2_ASAP7_75t_L g493 ( 
.A1(n_417),
.A2(n_181),
.B(n_178),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_429),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_429),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_366),
.B(n_191),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_384),
.Y(n_497)
);

AND2x2_ASAP7_75t_SL g498 ( 
.A(n_387),
.B(n_309),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_R g499 ( 
.A(n_376),
.B(n_228),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_361),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_386),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_388),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_393),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_SL g504 ( 
.A1(n_498),
.A2(n_410),
.B1(n_186),
.B2(n_230),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_498),
.B(n_354),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_455),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_498),
.B(n_309),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_376),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_464),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_378),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_464),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_438),
.B(n_408),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_444),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g514 ( 
.A(n_494),
.B(n_495),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_494),
.A2(n_425),
.B1(n_426),
.B2(n_400),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_494),
.B(n_378),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_392),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_448),
.Y(n_519)
);

INVxp33_ASAP7_75t_L g520 ( 
.A(n_446),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_488),
.B(n_368),
.Y(n_521)
);

BUFx10_ASAP7_75t_L g522 ( 
.A(n_492),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_392),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_495),
.B(n_309),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_495),
.B(n_395),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_449),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_398),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_424),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_443),
.B(n_428),
.Y(n_532)
);

BUFx10_ASAP7_75t_L g533 ( 
.A(n_437),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_444),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_482),
.B(n_398),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_493),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_479),
.B(n_427),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_471),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_493),
.A2(n_400),
.B1(n_371),
.B2(n_427),
.Y(n_540)
);

INVx4_ASAP7_75t_SL g541 ( 
.A(n_471),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_493),
.A2(n_419),
.B1(n_396),
.B2(n_397),
.Y(n_542)
);

NAND3xp33_ASAP7_75t_L g543 ( 
.A(n_485),
.B(n_411),
.C(n_407),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_465),
.B(n_310),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_453),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g546 ( 
.A(n_484),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g547 ( 
.A(n_469),
.B(n_411),
.C(n_407),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_447),
.B(n_348),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_479),
.B(n_399),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_458),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_465),
.B(n_310),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_468),
.B(n_414),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_496),
.Y(n_553)
);

NAND2x1p5_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_245),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_471),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_458),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_458),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_459),
.Y(n_558)
);

INVx1_ASAP7_75t_SL g559 ( 
.A(n_462),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_479),
.B(n_401),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_465),
.B(n_310),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_444),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_465),
.B(n_310),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_499),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_470),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_503),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_452),
.Y(n_567)
);

INVx5_ASAP7_75t_L g568 ( 
.A(n_444),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_477),
.B(n_413),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_460),
.B(n_474),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_460),
.B(n_416),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_474),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_474),
.B(n_310),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_474),
.B(n_416),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_418),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_500),
.Y(n_577)
);

AO22x2_ASAP7_75t_L g578 ( 
.A1(n_496),
.A2(n_237),
.B1(n_324),
.B2(n_337),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_461),
.A2(n_422),
.B1(n_421),
.B2(n_420),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_445),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_475),
.B(n_418),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_434),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_440),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_459),
.Y(n_584)
);

INVx4_ASAP7_75t_SL g585 ( 
.A(n_445),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_475),
.B(n_194),
.Y(n_586)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_432),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_459),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_L g589 ( 
.A1(n_487),
.A2(n_415),
.B1(n_405),
.B2(n_242),
.Y(n_589)
);

NAND3xp33_ASAP7_75t_L g590 ( 
.A(n_432),
.B(n_278),
.C(n_275),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_497),
.A2(n_280),
.B1(n_195),
.B2(n_269),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_434),
.B(n_201),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_475),
.B(n_206),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_450),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_451),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_497),
.B(n_374),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_497),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_435),
.Y(n_598)
);

AO22x2_ASAP7_75t_L g599 ( 
.A1(n_435),
.A2(n_220),
.B1(n_239),
.B2(n_246),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_440),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_445),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_436),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_477),
.B(n_372),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_501),
.B(n_362),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_501),
.B(n_255),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_502),
.B(n_282),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_440),
.B(n_232),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_433),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_436),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_501),
.A2(n_290),
.B1(n_325),
.B2(n_322),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_439),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_475),
.B(n_262),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_481),
.B(n_199),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_445),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_445),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_457),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_502),
.B(n_481),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_502),
.Y(n_618)
);

AOI22xp33_ASAP7_75t_L g619 ( 
.A1(n_491),
.A2(n_265),
.B1(n_306),
.B2(n_338),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_440),
.B(n_233),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_441),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_L g623 ( 
.A1(n_491),
.A2(n_288),
.B1(n_258),
.B2(n_283),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_442),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_457),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_454),
.A2(n_369),
.B1(n_343),
.B2(n_342),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_441),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_483),
.B(n_174),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_451),
.B(n_235),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_531),
.A2(n_491),
.B(n_490),
.C(n_489),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_576),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_508),
.B(n_480),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_520),
.B(n_603),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_505),
.B(n_475),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_SL g635 ( 
.A(n_564),
.B(n_480),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_507),
.A2(n_312),
.B1(n_328),
.B2(n_314),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_521),
.B(n_174),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_527),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_510),
.B(n_177),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_505),
.B(n_476),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_517),
.A2(n_238),
.B1(n_248),
.B2(n_257),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_518),
.B(n_456),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_506),
.B(n_476),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_509),
.B(n_511),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_514),
.B(n_260),
.Y(n_645)
);

BUFx8_ASAP7_75t_L g646 ( 
.A(n_608),
.Y(n_646)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_520),
.Y(n_647)
);

AOI221xp5_ASAP7_75t_L g648 ( 
.A1(n_578),
.A2(n_320),
.B1(n_344),
.B2(n_268),
.C(n_196),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_524),
.B(n_466),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_529),
.B(n_472),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_512),
.B(n_180),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_532),
.B(n_180),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_606),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_535),
.B(n_478),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_594),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_540),
.B(n_185),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_569),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_554),
.B(n_185),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_597),
.B(n_478),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_531),
.B(n_271),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_597),
.B(n_457),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_512),
.B(n_188),
.Y(n_662)
);

AND2x6_ASAP7_75t_SL g663 ( 
.A(n_536),
.B(n_184),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_618),
.B(n_457),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_606),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_507),
.A2(n_254),
.B1(n_336),
.B2(n_207),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_537),
.A2(n_207),
.B1(n_344),
.B2(n_341),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_546),
.B(n_463),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_624),
.B(n_473),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_554),
.B(n_188),
.Y(n_670)
);

AND2x2_ASAP7_75t_SL g671 ( 
.A(n_531),
.B(n_483),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_552),
.B(n_189),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_595),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_605),
.B(n_463),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_617),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_575),
.B(n_190),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_548),
.B(n_190),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_617),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_551),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_L g681 ( 
.A1(n_515),
.A2(n_490),
.B1(n_489),
.B2(n_486),
.C(n_301),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_560),
.B(n_486),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_582),
.B(n_272),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_598),
.B(n_602),
.Y(n_684)
);

BUFx8_ASAP7_75t_L g685 ( 
.A(n_587),
.Y(n_685)
);

AO221x1_ASAP7_75t_L g686 ( 
.A1(n_578),
.A2(n_313),
.B1(n_288),
.B2(n_283),
.C(n_258),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_609),
.B(n_274),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_560),
.B(n_197),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_621),
.B(n_627),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_592),
.B(n_279),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_604),
.B(n_197),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_596),
.B(n_198),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_617),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_603),
.B(n_198),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_565),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_566),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_537),
.B(n_281),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_572),
.B(n_203),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_542),
.A2(n_196),
.B1(n_204),
.B2(n_341),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_538),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_548),
.B(n_203),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_538),
.B(n_204),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_613),
.B(n_209),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_613),
.B(n_209),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_567),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_583),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_581),
.B(n_212),
.Y(n_707)
);

NAND2x1p5_ASAP7_75t_L g708 ( 
.A(n_573),
.B(n_65),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_530),
.B(n_286),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_522),
.B(n_258),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_599),
.A2(n_210),
.B1(n_268),
.B2(n_305),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_504),
.B(n_292),
.C(n_289),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_516),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_L g714 ( 
.A1(n_547),
.A2(n_305),
.B1(n_210),
.B2(n_317),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_530),
.B(n_570),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_581),
.B(n_212),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_549),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_549),
.B(n_285),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_628),
.B(n_287),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_519),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_553),
.A2(n_304),
.B1(n_342),
.B2(n_339),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_573),
.A2(n_343),
.B(n_339),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_526),
.B(n_267),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_526),
.B(n_573),
.Y(n_724)
);

BUFx5_ASAP7_75t_L g725 ( 
.A(n_592),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_519),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_599),
.A2(n_578),
.B1(n_592),
.B2(n_561),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_523),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_533),
.B(n_293),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_583),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_590),
.B(n_267),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_523),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_525),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_600),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_600),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_629),
.B(n_626),
.Y(n_736)
);

A2O1A1Ixp33_ASAP7_75t_L g737 ( 
.A1(n_555),
.A2(n_334),
.B(n_270),
.C(n_307),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_534),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_553),
.Y(n_739)
);

CKINVDCx8_ASAP7_75t_R g740 ( 
.A(n_577),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_607),
.B(n_270),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_620),
.B(n_307),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_623),
.B(n_311),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_534),
.B(n_311),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_577),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_SL g746 ( 
.A1(n_522),
.A2(n_283),
.B1(n_288),
.B2(n_313),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_562),
.B(n_315),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_619),
.A2(n_318),
.B1(n_323),
.B2(n_294),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_533),
.B(n_522),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_591),
.A2(n_323),
.B1(n_318),
.B2(n_300),
.Y(n_750)
);

INVxp33_ASAP7_75t_L g751 ( 
.A(n_599),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_624),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_571),
.B(n_299),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_539),
.B(n_333),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_513),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_528),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_539),
.B(n_333),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_545),
.Y(n_758)
);

A2O1A1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_544),
.A2(n_330),
.B(n_329),
.C(n_321),
.Y(n_759)
);

AND2x6_ASAP7_75t_L g760 ( 
.A(n_550),
.B(n_313),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_539),
.B(n_330),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_675),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_715),
.B(n_550),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_637),
.B(n_556),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_675),
.Y(n_765)
);

AO22x1_ASAP7_75t_L g766 ( 
.A1(n_637),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

OAI21xp5_ASAP7_75t_L g768 ( 
.A1(n_630),
.A2(n_588),
.B(n_557),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_639),
.B(n_556),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_679),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_639),
.B(n_557),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_667),
.A2(n_610),
.B(n_321),
.C(n_329),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_672),
.B(n_558),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_672),
.B(n_584),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_611),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_674),
.A2(n_580),
.B(n_601),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_SL g777 ( 
.A1(n_656),
.A2(n_544),
.B(n_561),
.C(n_563),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_679),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_669),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_693),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_706),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_706),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_693),
.Y(n_783)
);

OA21x2_ASAP7_75t_L g784 ( 
.A1(n_697),
.A2(n_586),
.B(n_593),
.Y(n_784)
);

NAND2x1p5_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_671),
.Y(n_785)
);

OAI321xp33_ASAP7_75t_L g786 ( 
.A1(n_667),
.A2(n_589),
.A3(n_579),
.B1(n_574),
.B2(n_563),
.C(n_612),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_676),
.B(n_559),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_645),
.A2(n_622),
.B(n_574),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_653),
.B(n_533),
.Y(n_789)
);

O2A1O1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_700),
.A2(n_593),
.B(n_612),
.C(n_586),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_671),
.B(n_736),
.Y(n_791)
);

O2A1O1Ixp5_ASAP7_75t_L g792 ( 
.A1(n_645),
.A2(n_625),
.B(n_571),
.C(n_614),
.Y(n_792)
);

AOI21xp33_ASAP7_75t_L g793 ( 
.A1(n_707),
.A2(n_9),
.B(n_10),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_677),
.B(n_736),
.Y(n_794)
);

OAI22xp5_ASAP7_75t_L g795 ( 
.A1(n_638),
.A2(n_614),
.B1(n_571),
.B2(n_616),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_SL g796 ( 
.A(n_752),
.B(n_624),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_755),
.A2(n_622),
.B(n_616),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_665),
.B(n_615),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_716),
.B(n_644),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_717),
.A2(n_592),
.B1(n_551),
.B2(n_541),
.Y(n_800)
);

OAI21xp33_ASAP7_75t_L g801 ( 
.A1(n_666),
.A2(n_11),
.B(n_12),
.Y(n_801)
);

AOI21x1_ASAP7_75t_L g802 ( 
.A1(n_659),
.A2(n_541),
.B(n_585),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_684),
.B(n_551),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_689),
.B(n_551),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_655),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_706),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_651),
.B(n_551),
.Y(n_807)
);

O2A1O1Ixp5_ASAP7_75t_L g808 ( 
.A1(n_741),
.A2(n_568),
.B(n_71),
.C(n_72),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_725),
.B(n_568),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_633),
.B(n_13),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_737),
.A2(n_16),
.B(n_19),
.C(n_21),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_651),
.B(n_22),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_662),
.A2(n_751),
.B(n_731),
.C(n_657),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_SL g814 ( 
.A(n_636),
.B(n_22),
.C(n_23),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_676),
.A2(n_137),
.B1(n_136),
.B2(n_132),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_662),
.B(n_24),
.Y(n_816)
);

O2A1O1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_759),
.A2(n_28),
.B(n_31),
.C(n_33),
.Y(n_817)
);

O2A1O1Ixp5_ASAP7_75t_L g818 ( 
.A1(n_741),
.A2(n_127),
.B(n_126),
.C(n_122),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_695),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_753),
.A2(n_117),
.B(n_115),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_648),
.A2(n_36),
.B1(n_39),
.B2(n_44),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_725),
.B(n_101),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_SL g823 ( 
.A1(n_652),
.A2(n_36),
.B(n_39),
.C(n_44),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_SL g824 ( 
.A(n_740),
.B(n_86),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_702),
.B(n_45),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_SL g826 ( 
.A1(n_725),
.A2(n_80),
.B(n_48),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_681),
.A2(n_45),
.B(n_50),
.C(n_54),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_642),
.B(n_54),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_643),
.A2(n_56),
.B(n_57),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_756),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_673),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_709),
.A2(n_636),
.B1(n_719),
.B2(n_734),
.Y(n_832)
);

O2A1O1Ixp5_ASAP7_75t_L g833 ( 
.A1(n_742),
.A2(n_692),
.B(n_691),
.C(n_698),
.Y(n_833)
);

A2O1A1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_678),
.A2(n_699),
.B(n_711),
.C(n_712),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_649),
.B(n_650),
.Y(n_835)
);

NAND2xp33_ASAP7_75t_L g836 ( 
.A(n_725),
.B(n_706),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_701),
.B(n_694),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_696),
.B(n_705),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_678),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_735),
.A2(n_744),
.B(n_747),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_754),
.B(n_761),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_738),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_699),
.A2(n_710),
.B(n_711),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_739),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_754),
.B(n_761),
.Y(n_845)
);

OAI22xp33_ASAP7_75t_SL g846 ( 
.A1(n_743),
.A2(n_670),
.B1(n_658),
.B2(n_704),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_727),
.A2(n_757),
.B(n_718),
.C(n_682),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_680),
.A2(n_654),
.B(n_690),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_757),
.B(n_682),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_727),
.A2(n_686),
.B1(n_758),
.B2(n_713),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_730),
.B(n_726),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_680),
.A2(n_687),
.B(n_683),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_703),
.B(n_635),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_720),
.B(n_728),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_720),
.B(n_726),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_732),
.B(n_733),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_723),
.A2(n_722),
.B(n_641),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_688),
.A2(n_708),
.B(n_725),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_688),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_708),
.A2(n_739),
.B(n_729),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_714),
.B(n_749),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_760),
.A2(n_746),
.B1(n_721),
.B2(n_745),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_760),
.B(n_748),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_750),
.A2(n_739),
.B(n_663),
.C(n_760),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_646),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_760),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_685),
.B(n_646),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_685),
.A2(n_573),
.B(n_531),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_637),
.A2(n_667),
.B(n_716),
.C(n_707),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_736),
.A2(n_505),
.B1(n_637),
.B2(n_671),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_675),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_724),
.A2(n_573),
.B(n_531),
.Y(n_872)
);

AOI21x1_ASAP7_75t_L g873 ( 
.A1(n_660),
.A2(n_507),
.B(n_697),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_715),
.B(n_637),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_715),
.B(n_637),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_637),
.A2(n_507),
.B(n_715),
.C(n_700),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_630),
.A2(n_531),
.B(n_507),
.Y(n_877)
);

NOR2x1_ASAP7_75t_L g878 ( 
.A(n_632),
.B(n_543),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_637),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_647),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_634),
.A2(n_505),
.B1(n_640),
.B2(n_671),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_724),
.A2(n_573),
.B(n_531),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_715),
.B(n_637),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_630),
.A2(n_531),
.B(n_507),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_715),
.B(n_637),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_637),
.A2(n_707),
.B(n_716),
.C(n_736),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_630),
.A2(n_531),
.B(n_507),
.Y(n_887)
);

INVxp67_ASAP7_75t_SL g888 ( 
.A(n_638),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_668),
.A2(n_664),
.B(n_661),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_669),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_630),
.A2(n_531),
.B(n_507),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_671),
.B(n_634),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_646),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_631),
.B(n_637),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_637),
.A2(n_507),
.B(n_715),
.C(n_700),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_724),
.A2(n_573),
.B(n_531),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_634),
.A2(n_505),
.B1(n_640),
.B2(n_671),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_794),
.A2(n_894),
.B(n_869),
.Y(n_898)
);

OAI21xp5_ASAP7_75t_L g899 ( 
.A1(n_841),
.A2(n_845),
.B(n_877),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_844),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_874),
.B(n_875),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_870),
.A2(n_843),
.B(n_834),
.C(n_894),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_839),
.B(n_775),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_879),
.B(n_883),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_785),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_885),
.A2(n_791),
.B1(n_799),
.B2(n_897),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_872),
.A2(n_896),
.B(n_882),
.Y(n_907)
);

OAI22xp5_ASAP7_75t_L g908 ( 
.A1(n_791),
.A2(n_881),
.B1(n_847),
.B2(n_834),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_813),
.B(n_849),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_884),
.A2(n_891),
.B(n_887),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_762),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_830),
.Y(n_912)
);

AOI221x1_ASAP7_75t_L g913 ( 
.A1(n_813),
.A2(n_816),
.B1(n_847),
.B2(n_832),
.C(n_846),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_844),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_780),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_764),
.B(n_892),
.Y(n_916)
);

O2A1O1Ixp5_ASAP7_75t_L g917 ( 
.A1(n_857),
.A2(n_833),
.B(n_807),
.C(n_873),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_775),
.B(n_767),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_892),
.B(n_763),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_830),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_767),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_787),
.Y(n_922)
);

NOR2xp67_ASAP7_75t_L g923 ( 
.A(n_779),
.B(n_890),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_876),
.A2(n_895),
.B(n_792),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_773),
.B(n_774),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_871),
.Y(n_926)
);

AO31x2_ASAP7_75t_L g927 ( 
.A1(n_866),
.A2(n_840),
.A3(n_795),
.B(n_788),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_836),
.A2(n_858),
.B(n_776),
.Y(n_928)
);

O2A1O1Ixp5_ASAP7_75t_L g929 ( 
.A1(n_863),
.A2(n_771),
.B(n_769),
.C(n_848),
.Y(n_929)
);

INVx5_ASAP7_75t_L g930 ( 
.A(n_844),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_787),
.Y(n_931)
);

OAI21xp33_ASAP7_75t_L g932 ( 
.A1(n_801),
.A2(n_821),
.B(n_828),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_819),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_880),
.B(n_819),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_814),
.A2(n_793),
.B(n_772),
.C(n_827),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_861),
.B(n_837),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_812),
.B(n_838),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_781),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_785),
.A2(n_888),
.B1(n_861),
.B2(n_835),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_844),
.B(n_868),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_831),
.B(n_810),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_765),
.Y(n_942)
);

OAI21x1_ASAP7_75t_L g943 ( 
.A1(n_797),
.A2(n_809),
.B(n_855),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_777),
.A2(n_852),
.B(n_804),
.Y(n_944)
);

OAI21x1_ASAP7_75t_L g945 ( 
.A1(n_809),
.A2(n_854),
.B(n_856),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_777),
.A2(n_803),
.B(n_784),
.Y(n_946)
);

BUFx10_ASAP7_75t_L g947 ( 
.A(n_789),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_825),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_784),
.A2(n_790),
.B(n_822),
.Y(n_949)
);

AOI21xp33_ASAP7_75t_L g950 ( 
.A1(n_835),
.A2(n_853),
.B(n_828),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_770),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_859),
.B(n_878),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_860),
.A2(n_851),
.B(n_786),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_778),
.A2(n_783),
.B(n_798),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_850),
.A2(n_808),
.B(n_805),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_893),
.Y(n_956)
);

OAI22x1_ASAP7_75t_L g957 ( 
.A1(n_862),
.A2(n_853),
.B1(n_789),
.B2(n_810),
.Y(n_957)
);

OAI21xp5_ASAP7_75t_L g958 ( 
.A1(n_800),
.A2(n_818),
.B(n_772),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_842),
.A2(n_806),
.B(n_820),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_806),
.Y(n_960)
);

NAND2x1p5_ASAP7_75t_L g961 ( 
.A(n_781),
.B(n_782),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_798),
.B(n_821),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_826),
.Y(n_963)
);

AO31x2_ASAP7_75t_L g964 ( 
.A1(n_829),
.A2(n_864),
.A3(n_815),
.B(n_823),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_811),
.A2(n_817),
.B(n_823),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_766),
.B(n_796),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_865),
.B(n_824),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_867),
.A2(n_531),
.B(n_886),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_867),
.B(n_633),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_894),
.B(n_633),
.Y(n_970)
);

AND2x2_ASAP7_75t_SL g971 ( 
.A(n_821),
.B(n_710),
.Y(n_971)
);

INVx4_ASAP7_75t_L g972 ( 
.A(n_844),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_844),
.Y(n_973)
);

INVx6_ASAP7_75t_L g974 ( 
.A(n_844),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_762),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_872),
.A2(n_573),
.B(n_531),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_762),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_886),
.A2(n_869),
.B(n_794),
.C(n_834),
.Y(n_978)
);

OAI22xp5_ASAP7_75t_L g979 ( 
.A1(n_886),
.A2(n_870),
.B1(n_869),
.B2(n_794),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_794),
.B(n_874),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_886),
.A2(n_531),
.B(n_573),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_886),
.A2(n_870),
.B1(n_794),
.B2(n_637),
.Y(n_982)
);

AO21x1_ASAP7_75t_L g983 ( 
.A1(n_794),
.A2(n_845),
.B(n_841),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_886),
.A2(n_870),
.B1(n_869),
.B2(n_794),
.Y(n_984)
);

AOI21x1_ASAP7_75t_L g985 ( 
.A1(n_872),
.A2(n_896),
.B(n_882),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_794),
.B(n_874),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_794),
.B(n_874),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_886),
.A2(n_531),
.B(n_573),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_794),
.B(n_874),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_886),
.A2(n_870),
.B1(n_869),
.B2(n_794),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_830),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_794),
.B(n_874),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_765),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_794),
.B(n_874),
.Y(n_994)
);

AO31x2_ASAP7_75t_L g995 ( 
.A1(n_869),
.A2(n_847),
.A3(n_886),
.B(n_881),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_844),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_886),
.A2(n_531),
.B(n_573),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_859),
.B(n_844),
.Y(n_998)
);

BUFx12f_ASAP7_75t_L g999 ( 
.A(n_865),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_794),
.B(n_874),
.Y(n_1000)
);

INVx4_ASAP7_75t_L g1001 ( 
.A(n_844),
.Y(n_1001)
);

NAND3xp33_ASAP7_75t_L g1002 ( 
.A(n_886),
.B(n_637),
.C(n_869),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_830),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_889),
.A2(n_768),
.B(n_802),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_844),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_844),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_844),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_889),
.A2(n_768),
.B(n_802),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_794),
.A2(n_637),
.B(n_636),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_781),
.Y(n_1010)
);

AND2x4_ASAP7_75t_L g1011 ( 
.A(n_859),
.B(n_844),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_894),
.B(n_631),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_794),
.B(n_874),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_872),
.A2(n_573),
.B(n_531),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_794),
.B(n_874),
.Y(n_1015)
);

NAND3xp33_ASAP7_75t_L g1016 ( 
.A(n_886),
.B(n_637),
.C(n_869),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_SL g1017 ( 
.A1(n_886),
.A2(n_869),
.B(n_514),
.Y(n_1017)
);

AOI221xp5_ASAP7_75t_L g1018 ( 
.A1(n_869),
.A2(n_834),
.B1(n_793),
.B2(n_843),
.C(n_886),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_794),
.B(n_874),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_794),
.B(n_874),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_911),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_901),
.B(n_904),
.Y(n_1022)
);

AND2x6_ASAP7_75t_L g1023 ( 
.A(n_916),
.B(n_909),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_1009),
.A2(n_971),
.B1(n_932),
.B2(n_936),
.Y(n_1024)
);

AOI222xp33_ASAP7_75t_L g1025 ( 
.A1(n_898),
.A2(n_1018),
.B1(n_979),
.B2(n_984),
.C1(n_990),
.C2(n_1016),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_982),
.A2(n_1002),
.B1(n_1012),
.B2(n_970),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_1011),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_903),
.B(n_918),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_969),
.B(n_948),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_915),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_998),
.B(n_1011),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_938),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_981),
.A2(n_997),
.B(n_988),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_901),
.B(n_904),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_926),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1005),
.B(n_1006),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_L g1037 ( 
.A(n_923),
.B(n_972),
.Y(n_1037)
);

A2O1A1Ixp33_ASAP7_75t_SL g1038 ( 
.A1(n_924),
.A2(n_958),
.B(n_899),
.C(n_955),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_900),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_991),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_975),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_980),
.B(n_986),
.Y(n_1042)
);

AOI21xp33_ASAP7_75t_L g1043 ( 
.A1(n_978),
.A2(n_935),
.B(n_1018),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_977),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_SL g1045 ( 
.A(n_1003),
.B(n_934),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_980),
.B(n_986),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_987),
.B(n_989),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_922),
.B(n_931),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_900),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_902),
.B(n_913),
.C(n_992),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_987),
.B(n_989),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_933),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_992),
.B(n_994),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_994),
.B(n_1000),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_988),
.A2(n_997),
.B(n_953),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_1000),
.A2(n_1020),
.B(n_1019),
.C(n_1015),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_956),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_953),
.A2(n_976),
.B(n_1014),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_912),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_942),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_949),
.A2(n_925),
.B(n_944),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_993),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_949),
.A2(n_925),
.B(n_944),
.Y(n_1063)
);

AND2x6_ASAP7_75t_L g1064 ( 
.A(n_916),
.B(n_909),
.Y(n_1064)
);

AO21x2_ASAP7_75t_L g1065 ( 
.A1(n_907),
.A2(n_946),
.B(n_985),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_920),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_900),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_1013),
.A2(n_1020),
.B1(n_1019),
.B2(n_1015),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_921),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_938),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1013),
.A2(n_962),
.B1(n_937),
.B2(n_906),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_940),
.B(n_972),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_940),
.B(n_1001),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_919),
.B(n_962),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_908),
.A2(n_929),
.B(n_917),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_951),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_905),
.B(n_952),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_914),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_952),
.B(n_1001),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_941),
.B(n_939),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_968),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_SL g1082 ( 
.A(n_930),
.B(n_966),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_914),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_947),
.B(n_957),
.Y(n_1084)
);

OR2x2_ASAP7_75t_L g1085 ( 
.A(n_966),
.B(n_995),
.Y(n_1085)
);

HB1xp67_ASAP7_75t_L g1086 ( 
.A(n_930),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_947),
.B(n_983),
.Y(n_1087)
);

OR2x2_ASAP7_75t_L g1088 ( 
.A(n_995),
.B(n_960),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_930),
.B(n_973),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_965),
.A2(n_954),
.B(n_963),
.C(n_959),
.Y(n_1090)
);

CKINVDCx6p67_ASAP7_75t_R g1091 ( 
.A(n_914),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_973),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1010),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_973),
.Y(n_1094)
);

INVxp67_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_L g1096 ( 
.A(n_1010),
.B(n_940),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_996),
.B(n_1007),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_964),
.B(n_945),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_974),
.A2(n_1007),
.B1(n_961),
.B2(n_943),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_961),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_927),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_927),
.Y(n_1102)
);

NAND2x1p5_ASAP7_75t_L g1103 ( 
.A(n_1004),
.B(n_1008),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_903),
.B(n_631),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_911),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_970),
.B(n_936),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_933),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_901),
.B(n_904),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_970),
.B(n_936),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_970),
.B(n_936),
.Y(n_1110)
);

BUFx4_ASAP7_75t_SL g1111 ( 
.A(n_956),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_928),
.A2(n_886),
.B(n_1017),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_911),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_933),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_998),
.B(n_1011),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_933),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_911),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_970),
.B(n_936),
.Y(n_1118)
);

HB1xp67_ASAP7_75t_L g1119 ( 
.A(n_933),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_980),
.B(n_986),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_970),
.B(n_528),
.Y(n_1121)
);

BUFx8_ASAP7_75t_SL g1122 ( 
.A(n_999),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_999),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_940),
.B(n_844),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_950),
.B(n_775),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_900),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_933),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_928),
.A2(n_886),
.B(n_1017),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_900),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_970),
.B(n_936),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_900),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1009),
.A2(n_794),
.B(n_886),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_903),
.B(n_631),
.Y(n_1133)
);

INVx1_ASAP7_75t_SL g1134 ( 
.A(n_933),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_900),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_933),
.Y(n_1136)
);

BUFx5_ASAP7_75t_L g1137 ( 
.A(n_960),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_928),
.A2(n_886),
.B(n_1017),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_933),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_SL g1140 ( 
.A1(n_910),
.A2(n_886),
.B(n_869),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_928),
.A2(n_886),
.B(n_1017),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_933),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1009),
.A2(n_971),
.B1(n_870),
.B2(n_843),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_901),
.A2(n_886),
.B1(n_870),
.B2(n_869),
.Y(n_1144)
);

AND2x4_ASAP7_75t_L g1145 ( 
.A(n_998),
.B(n_1011),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_980),
.B(n_986),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1002),
.A2(n_886),
.B(n_1016),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_991),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_928),
.A2(n_886),
.B(n_1017),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_R g1150 ( 
.A(n_967),
.B(n_449),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_901),
.B(n_904),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_938),
.Y(n_1152)
);

CKINVDCx11_ASAP7_75t_R g1153 ( 
.A(n_1078),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1032),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_1135),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_1025),
.A2(n_1125),
.B1(n_1024),
.B2(n_1143),
.Y(n_1156)
);

BUFx12f_ASAP7_75t_L g1157 ( 
.A(n_1123),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1111),
.Y(n_1158)
);

INVx1_ASAP7_75t_SL g1159 ( 
.A(n_1029),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1025),
.A2(n_1024),
.B1(n_1143),
.B2(n_1043),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_1119),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_SL g1162 ( 
.A1(n_1150),
.A2(n_1144),
.B1(n_1133),
.B2(n_1104),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_1122),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_1081),
.B(n_1096),
.Y(n_1164)
);

OAI22xp33_ASAP7_75t_L g1165 ( 
.A1(n_1022),
.A2(n_1151),
.B1(n_1108),
.B2(n_1046),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_1057),
.Y(n_1166)
);

BUFx2_ASAP7_75t_L g1167 ( 
.A(n_1023),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1044),
.Y(n_1168)
);

NAND2x1p5_ASAP7_75t_L g1169 ( 
.A(n_1081),
.B(n_1088),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1034),
.A2(n_1047),
.B1(n_1054),
.B2(n_1120),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1171)
);

CKINVDCx14_ASAP7_75t_R g1172 ( 
.A(n_1048),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_1043),
.A2(n_1144),
.B1(n_1147),
.B2(n_1118),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1113),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1107),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1117),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1110),
.B(n_1130),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1077),
.B(n_1027),
.Y(n_1178)
);

CKINVDCx6p67_ASAP7_75t_R g1179 ( 
.A(n_1135),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1107),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1101),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1021),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1035),
.Y(n_1184)
);

AOI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1112),
.A2(n_1149),
.B(n_1128),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1026),
.B(n_1053),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1116),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1026),
.A2(n_1068),
.B1(n_1077),
.B2(n_1084),
.Y(n_1188)
);

BUFx6f_ASAP7_75t_L g1189 ( 
.A(n_1135),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1116),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1102),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1121),
.A2(n_1054),
.B1(n_1053),
.B2(n_1120),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1146),
.B(n_1042),
.Y(n_1193)
);

INVx3_ASAP7_75t_L g1194 ( 
.A(n_1032),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1052),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1114),
.Y(n_1196)
);

INVx4_ASAP7_75t_SL g1197 ( 
.A(n_1023),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_1023),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1027),
.B(n_1031),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_1127),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1134),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1041),
.Y(n_1202)
);

BUFx2_ASAP7_75t_R g1203 ( 
.A(n_1094),
.Y(n_1203)
);

BUFx2_ASAP7_75t_R g1204 ( 
.A(n_1136),
.Y(n_1204)
);

OAI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1051),
.A2(n_1146),
.B1(n_1082),
.B2(n_1068),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1105),
.Y(n_1206)
);

AO21x2_ASAP7_75t_L g1207 ( 
.A1(n_1058),
.A2(n_1033),
.B(n_1055),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1147),
.A2(n_1132),
.B1(n_1050),
.B2(n_1064),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1103),
.A2(n_1141),
.B(n_1138),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1134),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1076),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1082),
.A2(n_1050),
.B1(n_1028),
.B2(n_1071),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1132),
.A2(n_1023),
.B1(n_1064),
.B2(n_1071),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1060),
.Y(n_1214)
);

BUFx8_ASAP7_75t_L g1215 ( 
.A(n_1139),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1062),
.Y(n_1216)
);

AO21x2_ASAP7_75t_L g1217 ( 
.A1(n_1075),
.A2(n_1061),
.B(n_1063),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1080),
.A2(n_1045),
.B1(n_1074),
.B2(n_1087),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1093),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1074),
.B(n_1056),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1152),
.Y(n_1221)
);

BUFx4f_ASAP7_75t_SL g1222 ( 
.A(n_1091),
.Y(n_1222)
);

CKINVDCx8_ASAP7_75t_R g1223 ( 
.A(n_1142),
.Y(n_1223)
);

BUFx4_ASAP7_75t_R g1224 ( 
.A(n_1137),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1059),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1098),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1070),
.Y(n_1227)
);

AO21x2_ASAP7_75t_L g1228 ( 
.A1(n_1075),
.A2(n_1090),
.B(n_1038),
.Y(n_1228)
);

BUFx12f_ASAP7_75t_L g1229 ( 
.A(n_1036),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1031),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1152),
.Y(n_1231)
);

BUFx4f_ASAP7_75t_SL g1232 ( 
.A(n_1036),
.Y(n_1232)
);

BUFx8_ASAP7_75t_L g1233 ( 
.A(n_1083),
.Y(n_1233)
);

AO21x2_ASAP7_75t_L g1234 ( 
.A1(n_1140),
.A2(n_1098),
.B(n_1065),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_1066),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1064),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1115),
.B(n_1145),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1097),
.Y(n_1238)
);

INVxp33_ASAP7_75t_L g1239 ( 
.A(n_1069),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1099),
.B(n_1100),
.Y(n_1240)
);

BUFx12f_ASAP7_75t_L g1241 ( 
.A(n_1040),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1148),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1145),
.B(n_1124),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1095),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1124),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_1039),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1079),
.A2(n_1073),
.B1(n_1072),
.B2(n_1037),
.Y(n_1247)
);

AO21x1_ASAP7_75t_SL g1248 ( 
.A1(n_1099),
.A2(n_1086),
.B(n_1072),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1089),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1072),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_1073),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1039),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1049),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1067),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1097),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1092),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1092),
.B(n_1131),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1126),
.A2(n_971),
.B1(n_1009),
.B2(n_932),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1126),
.A2(n_971),
.B1(n_1009),
.B2(n_932),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1126),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1129),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1129),
.A2(n_971),
.B1(n_1009),
.B2(n_932),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1129),
.Y(n_1263)
);

BUFx8_ASAP7_75t_L g1264 ( 
.A(n_1052),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1030),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1106),
.B(n_1109),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1150),
.A2(n_971),
.B1(n_710),
.B2(n_936),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1034),
.A2(n_886),
.B1(n_870),
.B2(n_1151),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1171),
.B(n_1177),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1191),
.Y(n_1270)
);

BUFx2_ASAP7_75t_L g1271 ( 
.A(n_1169),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1226),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1175),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1186),
.B(n_1180),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1169),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1181),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1162),
.B(n_1267),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1186),
.B(n_1180),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1236),
.Y(n_1279)
);

HB1xp67_ASAP7_75t_L g1280 ( 
.A(n_1187),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1201),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1210),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1248),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1167),
.B(n_1198),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1182),
.Y(n_1285)
);

OR2x6_ASAP7_75t_L g1286 ( 
.A(n_1185),
.B(n_1209),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1193),
.B(n_1170),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1250),
.B(n_1251),
.Y(n_1288)
);

BUFx4f_ASAP7_75t_L g1289 ( 
.A(n_1155),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1218),
.B(n_1208),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1161),
.Y(n_1291)
);

INVxp67_ASAP7_75t_R g1292 ( 
.A(n_1192),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1183),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1165),
.B(n_1177),
.Y(n_1294)
);

OR2x6_ASAP7_75t_L g1295 ( 
.A(n_1167),
.B(n_1198),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1184),
.Y(n_1296)
);

INVx3_ASAP7_75t_SL g1297 ( 
.A(n_1179),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1188),
.B(n_1234),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1220),
.Y(n_1299)
);

HB1xp67_ASAP7_75t_L g1300 ( 
.A(n_1190),
.Y(n_1300)
);

BUFx4f_ASAP7_75t_L g1301 ( 
.A(n_1155),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1240),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_SL g1303 ( 
.A1(n_1268),
.A2(n_1164),
.B(n_1189),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1240),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1173),
.B(n_1266),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1217),
.A2(n_1207),
.B(n_1205),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1266),
.B(n_1159),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1240),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1248),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1158),
.Y(n_1310)
);

BUFx2_ASAP7_75t_L g1311 ( 
.A(n_1164),
.Y(n_1311)
);

OR2x2_ASAP7_75t_L g1312 ( 
.A(n_1234),
.B(n_1213),
.Y(n_1312)
);

OAI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1160),
.A2(n_1156),
.B(n_1259),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_1224),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1202),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1206),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1163),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1195),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1234),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1228),
.B(n_1212),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_SL g1322 ( 
.A(n_1158),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1228),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1197),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1217),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1197),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1243),
.B(n_1219),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1217),
.A2(n_1249),
.B(n_1221),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_L g1329 ( 
.A(n_1195),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1197),
.Y(n_1330)
);

AND2x4_ASAP7_75t_L g1331 ( 
.A(n_1245),
.B(n_1243),
.Y(n_1331)
);

BUFx3_ASAP7_75t_R g1332 ( 
.A(n_1204),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1168),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_1235),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1258),
.A2(n_1262),
.B(n_1211),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1239),
.A2(n_1247),
.B(n_1242),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1174),
.B(n_1265),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1270),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1313),
.A2(n_1178),
.B1(n_1172),
.B2(n_1199),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1323),
.B(n_1176),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_1314),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1273),
.Y(n_1342)
);

AOI33xp33_ASAP7_75t_L g1343 ( 
.A1(n_1320),
.A2(n_1214),
.A3(n_1216),
.B1(n_1255),
.B2(n_1263),
.B3(n_1253),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1274),
.B(n_1231),
.Y(n_1344)
);

OA21x2_ASAP7_75t_L g1345 ( 
.A1(n_1306),
.A2(n_1252),
.B(n_1254),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1278),
.B(n_1231),
.Y(n_1346)
);

NAND2x1_ASAP7_75t_L g1347 ( 
.A(n_1303),
.B(n_1231),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1278),
.B(n_1227),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1287),
.B(n_1200),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1320),
.B(n_1227),
.Y(n_1350)
);

NOR4xp25_ASAP7_75t_SL g1351 ( 
.A(n_1277),
.B(n_1246),
.C(n_1235),
.D(n_1225),
.Y(n_1351)
);

INVx11_ASAP7_75t_L g1352 ( 
.A(n_1332),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1295),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1285),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1290),
.A2(n_1225),
.B1(n_1196),
.B2(n_1244),
.C(n_1178),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1312),
.B(n_1154),
.Y(n_1356)
);

INVx5_ASAP7_75t_L g1357 ( 
.A(n_1286),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1312),
.B(n_1194),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1276),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1290),
.A2(n_1178),
.B(n_1199),
.C(n_1155),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1325),
.B(n_1257),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1272),
.B(n_1257),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1303),
.B(n_1189),
.Y(n_1363)
);

AOI221xp5_ASAP7_75t_L g1364 ( 
.A1(n_1294),
.A2(n_1196),
.B1(n_1244),
.B2(n_1199),
.C(n_1237),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1295),
.Y(n_1365)
);

OR2x2_ASAP7_75t_L g1366 ( 
.A(n_1298),
.B(n_1256),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1305),
.A2(n_1237),
.B1(n_1230),
.B2(n_1264),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1328),
.Y(n_1368)
);

INVxp67_ASAP7_75t_L g1369 ( 
.A(n_1299),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1328),
.Y(n_1370)
);

OAI31xp33_ASAP7_75t_L g1371 ( 
.A1(n_1300),
.A2(n_1238),
.A3(n_1260),
.B(n_1261),
.Y(n_1371)
);

AOI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1292),
.A2(n_1230),
.B1(n_1166),
.B2(n_1229),
.Y(n_1372)
);

NAND2x1_ASAP7_75t_L g1373 ( 
.A(n_1314),
.B(n_1302),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1299),
.B(n_1223),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1338),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1364),
.A2(n_1314),
.B1(n_1305),
.B2(n_1331),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1342),
.B(n_1280),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1355),
.B(n_1336),
.C(n_1282),
.Y(n_1378)
);

NOR3xp33_ASAP7_75t_SL g1379 ( 
.A(n_1374),
.B(n_1310),
.C(n_1246),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1342),
.B(n_1281),
.Y(n_1380)
);

NAND3xp33_ASAP7_75t_L g1381 ( 
.A(n_1355),
.B(n_1343),
.C(n_1364),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1372),
.B(n_1283),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1339),
.A2(n_1292),
.B1(n_1334),
.B2(n_1223),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1359),
.B(n_1291),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1350),
.B(n_1271),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1361),
.B(n_1275),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1343),
.B(n_1269),
.C(n_1335),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1341),
.A2(n_1309),
.B1(n_1283),
.B2(n_1321),
.Y(n_1388)
);

NAND3xp33_ASAP7_75t_L g1389 ( 
.A(n_1371),
.B(n_1304),
.C(n_1308),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1361),
.B(n_1275),
.Y(n_1390)
);

AOI221x1_ASAP7_75t_SL g1391 ( 
.A1(n_1349),
.A2(n_1307),
.B1(n_1332),
.B2(n_1316),
.C(n_1333),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1339),
.A2(n_1297),
.B1(n_1326),
.B2(n_1309),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1349),
.B(n_1315),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1361),
.B(n_1295),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1338),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1367),
.A2(n_1331),
.B1(n_1309),
.B2(n_1283),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1356),
.B(n_1358),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1356),
.B(n_1284),
.Y(n_1398)
);

OAI21xp33_ASAP7_75t_L g1399 ( 
.A1(n_1372),
.A2(n_1327),
.B(n_1337),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1356),
.B(n_1284),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1352),
.A2(n_1297),
.B1(n_1326),
.B2(n_1283),
.Y(n_1401)
);

OA211x2_ASAP7_75t_L g1402 ( 
.A1(n_1371),
.A2(n_1347),
.B(n_1373),
.C(n_1374),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1362),
.B(n_1288),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1363),
.B(n_1283),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1297),
.B1(n_1309),
.B2(n_1283),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1352),
.A2(n_1309),
.B1(n_1289),
.B2(n_1301),
.Y(n_1406)
);

NAND3xp33_ASAP7_75t_L g1407 ( 
.A(n_1367),
.B(n_1351),
.C(n_1369),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1362),
.B(n_1288),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1362),
.B(n_1288),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1358),
.B(n_1279),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1358),
.B(n_1279),
.Y(n_1411)
);

NAND3xp33_ASAP7_75t_L g1412 ( 
.A(n_1351),
.B(n_1311),
.C(n_1335),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1360),
.A2(n_1309),
.B1(n_1289),
.B2(n_1301),
.Y(n_1413)
);

OAI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1360),
.A2(n_1301),
.B1(n_1289),
.B2(n_1318),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1366),
.B(n_1319),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1363),
.A2(n_1286),
.B(n_1302),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1341),
.A2(n_1329),
.B1(n_1324),
.B2(n_1330),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1348),
.B(n_1293),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1348),
.B(n_1296),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1348),
.B(n_1296),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1375),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1375),
.Y(n_1423)
);

NAND2x1_ASAP7_75t_L g1424 ( 
.A(n_1416),
.B(n_1353),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1395),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1395),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1397),
.B(n_1345),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1415),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1415),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1393),
.B(n_1369),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1397),
.B(n_1345),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1394),
.B(n_1345),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1394),
.B(n_1345),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1398),
.B(n_1345),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1384),
.B(n_1322),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1404),
.B(n_1357),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1377),
.B(n_1317),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1410),
.Y(n_1438)
);

BUFx2_ASAP7_75t_L g1439 ( 
.A(n_1411),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1419),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1420),
.B(n_1368),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1421),
.B(n_1368),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1400),
.B(n_1386),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1380),
.B(n_1340),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1417),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1390),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1378),
.B(n_1215),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1403),
.B(n_1370),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1408),
.B(n_1370),
.Y(n_1449)
);

NAND2x1_ASAP7_75t_L g1450 ( 
.A(n_1387),
.B(n_1353),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1427),
.B(n_1385),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1427),
.B(n_1385),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1440),
.B(n_1391),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1422),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1441),
.B(n_1409),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1422),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1427),
.B(n_1357),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1423),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1423),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1441),
.B(n_1387),
.Y(n_1460)
);

NOR2x1_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_1407),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1441),
.B(n_1366),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1431),
.B(n_1357),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1423),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1447),
.B(n_1157),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1436),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1431),
.B(n_1434),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1436),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_SL g1469 ( 
.A1(n_1435),
.A2(n_1381),
.B1(n_1378),
.B2(n_1383),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1431),
.B(n_1357),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1425),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1366),
.Y(n_1472)
);

AND3x2_ASAP7_75t_L g1473 ( 
.A(n_1437),
.B(n_1402),
.C(n_1311),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1430),
.B(n_1381),
.Y(n_1474)
);

OAI221xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1450),
.A2(n_1399),
.B1(n_1376),
.B2(n_1396),
.C(n_1412),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1425),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1434),
.B(n_1357),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1425),
.Y(n_1478)
);

AND2x4_ASAP7_75t_SL g1479 ( 
.A(n_1438),
.B(n_1341),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1426),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1432),
.B(n_1357),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1426),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1436),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1440),
.B(n_1354),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1434),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1429),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1432),
.B(n_1357),
.Y(n_1487)
);

NAND2x1_ASAP7_75t_L g1488 ( 
.A(n_1432),
.B(n_1365),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1445),
.B(n_1354),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1460),
.B(n_1448),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1480),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1451),
.B(n_1433),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1454),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1451),
.B(n_1433),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1451),
.B(n_1452),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1480),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1474),
.B(n_1445),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1480),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1482),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1454),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1482),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1486),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1504)
);

AOI22xp5_ASAP7_75t_L g1505 ( 
.A1(n_1469),
.A2(n_1402),
.B1(n_1382),
.B2(n_1450),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1486),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1456),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1489),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1474),
.B(n_1430),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1456),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1453),
.B(n_1429),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1452),
.B(n_1439),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1439),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1453),
.B(n_1444),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1464),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1516)
);

BUFx2_ASAP7_75t_L g1517 ( 
.A(n_1461),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1464),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1460),
.B(n_1448),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1454),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1484),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1484),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1460),
.B(n_1448),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1462),
.B(n_1449),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1469),
.B(n_1444),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1489),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1461),
.B(n_1428),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1529)
);

INVx6_ASAP7_75t_L g1530 ( 
.A(n_1468),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1462),
.B(n_1449),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1466),
.B(n_1446),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1458),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1473),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1511),
.B(n_1490),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1528),
.A2(n_1488),
.B(n_1424),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1512),
.B(n_1483),
.Y(n_1539)
);

NOR2x1_ASAP7_75t_L g1540 ( 
.A(n_1517),
.B(n_1497),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1506),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1490),
.B(n_1455),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1530),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1503),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1514),
.B(n_1473),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1519),
.B(n_1455),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1524),
.B(n_1462),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1495),
.B(n_1468),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1503),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1491),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1524),
.B(n_1472),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1443),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_L g1554 ( 
.A(n_1517),
.B(n_1465),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1491),
.Y(n_1555)
);

NAND2x1p5_ASAP7_75t_L g1556 ( 
.A(n_1505),
.B(n_1468),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1496),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1513),
.B(n_1487),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1505),
.B(n_1508),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1496),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1507),
.B(n_1475),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1498),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1493),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1498),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1525),
.B(n_1472),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1522),
.B(n_1523),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1530),
.A2(n_1392),
.B1(n_1399),
.B2(n_1414),
.Y(n_1568)
);

AO21x2_ASAP7_75t_L g1569 ( 
.A1(n_1507),
.A2(n_1471),
.B(n_1458),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1537),
.B(n_1516),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1562),
.B(n_1541),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1544),
.Y(n_1572)
);

XNOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1556),
.B(n_1401),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1562),
.A2(n_1530),
.B1(n_1405),
.B2(n_1521),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1553),
.B(n_1522),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1554),
.B(n_1436),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1550),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1551),
.Y(n_1578)
);

OAI221xp5_ASAP7_75t_L g1579 ( 
.A1(n_1556),
.A2(n_1475),
.B1(n_1530),
.B2(n_1523),
.C(n_1527),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1543),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1535),
.B(n_1525),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1540),
.B(n_1515),
.C(n_1510),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1535),
.B(n_1527),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1555),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1543),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1537),
.B(n_1531),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1568),
.B(n_1516),
.Y(n_1587)
);

NAND4xp25_ASAP7_75t_SL g1588 ( 
.A(n_1560),
.B(n_1163),
.C(n_1487),
.D(n_1529),
.Y(n_1588)
);

A2O1A1Ixp33_ASAP7_75t_L g1589 ( 
.A1(n_1546),
.A2(n_1379),
.B(n_1488),
.C(n_1529),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1567),
.B(n_1510),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1558),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1534),
.B(n_1531),
.Y(n_1592)
);

INVxp33_ASAP7_75t_L g1593 ( 
.A(n_1536),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_SL g1594 ( 
.A1(n_1543),
.A2(n_1166),
.B1(n_1157),
.B2(n_1515),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1561),
.Y(n_1595)
);

NAND2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1580),
.B(n_1538),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1571),
.B(n_1536),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1571),
.B(n_1539),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1543),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1585),
.B(n_1539),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1593),
.B(n_1549),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1549),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1587),
.B(n_1557),
.Y(n_1603)
);

AOI222xp33_ASAP7_75t_L g1604 ( 
.A1(n_1579),
.A2(n_1518),
.B1(n_1557),
.B2(n_1559),
.C1(n_1532),
.C2(n_1538),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1574),
.B(n_1542),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1578),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1570),
.B(n_1559),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1573),
.A2(n_1542),
.B1(n_1547),
.B2(n_1545),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1584),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1570),
.B(n_1545),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1572),
.B(n_1577),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1591),
.B(n_1547),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1595),
.B(n_1548),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1581),
.B(n_1548),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1586),
.Y(n_1615)
);

AOI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1599),
.A2(n_1594),
.B1(n_1582),
.B2(n_1589),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_R g1617 ( 
.A(n_1597),
.B(n_1153),
.Y(n_1617)
);

XOR2x2_ASAP7_75t_L g1618 ( 
.A(n_1605),
.B(n_1576),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1615),
.B(n_1575),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1604),
.A2(n_1590),
.B(n_1575),
.C(n_1583),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1608),
.A2(n_1590),
.B(n_1583),
.Y(n_1621)
);

O2A1O1Ixp33_ASAP7_75t_L g1622 ( 
.A1(n_1598),
.A2(n_1518),
.B(n_1565),
.C(n_1563),
.Y(n_1622)
);

NAND4xp75_ASAP7_75t_L g1623 ( 
.A(n_1603),
.B(n_1564),
.C(n_1532),
.D(n_1521),
.Y(n_1623)
);

AOI222xp33_ASAP7_75t_L g1624 ( 
.A1(n_1602),
.A2(n_1564),
.B1(n_1492),
.B2(n_1494),
.C1(n_1504),
.C2(n_1499),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1611),
.A2(n_1552),
.B(n_1569),
.C(n_1566),
.Y(n_1625)
);

AOI221xp5_ASAP7_75t_L g1626 ( 
.A1(n_1601),
.A2(n_1552),
.B1(n_1566),
.B2(n_1569),
.C(n_1533),
.Y(n_1626)
);

AOI222xp33_ASAP7_75t_L g1627 ( 
.A1(n_1612),
.A2(n_1613),
.B1(n_1609),
.B2(n_1606),
.C1(n_1614),
.C2(n_1610),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1616),
.A2(n_1600),
.B1(n_1607),
.B2(n_1596),
.Y(n_1628)
);

NAND3xp33_ASAP7_75t_L g1629 ( 
.A(n_1625),
.B(n_1264),
.C(n_1215),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1619),
.B(n_1596),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1621),
.B(n_1492),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1620),
.A2(n_1481),
.B1(n_1500),
.B2(n_1499),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1617),
.Y(n_1633)
);

NAND2x1_ASAP7_75t_SL g1634 ( 
.A(n_1618),
.B(n_1494),
.Y(n_1634)
);

NAND4xp75_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1533),
.C(n_1457),
.D(n_1470),
.Y(n_1635)
);

NOR2xp67_ASAP7_75t_L g1636 ( 
.A(n_1623),
.B(n_1500),
.Y(n_1636)
);

NAND3xp33_ASAP7_75t_L g1637 ( 
.A(n_1627),
.B(n_1264),
.C(n_1215),
.Y(n_1637)
);

NOR2x1_ASAP7_75t_L g1638 ( 
.A(n_1622),
.B(n_1569),
.Y(n_1638)
);

NAND4xp75_ASAP7_75t_L g1639 ( 
.A(n_1624),
.B(n_1470),
.C(n_1463),
.D(n_1457),
.Y(n_1639)
);

NAND4xp25_ASAP7_75t_SL g1640 ( 
.A(n_1637),
.B(n_1504),
.C(n_1457),
.D(n_1463),
.Y(n_1640)
);

NAND4xp25_ASAP7_75t_SL g1641 ( 
.A(n_1638),
.B(n_1463),
.C(n_1470),
.D(n_1477),
.Y(n_1641)
);

NAND4xp75_ASAP7_75t_L g1642 ( 
.A(n_1630),
.B(n_1153),
.C(n_1502),
.D(n_1477),
.Y(n_1642)
);

NOR2x1_ASAP7_75t_L g1643 ( 
.A(n_1628),
.B(n_1502),
.Y(n_1643)
);

NAND4xp25_ASAP7_75t_L g1644 ( 
.A(n_1633),
.B(n_1406),
.C(n_1388),
.D(n_1481),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1629),
.A2(n_1520),
.B(n_1493),
.C(n_1501),
.Y(n_1645)
);

NAND4xp25_ASAP7_75t_L g1646 ( 
.A(n_1631),
.B(n_1636),
.C(n_1632),
.D(n_1634),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1643),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1646),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1642),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1644),
.B(n_1640),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1641),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1645),
.Y(n_1652)
);

AOI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1640),
.A2(n_1639),
.B1(n_1635),
.B2(n_1481),
.Y(n_1653)
);

OAI321xp33_ASAP7_75t_L g1654 ( 
.A1(n_1648),
.A2(n_1520),
.A3(n_1501),
.B1(n_1413),
.B2(n_1477),
.C(n_1418),
.Y(n_1654)
);

AOI32xp33_ASAP7_75t_L g1655 ( 
.A1(n_1651),
.A2(n_1481),
.A3(n_1467),
.B1(n_1485),
.B2(n_1446),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1647),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1649),
.B(n_1222),
.C(n_1241),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1652),
.B(n_1467),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1650),
.B(n_1241),
.C(n_1389),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1658),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1656),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1655),
.Y(n_1662)
);

XNOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1662),
.B(n_1657),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1663),
.A2(n_1660),
.B(n_1661),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1660),
.B1(n_1659),
.B2(n_1653),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_1664),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1666),
.Y(n_1667)
);

XOR2xp5_ASAP7_75t_L g1668 ( 
.A(n_1665),
.B(n_1203),
.Y(n_1668)
);

AOI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1668),
.A2(n_1654),
.B1(n_1481),
.B2(n_1485),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1667),
.A2(n_1485),
.B(n_1471),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1669),
.A2(n_1179),
.B1(n_1467),
.B2(n_1232),
.Y(n_1671)
);

AOI322xp5_ASAP7_75t_L g1672 ( 
.A1(n_1671),
.A2(n_1670),
.A3(n_1458),
.B1(n_1471),
.B2(n_1476),
.C1(n_1459),
.C2(n_1478),
.Y(n_1672)
);

OAI221xp5_ASAP7_75t_R g1673 ( 
.A1(n_1672),
.A2(n_1233),
.B1(n_1229),
.B2(n_1476),
.C(n_1478),
.Y(n_1673)
);

AOI211xp5_ASAP7_75t_L g1674 ( 
.A1(n_1673),
.A2(n_1155),
.B(n_1189),
.C(n_1260),
.Y(n_1674)
);


endmodule