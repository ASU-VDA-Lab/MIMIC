module fake_jpeg_3220_n_153 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_153);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_153;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_58),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_52),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_57),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_64),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_51),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_45),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_69),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_50),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_1),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_55),
.B1(n_57),
.B2(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_57),
.B1(n_38),
.B2(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_66),
.B1(n_43),
.B2(n_38),
.Y(n_75)
);

OAI22x1_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_56),
.B1(n_48),
.B2(n_44),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_4),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_56),
.B1(n_48),
.B2(n_44),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_46),
.B1(n_40),
.B2(n_41),
.Y(n_87)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_48),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_61),
.B1(n_52),
.B2(n_49),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_41),
.B1(n_19),
.B2(n_21),
.Y(n_97)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_97),
.B1(n_91),
.B2(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_90),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_78),
.B(n_2),
.Y(n_90)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_81),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_91),
.A2(n_23),
.B(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_94),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_4),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_16),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_20),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_9),
.Y(n_112)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_112),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_76),
.B1(n_7),
.B2(n_8),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_108),
.B1(n_109),
.B2(n_10),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_6),
.B(n_8),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_11),
.B(n_14),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_9),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_26),
.B(n_27),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_17),
.B1(n_32),
.B2(n_30),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_126)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_14),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_93),
.B1(n_92),
.B2(n_12),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_116),
.A2(n_126),
.B1(n_110),
.B2(n_115),
.Y(n_134)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_104),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_24),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_107),
.C(n_112),
.Y(n_131)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_37),
.B(n_29),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_128),
.B(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_105),
.C(n_15),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_122),
.C(n_115),
.Y(n_142)
);

XNOR2x2_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_117),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_124),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_143),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_130),
.C(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_141),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_145),
.A2(n_139),
.B1(n_140),
.B2(n_124),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_126),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_146),
.C(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_118),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_150),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_151),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_15),
.Y(n_153)
);


endmodule