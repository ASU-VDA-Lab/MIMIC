module fake_jpeg_5409_n_160 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_160);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_2),
.B(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_25),
.Y(n_30)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_23),
.A2(n_11),
.B1(n_21),
.B2(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_26),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_11),
.B1(n_21),
.B2(n_14),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_38),
.B1(n_26),
.B2(n_28),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_27),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_23),
.A2(n_11),
.B1(n_21),
.B2(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_44),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_24),
.B(n_26),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_47),
.B1(n_36),
.B2(n_23),
.Y(n_55)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_26),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_29),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_45),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_51),
.B1(n_47),
.B2(n_42),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_23),
.B1(n_22),
.B2(n_25),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_25),
.B1(n_32),
.B2(n_33),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_47),
.A2(n_28),
.B1(n_32),
.B2(n_36),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_43),
.B(n_44),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_39),
.A2(n_32),
.B1(n_36),
.B2(n_35),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_75),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_77),
.B(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_63),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_70),
.B(n_71),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_65),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_52),
.B(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_45),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_58),
.B(n_54),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_45),
.B(n_49),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_61),
.B(n_15),
.Y(n_100)
);

NAND2xp67_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_58),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_82),
.B(n_76),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_57),
.C(n_56),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_75),
.C(n_73),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_84),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_72),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_64),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_28),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_68),
.B1(n_73),
.B2(n_59),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_91),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_53),
.B1(n_74),
.B2(n_73),
.Y(n_94)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_97),
.C(n_81),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_57),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_82),
.A2(n_61),
.B1(n_40),
.B2(n_12),
.Y(n_98)
);

AO32x1_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_79),
.A3(n_87),
.B1(n_89),
.B2(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_99),
.B(n_101),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_85),
.A2(n_13),
.B1(n_16),
.B2(n_20),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_103),
.A2(n_18),
.B(n_19),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_113),
.C(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_89),
.C(n_29),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_111),
.C(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_18),
.Y(n_109)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_109),
.Y(n_125)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_110),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_28),
.C(n_15),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_18),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_8),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g115 ( 
.A(n_95),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_90),
.C(n_94),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_122),
.C(n_106),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_91),
.C(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_91),
.B1(n_102),
.B2(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_102),
.B1(n_20),
.B2(n_16),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_127),
.Y(n_136)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_116),
.A2(n_20),
.B1(n_16),
.B2(n_13),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_130),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_113),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_0),
.C(n_1),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_116),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_134),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_110),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_9),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_133),
.A3(n_135),
.B1(n_136),
.B2(n_132),
.C1(n_134),
.C2(n_128),
.Y(n_139)
);

AOI211xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_142),
.B(n_7),
.C(n_2),
.Y(n_146)
);

AOI322xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_117),
.A3(n_125),
.B1(n_126),
.B2(n_120),
.C1(n_19),
.C2(n_28),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_144),
.B(n_6),
.Y(n_149)
);

OAI31xp33_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_8),
.A3(n_7),
.B(n_3),
.Y(n_145)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_146),
.B(n_6),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_0),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_0),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_148),
.A2(n_149),
.B(n_4),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_4),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_155),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_5),
.B1(n_6),
.B2(n_154),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_5),
.B1(n_157),
.B2(n_156),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_156),
.Y(n_160)
);


endmodule