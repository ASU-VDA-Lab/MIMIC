module fake_jpeg_18526_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx12_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_5),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g110 ( 
.A(n_86),
.Y(n_110)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_90),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_79),
.B(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_73),
.Y(n_91)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_60),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_72),
.Y(n_122)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_117),
.Y(n_125)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_93),
.A2(n_55),
.B(n_49),
.Y(n_107)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_115),
.CI(n_67),
.CON(n_126),
.SN(n_126)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_113),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_95),
.A2(n_62),
.B1(n_50),
.B2(n_66),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_112),
.B1(n_116),
.B2(n_121),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_58),
.B1(n_65),
.B2(n_68),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_69),
.C(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_59),
.B1(n_49),
.B2(n_55),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_122),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_83),
.A2(n_55),
.B1(n_63),
.B2(n_56),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_105),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_126),
.Y(n_139)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_127),
.A2(n_110),
.B1(n_99),
.B2(n_111),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_105),
.B(n_57),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_134),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_107),
.A2(n_57),
.B1(n_72),
.B2(n_23),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_130),
.A2(n_128),
.B1(n_125),
.B2(n_126),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_128),
.B1(n_133),
.B2(n_132),
.Y(n_147)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_142),
.Y(n_145)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_135),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_144),
.A2(n_139),
.B1(n_100),
.B2(n_137),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_145),
.B1(n_139),
.B2(n_146),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_150),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_151),
.B(n_153),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_101),
.B1(n_102),
.B2(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_19),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_24),
.Y(n_154)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_145),
.B(n_106),
.C(n_17),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_155),
.B1(n_25),
.B2(n_28),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_160),
.A2(n_161),
.B1(n_155),
.B2(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_158),
.B(n_159),
.Y(n_161)
);

OAI322xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_14),
.A3(n_47),
.B1(n_46),
.B2(n_40),
.C1(n_39),
.C2(n_38),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_6),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_7),
.C(n_37),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_48),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_34),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_33),
.C(n_32),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_168),
.A2(n_31),
.B(n_30),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_15),
.C(n_9),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_171),
.Y(n_172)
);

AOI31xp33_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_0),
.A3(n_1),
.B(n_2),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_173),
.Y(n_174)
);


endmodule