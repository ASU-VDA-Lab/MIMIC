module fake_netlist_5_2398_n_2628 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_547, n_43, n_116, n_22, n_467, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_382, n_254, n_33, n_23, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_106, n_209, n_259, n_448, n_375, n_301, n_68, n_93, n_186, n_537, n_134, n_191, n_51, n_63, n_492, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_221, n_178, n_386, n_287, n_344, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_384, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_504, n_511, n_12, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_340, n_207, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_113, n_246, n_179, n_125, n_410, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_426, n_520, n_409, n_500, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2628);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_382;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_51;
input n_63;
input n_492;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_221;
input n_178;
input n_386;
input n_287;
input n_344;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_384;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_504;
input n_511;
input n_12;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_426;
input n_520;
input n_409;
input n_500;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2628;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2031;
wire n_556;
wire n_2076;
wire n_2482;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_731;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2300;
wire n_1796;
wire n_2551;
wire n_1473;
wire n_680;
wire n_1587;
wire n_553;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_888;
wire n_1880;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_571;
wire n_1585;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_1053;
wire n_1224;
wire n_2557;
wire n_1926;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2616;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2331;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_1415;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_2577;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_2342;
wire n_633;
wire n_1832;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_1964;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_724;
wire n_2084;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_2168;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_1574;
wire n_2399;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2418;
wire n_829;
wire n_2519;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_2467;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2541;
wire n_1139;
wire n_2333;
wire n_885;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_2475;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2556;
wire n_2269;
wire n_2309;
wire n_2415;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2287;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2325;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2034;
wire n_1637;
wire n_1687;
wire n_1419;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_770;
wire n_1375;
wire n_2494;
wire n_1102;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_1399;
wire n_1543;
wire n_2224;
wire n_1991;
wire n_791;
wire n_732;
wire n_1533;
wire n_1979;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_1067;
wire n_1720;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2332;
wire n_1235;
wire n_980;
wire n_698;
wire n_1115;
wire n_703;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2497;
wire n_2006;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2456;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_1287;
wire n_1262;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2525;
wire n_2513;
wire n_1764;
wire n_712;
wire n_2414;
wire n_1583;
wire n_2426;
wire n_1042;
wire n_1402;
wire n_2049;
wire n_2273;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_2044;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_2599;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_1542;
wire n_1251;
wire n_2268;

INVx1_ASAP7_75t_L g550 ( 
.A(n_542),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_260),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_115),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_152),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_226),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_494),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_13),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_40),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_204),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_218),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_241),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_492),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_548),
.Y(n_562)
);

BUFx10_ASAP7_75t_L g563 ( 
.A(n_2),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_214),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_186),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_501),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_187),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_118),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_80),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_515),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_255),
.Y(n_571)
);

BUFx10_ASAP7_75t_L g572 ( 
.A(n_380),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_398),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_446),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_532),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_335),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_522),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_43),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_546),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_445),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_138),
.Y(n_581)
);

INVx1_ASAP7_75t_SL g582 ( 
.A(n_110),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_219),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_497),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_41),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_422),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_339),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_253),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_47),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_259),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_477),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_457),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_4),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_426),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_471),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_549),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_229),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_125),
.Y(n_598)
);

CKINVDCx16_ASAP7_75t_R g599 ( 
.A(n_325),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_421),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_235),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_313),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_60),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_528),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_35),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_294),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_403),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_7),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_289),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_50),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_289),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_124),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_328),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_140),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_418),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_383),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_133),
.Y(n_617)
);

CKINVDCx14_ASAP7_75t_R g618 ( 
.A(n_505),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_14),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_479),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_28),
.Y(n_621)
);

BUFx2_ASAP7_75t_SL g622 ( 
.A(n_366),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_392),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_411),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_43),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_400),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_419),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_434),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_164),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_443),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_343),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_78),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_355),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_197),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_238),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_390),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_90),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_539),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_30),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_370),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_506),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_437),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_152),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_97),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_534),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_71),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_203),
.Y(n_648)
);

BUFx8_ASAP7_75t_SL g649 ( 
.A(n_507),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_480),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_473),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_219),
.Y(n_652)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_531),
.Y(n_653)
);

INVx1_ASAP7_75t_SL g654 ( 
.A(n_236),
.Y(n_654)
);

BUFx10_ASAP7_75t_L g655 ( 
.A(n_313),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_397),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_387),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_389),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_358),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_346),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_114),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_524),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_116),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_305),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_243),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_350),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_485),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_130),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_169),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_283),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_301),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_367),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_263),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_36),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_38),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_173),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_394),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_23),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_55),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_29),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_291),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_45),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_502),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_171),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_35),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_227),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_529),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_302),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_424),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_61),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_326),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_412),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_530),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_255),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_206),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_503),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_133),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_264),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_87),
.Y(n_699)
);

CKINVDCx20_ASAP7_75t_R g700 ( 
.A(n_48),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_535),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_368),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_294),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_423),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_472),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_358),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_25),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_511),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_230),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_319),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_514),
.Y(n_711)
);

CKINVDCx16_ASAP7_75t_R g712 ( 
.A(n_428),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_495),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_91),
.Y(n_714)
);

CKINVDCx16_ASAP7_75t_R g715 ( 
.A(n_543),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_410),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_422),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_226),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_153),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_201),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_388),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_343),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_486),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_425),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_220),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_13),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_80),
.Y(n_727)
);

CKINVDCx16_ASAP7_75t_R g728 ( 
.A(n_533),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_424),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_359),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_487),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_250),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_541),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_20),
.Y(n_734)
);

HB1xp67_ASAP7_75t_L g735 ( 
.A(n_160),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_526),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_163),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_253),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_415),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_78),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_265),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_399),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_398),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_238),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_440),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_134),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_454),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_217),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_427),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_240),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_153),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_540),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_537),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_496),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_55),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_230),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_468),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_169),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_425),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_342),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_47),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_212),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_470),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_527),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_536),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_99),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_210),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_198),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_282),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_420),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_95),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_484),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_268),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_439),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_189),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_504),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_547),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_463),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_574),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_571),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_571),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_599),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_588),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_588),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_589),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_589),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_560),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_668),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_668),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_681),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_681),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_560),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_560),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_560),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_623),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_623),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_623),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_623),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_631),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_631),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_631),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_631),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_640),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_557),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_678),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_712),
.Y(n_806)
);

INVxp33_ASAP7_75t_SL g807 ( 
.A(n_735),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_678),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_678),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_678),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_695),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_695),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_567),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_567),
.Y(n_814)
);

NOR2xp67_ASAP7_75t_L g815 ( 
.A(n_597),
.B(n_0),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_551),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_695),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_695),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_552),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_556),
.B(n_0),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_672),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_553),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_564),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_574),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_672),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_565),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_568),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_581),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_583),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_690),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_593),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_554),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_563),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_557),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_594),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_559),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_690),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_653),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_702),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_612),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_613),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_616),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_653),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_626),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_632),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_647),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_665),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_669),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_670),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_671),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_673),
.Y(n_851)
);

HB1xp67_ASAP7_75t_L g852 ( 
.A(n_568),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_611),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_676),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_679),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_711),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_680),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_685),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_597),
.B(n_1),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_569),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_686),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_576),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_688),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_689),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_691),
.Y(n_865)
);

CKINVDCx14_ASAP7_75t_R g866 ( 
.A(n_618),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_692),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_578),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_569),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_698),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_706),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_707),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_586),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_702),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_587),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_709),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_816),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_811),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_824),
.B(n_711),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_804),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_812),
.Y(n_881)
);

NOR2xp67_ASAP7_75t_L g882 ( 
.A(n_816),
.B(n_550),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_555),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_817),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_866),
.Y(n_885)
);

INVxp33_ASAP7_75t_SL g886 ( 
.A(n_803),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_818),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_787),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_822),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_832),
.Y(n_890)
);

INVxp67_ASAP7_75t_SL g891 ( 
.A(n_779),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_832),
.B(n_715),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_787),
.Y(n_893)
);

INVxp33_ASAP7_75t_L g894 ( 
.A(n_813),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_804),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_798),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_834),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_836),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_798),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_834),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_782),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_836),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_862),
.Y(n_903)
);

NOR2xp67_ASAP7_75t_L g904 ( 
.A(n_862),
.B(n_561),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_808),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_868),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_868),
.B(n_728),
.Y(n_907)
);

BUFx6f_ASAP7_75t_SL g908 ( 
.A(n_779),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_808),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_810),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_810),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_873),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_792),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_792),
.Y(n_914)
);

CKINVDCx16_ASAP7_75t_R g915 ( 
.A(n_853),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_853),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_875),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_875),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_793),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_793),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_803),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_833),
.B(n_566),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_794),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_795),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_806),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_806),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_852),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_795),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_807),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_807),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_814),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_814),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_796),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_797),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_797),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_827),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_799),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_827),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_913),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_891),
.B(n_757),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_894),
.B(n_892),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_914),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_879),
.B(n_856),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_919),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_907),
.A2(n_595),
.B1(n_683),
.B2(n_575),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_923),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_927),
.B(n_860),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_901),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_933),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_882),
.B(n_883),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_904),
.B(n_757),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_934),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_931),
.A2(n_932),
.B1(n_886),
.B2(n_930),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_935),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_878),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_936),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_877),
.B(n_869),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_919),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_881),
.Y(n_960)
);

AND2x6_ASAP7_75t_L g961 ( 
.A(n_888),
.B(n_650),
.Y(n_961)
);

BUFx8_ASAP7_75t_L g962 ( 
.A(n_908),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_884),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_887),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_920),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_893),
.B(n_799),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_896),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_920),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_899),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_885),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_885),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_924),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_905),
.B(n_800),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_909),
.Y(n_974)
);

BUFx8_ASAP7_75t_L g975 ( 
.A(n_908),
.Y(n_975)
);

BUFx8_ASAP7_75t_L g976 ( 
.A(n_908),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_910),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_924),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_911),
.Y(n_980)
);

CKINVDCx16_ASAP7_75t_R g981 ( 
.A(n_915),
.Y(n_981)
);

CKINVDCx8_ASAP7_75t_R g982 ( 
.A(n_921),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_937),
.Y(n_983)
);

AND2x4_ASAP7_75t_L g984 ( 
.A(n_922),
.B(n_777),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_931),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_932),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_889),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_890),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_898),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_902),
.Y(n_990)
);

NOR2x1_ASAP7_75t_L g991 ( 
.A(n_926),
.B(n_838),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_925),
.Y(n_992)
);

AOI22xp5_ASAP7_75t_L g993 ( 
.A1(n_886),
.A2(n_595),
.B1(n_683),
.B2(n_575),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_903),
.A2(n_815),
.B1(n_859),
.B2(n_663),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_906),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_880),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_912),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_L g998 ( 
.A(n_929),
.B(n_650),
.Y(n_998)
);

AND2x6_ASAP7_75t_L g999 ( 
.A(n_917),
.B(n_713),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_918),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_938),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_938),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_926),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_916),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_880),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_895),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_895),
.Y(n_1007)
);

INVxp67_ASAP7_75t_L g1008 ( 
.A(n_916),
.Y(n_1008)
);

AND2x2_ASAP7_75t_SL g1009 ( 
.A(n_897),
.B(n_713),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_897),
.B(n_838),
.Y(n_1010)
);

OA21x2_ASAP7_75t_L g1011 ( 
.A1(n_900),
.A2(n_802),
.B(n_801),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_919),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_913),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_919),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_919),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_894),
.B(n_843),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_891),
.B(n_777),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_919),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_913),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_SL g1020 ( 
.A1(n_936),
.A2(n_614),
.B1(n_645),
.B2(n_611),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_913),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_879),
.A2(n_754),
.B(n_620),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_953),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_944),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_944),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_941),
.B(n_754),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_979),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_942),
.B(n_651),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_959),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_1016),
.B(n_843),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_959),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_SL g1032 ( 
.A(n_1009),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_965),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_956),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_960),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_965),
.Y(n_1036)
);

INVx4_ASAP7_75t_L g1037 ( 
.A(n_979),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_947),
.B(n_791),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_968),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_958),
.B(n_791),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_1011),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_963),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_964),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_968),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1011),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_943),
.B(n_701),
.Y(n_1046)
);

INVx8_ASAP7_75t_L g1047 ( 
.A(n_999),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_998),
.B(n_781),
.C(n_780),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_972),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_939),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_946),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_972),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_978),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_942),
.B(n_592),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_942),
.B(n_628),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_949),
.B(n_584),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_978),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_983),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_985),
.B(n_783),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_1013),
.B(n_643),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1012),
.Y(n_1061)
);

CKINVDCx6p67_ASAP7_75t_R g1062 ( 
.A(n_981),
.Y(n_1062)
);

INVx2_ASAP7_75t_SL g1063 ( 
.A(n_1011),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_940),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_942),
.B(n_667),
.Y(n_1065)
);

INVxp67_ASAP7_75t_SL g1066 ( 
.A(n_979),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_948),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_985),
.B(n_784),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_948),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_1012),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_1010),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_961),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1014),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_950),
.B(n_687),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1014),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1015),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_951),
.B(n_945),
.Y(n_1077)
);

OR2x6_ASAP7_75t_L g1078 ( 
.A(n_988),
.B(n_820),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_953),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1015),
.Y(n_1080)
);

NOR3xp33_ASAP7_75t_L g1081 ( 
.A(n_1020),
.B(n_582),
.C(n_558),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_962),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1021),
.B(n_696),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1018),
.Y(n_1084)
);

NAND3x1_ASAP7_75t_L g1085 ( 
.A(n_993),
.B(n_718),
.C(n_717),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1018),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_982),
.B(n_649),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1018),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_1005),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_986),
.B(n_785),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_979),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_967),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_950),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_940),
.B(n_705),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_969),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_974),
.Y(n_1096)
);

OAI21xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1022),
.A2(n_1009),
.B(n_986),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_977),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_1004),
.B(n_786),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_980),
.Y(n_1100)
);

OR2x6_ASAP7_75t_L g1101 ( 
.A(n_988),
.B(n_820),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_950),
.B(n_733),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_940),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_966),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_950),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_973),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_955),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_1017),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_955),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_955),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_998),
.B(n_994),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1017),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_970),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_987),
.B(n_570),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_952),
.B(n_955),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1019),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_989),
.B(n_570),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1019),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1019),
.B(n_747),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1019),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_961),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_984),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_961),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_952),
.B(n_763),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_961),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_984),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_961),
.Y(n_1127)
);

AO21x2_ASAP7_75t_L g1128 ( 
.A1(n_995),
.A2(n_778),
.B(n_805),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_995),
.B(n_562),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_997),
.B(n_622),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_999),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_999),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_999),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_999),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_997),
.B(n_577),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1000),
.B(n_579),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1000),
.Y(n_1137)
);

NAND2xp33_ASAP7_75t_L g1138 ( 
.A(n_991),
.B(n_764),
.Y(n_1138)
);

NAND3xp33_ASAP7_75t_L g1139 ( 
.A(n_954),
.B(n_789),
.C(n_788),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_990),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_990),
.Y(n_1141)
);

BUFx10_ASAP7_75t_L g1142 ( 
.A(n_970),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_982),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_992),
.B(n_765),
.Y(n_1144)
);

INVx8_ASAP7_75t_L g1145 ( 
.A(n_971),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_962),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_962),
.Y(n_1147)
);

INVx1_ASAP7_75t_SL g1148 ( 
.A(n_996),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_975),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_992),
.B(n_580),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1003),
.Y(n_1151)
);

INVx4_ASAP7_75t_SL g1152 ( 
.A(n_1032),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1046),
.B(n_591),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1029),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_1089),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1062),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1111),
.A2(n_1003),
.B1(n_642),
.B2(n_645),
.Y(n_1157)
);

BUFx2_ASAP7_75t_L g1158 ( 
.A(n_1148),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_1062),
.Y(n_1159)
);

INVx8_ASAP7_75t_L g1160 ( 
.A(n_1145),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1023),
.Y(n_1161)
);

OR2x6_ASAP7_75t_L g1162 ( 
.A(n_1145),
.B(n_1005),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_1038),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1029),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1040),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1033),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1030),
.B(n_1002),
.Y(n_1167)
);

AND2x6_ASAP7_75t_L g1168 ( 
.A(n_1131),
.B(n_1005),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1033),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1036),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1079),
.B(n_1005),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1036),
.Y(n_1172)
);

INVx4_ASAP7_75t_SL g1173 ( 
.A(n_1032),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1039),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1039),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1023),
.B(n_971),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_1130),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1049),
.Y(n_1178)
);

INVxp33_ASAP7_75t_L g1179 ( 
.A(n_1099),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_1023),
.B(n_975),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_1130),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1023),
.B(n_975),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1049),
.Y(n_1183)
);

BUFx10_ASAP7_75t_L g1184 ( 
.A(n_1144),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1079),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1130),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1077),
.B(n_1008),
.Y(n_1187)
);

BUFx2_ASAP7_75t_L g1188 ( 
.A(n_1130),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1145),
.Y(n_1189)
);

INVxp67_ASAP7_75t_L g1190 ( 
.A(n_1078),
.Y(n_1190)
);

OR2x6_ASAP7_75t_L g1191 ( 
.A(n_1145),
.B(n_1006),
.Y(n_1191)
);

OAI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1064),
.A2(n_656),
.B1(n_700),
.B2(n_614),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1104),
.B(n_1106),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_1108),
.B(n_1006),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1093),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1067),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1104),
.B(n_596),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1067),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1137),
.B(n_976),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1064),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_1151),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1041),
.A2(n_642),
.B1(n_700),
.B2(n_656),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1071),
.Y(n_1203)
);

INVx1_ASAP7_75t_SL g1204 ( 
.A(n_1069),
.Y(n_1204)
);

INVxp67_ASAP7_75t_SL g1205 ( 
.A(n_1093),
.Y(n_1205)
);

AND2x2_ASAP7_75t_SL g1206 ( 
.A(n_1087),
.B(n_1006),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1103),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1052),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_L g1209 ( 
.A(n_1137),
.B(n_1001),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1069),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1053),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1057),
.Y(n_1212)
);

BUFx4f_ASAP7_75t_L g1213 ( 
.A(n_1143),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1106),
.B(n_604),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1057),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1103),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1140),
.Y(n_1217)
);

INVx4_ASAP7_75t_L g1218 ( 
.A(n_1093),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1058),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_L g1220 ( 
.A(n_1140),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1141),
.B(n_1006),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_1131),
.B(n_1007),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1141),
.B(n_1007),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1113),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1112),
.B(n_630),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1061),
.Y(n_1226)
);

INVx4_ASAP7_75t_SL g1227 ( 
.A(n_1032),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1061),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1059),
.B(n_638),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1070),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_1113),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1142),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1073),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1073),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1114),
.B(n_976),
.Y(n_1235)
);

NAND2x1p5_ASAP7_75t_L g1236 ( 
.A(n_1105),
.B(n_1002),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1105),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1075),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1091),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1109),
.Y(n_1240)
);

INVx6_ASAP7_75t_L g1241 ( 
.A(n_1142),
.Y(n_1241)
);

NAND2xp33_ASAP7_75t_L g1242 ( 
.A(n_1047),
.B(n_641),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1068),
.B(n_646),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1076),
.Y(n_1244)
);

HB1xp67_ASAP7_75t_L g1245 ( 
.A(n_1078),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1050),
.B(n_662),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1078),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1076),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1051),
.B(n_693),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1078),
.Y(n_1250)
);

HB1xp67_ASAP7_75t_L g1251 ( 
.A(n_1101),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1101),
.B(n_1002),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1080),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1080),
.Y(n_1254)
);

NAND2x1p5_ASAP7_75t_L g1255 ( 
.A(n_1105),
.B(n_1002),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1024),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1034),
.B(n_819),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1035),
.B(n_823),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1109),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1091),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1042),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1026),
.A2(n_720),
.B(n_666),
.C(n_585),
.Y(n_1262)
);

INVxp67_ASAP7_75t_SL g1263 ( 
.A(n_1107),
.Y(n_1263)
);

AND2x6_ASAP7_75t_L g1264 ( 
.A(n_1132),
.B(n_726),
.Y(n_1264)
);

INVx1_ASAP7_75t_SL g1265 ( 
.A(n_1090),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1092),
.B(n_708),
.Y(n_1266)
);

INVx2_ASAP7_75t_SL g1267 ( 
.A(n_1101),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1101),
.B(n_957),
.Y(n_1268)
);

INVxp67_ASAP7_75t_L g1269 ( 
.A(n_1117),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1150),
.B(n_996),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1098),
.B(n_723),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1142),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1043),
.B(n_1122),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1024),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1110),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1098),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1126),
.B(n_731),
.Y(n_1277)
);

INVx4_ASAP7_75t_L g1278 ( 
.A(n_1107),
.Y(n_1278)
);

AND2x4_ASAP7_75t_L g1279 ( 
.A(n_1095),
.B(n_826),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1096),
.Y(n_1280)
);

AND2x6_ASAP7_75t_L g1281 ( 
.A(n_1132),
.B(n_726),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1100),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1025),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1085),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1031),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1031),
.Y(n_1286)
);

AND2x6_ASAP7_75t_L g1287 ( 
.A(n_1133),
.B(n_761),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1044),
.Y(n_1288)
);

BUFx6f_ASAP7_75t_L g1289 ( 
.A(n_1110),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1136),
.B(n_737),
.Y(n_1290)
);

AND2x2_ASAP7_75t_L g1291 ( 
.A(n_1026),
.B(n_790),
.Y(n_1291)
);

AO22x2_ASAP7_75t_L g1292 ( 
.A1(n_1081),
.A2(n_1045),
.B1(n_1063),
.B2(n_1041),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1044),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_SL g1294 ( 
.A(n_1115),
.B(n_976),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1139),
.B(n_828),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1129),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1045),
.A2(n_1063),
.B1(n_1128),
.B2(n_1094),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1044),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1084),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1084),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1086),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1135),
.B(n_737),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1086),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1088),
.Y(n_1304)
);

BUFx10_ASAP7_75t_L g1305 ( 
.A(n_1138),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1085),
.A2(n_720),
.B1(n_666),
.B2(n_610),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1135),
.B(n_572),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1088),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1138),
.B(n_572),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1056),
.B(n_736),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1028),
.B(n_755),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1116),
.B(n_829),
.Y(n_1312)
);

AO22x2_ASAP7_75t_L g1313 ( 
.A1(n_1146),
.A2(n_654),
.B1(n_748),
.B2(n_761),
.Y(n_1313)
);

INVx6_ASAP7_75t_L g1314 ( 
.A(n_1082),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1118),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1028),
.B(n_572),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1120),
.Y(n_1317)
);

OR2x2_ASAP7_75t_L g1318 ( 
.A(n_1048),
.B(n_831),
.Y(n_1318)
);

CKINVDCx14_ASAP7_75t_R g1319 ( 
.A(n_1082),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1120),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1107),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1146),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1060),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1072),
.B(n_765),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1047),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1072),
.B(n_745),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1027),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1124),
.B(n_767),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1265),
.B(n_1124),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1224),
.Y(n_1330)
);

BUFx6f_ASAP7_75t_L g1331 ( 
.A(n_1161),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1193),
.B(n_1083),
.Y(n_1332)
);

BUFx10_ASAP7_75t_L g1333 ( 
.A(n_1210),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1226),
.Y(n_1334)
);

O2A1O1Ixp5_ASAP7_75t_L g1335 ( 
.A1(n_1153),
.A2(n_1134),
.B(n_1133),
.C(n_1055),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1269),
.B(n_1147),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1290),
.A2(n_1097),
.B(n_1055),
.C(n_1065),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1323),
.B(n_1187),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1302),
.B(n_1147),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1323),
.B(n_1066),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1226),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1179),
.B(n_1311),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1314),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1254),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1291),
.B(n_1027),
.Y(n_1345)
);

OAI221xp5_ASAP7_75t_L g1346 ( 
.A1(n_1328),
.A2(n_1149),
.B1(n_760),
.B2(n_762),
.C(n_756),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1209),
.B(n_1037),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_1296),
.B(n_1072),
.Y(n_1348)
);

AOI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1167),
.A2(n_1134),
.B1(n_1054),
.B2(n_1074),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1270),
.A2(n_1054),
.B1(n_1074),
.B2(n_1065),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1164),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1165),
.B(n_1149),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1163),
.B(n_1192),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1261),
.Y(n_1354)
);

INVx8_ASAP7_75t_L g1355 ( 
.A(n_1160),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1221),
.A2(n_1102),
.B1(n_1119),
.B2(n_1121),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1166),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1280),
.B(n_1282),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1197),
.B(n_1037),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1175),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1214),
.B(n_1102),
.Y(n_1361)
);

AND2x6_ASAP7_75t_L g1362 ( 
.A(n_1327),
.B(n_1121),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1185),
.B(n_1213),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1276),
.B(n_1123),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1273),
.A2(n_1125),
.B1(n_1127),
.B2(n_1123),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1195),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1215),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1229),
.B(n_1125),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1154),
.Y(n_1369)
);

INVx2_ASAP7_75t_SL g1370 ( 
.A(n_1203),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1184),
.B(n_1127),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1243),
.B(n_752),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_753),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1185),
.B(n_772),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1312),
.B(n_774),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1312),
.B(n_776),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1273),
.B(n_590),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1217),
.B(n_598),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1161),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1221),
.B(n_835),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1160),
.B(n_1162),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1231),
.A2(n_760),
.B1(n_756),
.B2(n_573),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1217),
.B(n_600),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1220),
.B(n_601),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1169),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1219),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1220),
.B(n_602),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1170),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1292),
.A2(n_1295),
.B1(n_1307),
.B2(n_1202),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1220),
.B(n_603),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1267),
.A2(n_841),
.B1(n_842),
.B2(n_840),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1172),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1200),
.B(n_605),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1200),
.B(n_606),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1200),
.B(n_1207),
.Y(n_1395)
);

AOI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1190),
.A2(n_1252),
.B1(n_1309),
.B2(n_1223),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1207),
.B(n_607),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1207),
.B(n_608),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1216),
.B(n_609),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1216),
.B(n_615),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1213),
.B(n_844),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_SL g1402 ( 
.A(n_1216),
.B(n_845),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1218),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1297),
.A2(n_617),
.B1(n_621),
.B2(n_619),
.Y(n_1404)
);

NAND2xp33_ASAP7_75t_L g1405 ( 
.A(n_1168),
.B(n_573),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1316),
.B(n_624),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1184),
.B(n_846),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1201),
.B(n_625),
.Y(n_1408)
);

INVx8_ASAP7_75t_L g1409 ( 
.A(n_1162),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1257),
.B(n_627),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1174),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1257),
.B(n_629),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1178),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1183),
.Y(n_1414)
);

INVx8_ASAP7_75t_L g1415 ( 
.A(n_1191),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1258),
.B(n_633),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1258),
.B(n_634),
.Y(n_1417)
);

INVxp67_ASAP7_75t_L g1418 ( 
.A(n_1158),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1279),
.B(n_635),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1208),
.Y(n_1420)
);

INVxp67_ASAP7_75t_L g1421 ( 
.A(n_1155),
.Y(n_1421)
);

INVx8_ASAP7_75t_L g1422 ( 
.A(n_1191),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1292),
.A2(n_649),
.B1(n_721),
.B2(n_719),
.Y(n_1423)
);

BUFx6f_ASAP7_75t_L g1424 ( 
.A(n_1161),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1171),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1279),
.B(n_636),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1171),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1194),
.B(n_847),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1194),
.B(n_848),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1295),
.B(n_637),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_1294),
.B(n_850),
.C(n_849),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1156),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1223),
.A2(n_854),
.B1(n_855),
.B2(n_851),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1248),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1253),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1189),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1159),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1222),
.B(n_639),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1256),
.Y(n_1439)
);

NOR2xp67_ASAP7_75t_L g1440 ( 
.A(n_1235),
.B(n_429),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1222),
.B(n_644),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1322),
.B(n_857),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1268),
.A2(n_1250),
.B1(n_1247),
.B2(n_1176),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1211),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1212),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1177),
.Y(n_1446)
);

INVxp67_ASAP7_75t_SL g1447 ( 
.A(n_1240),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_SL g1448 ( 
.A(n_1206),
.B(n_1305),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_SL g1449 ( 
.A(n_1305),
.B(n_858),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1181),
.B(n_861),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1222),
.B(n_648),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1196),
.B(n_652),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_L g1453 ( 
.A(n_1168),
.B(n_762),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1198),
.B(n_657),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1222),
.B(n_658),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1228),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1152),
.B(n_863),
.Y(n_1457)
);

A2O1A1Ixp33_ASAP7_75t_L g1458 ( 
.A1(n_1262),
.A2(n_725),
.B(n_749),
.C(n_722),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1230),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1233),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1152),
.B(n_864),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1204),
.B(n_659),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1186),
.B(n_865),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1234),
.Y(n_1464)
);

AND2x6_ASAP7_75t_L g1465 ( 
.A(n_1240),
.B(n_758),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1245),
.A2(n_870),
.B1(n_871),
.B2(n_867),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1238),
.Y(n_1467)
);

INVx5_ASAP7_75t_L g1468 ( 
.A(n_1241),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_SL g1469 ( 
.A(n_1241),
.B(n_655),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1168),
.B(n_660),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1284),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1244),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1188),
.B(n_872),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1251),
.A2(n_876),
.B1(n_661),
.B2(n_664),
.Y(n_1474)
);

BUFx5_ASAP7_75t_L g1475 ( 
.A(n_1264),
.Y(n_1475)
);

NOR2xp67_ASAP7_75t_L g1476 ( 
.A(n_1225),
.B(n_430),
.Y(n_1476)
);

O2A1O1Ixp5_ASAP7_75t_L g1477 ( 
.A1(n_1324),
.A2(n_759),
.B(n_768),
.C(n_750),
.Y(n_1477)
);

O2A1O1Ixp33_ASAP7_75t_L g1478 ( 
.A1(n_1199),
.A2(n_1271),
.B(n_1266),
.C(n_1249),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1173),
.B(n_874),
.Y(n_1479)
);

AND2x4_ASAP7_75t_SL g1480 ( 
.A(n_1240),
.B(n_655),
.Y(n_1480)
);

NAND2xp33_ASAP7_75t_L g1481 ( 
.A(n_1168),
.B(n_766),
.Y(n_1481)
);

NOR2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1232),
.B(n_766),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1157),
.B(n_655),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1236),
.B(n_821),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1246),
.B(n_674),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1255),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1299),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1315),
.B(n_675),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1173),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1325),
.A2(n_682),
.B1(n_684),
.B2(n_677),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1325),
.B(n_1218),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1300),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1301),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1227),
.B(n_694),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1227),
.B(n_697),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1272),
.B(n_699),
.Y(n_1496)
);

AOI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1277),
.A2(n_704),
.B1(n_710),
.B2(n_703),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1303),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1317),
.B(n_714),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1320),
.B(n_716),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1304),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1205),
.B(n_724),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_SL g1503 ( 
.A(n_1259),
.B(n_727),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1308),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1313),
.A2(n_1306),
.B1(n_775),
.B2(n_771),
.C(n_732),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1259),
.B(n_729),
.Y(n_1506)
);

INVxp67_ASAP7_75t_L g1507 ( 
.A(n_1313),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1319),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1418),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1353),
.A2(n_1306),
.B1(n_1182),
.B2(n_1180),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1354),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1338),
.B(n_1318),
.Y(n_1512)
);

INVx4_ASAP7_75t_L g1513 ( 
.A(n_1468),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1342),
.B(n_1272),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1334),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1341),
.Y(n_1516)
);

INVx2_ASAP7_75t_SL g1517 ( 
.A(n_1343),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1358),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1330),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1329),
.Y(n_1520)
);

INVx2_ASAP7_75t_SL g1521 ( 
.A(n_1468),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1339),
.B(n_1259),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1369),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1468),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1421),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1385),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1366),
.Y(n_1527)
);

INVxp67_ASAP7_75t_L g1528 ( 
.A(n_1352),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1485),
.B(n_1321),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1388),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_SL g1531 ( 
.A(n_1436),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1436),
.B(n_1237),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_SL g1533 ( 
.A(n_1336),
.B(n_1275),
.Y(n_1533)
);

CKINVDCx11_ASAP7_75t_R g1534 ( 
.A(n_1489),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1332),
.B(n_1263),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1446),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1344),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1392),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1389),
.B(n_1275),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1471),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1439),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1508),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1425),
.B(n_1427),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1340),
.B(n_1275),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1355),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1370),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_SL g1547 ( 
.A(n_1346),
.B(n_734),
.C(n_730),
.Y(n_1547)
);

NOR3xp33_ASAP7_75t_SL g1548 ( 
.A(n_1448),
.B(n_739),
.C(n_738),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_1442),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1411),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1333),
.Y(n_1551)
);

INVx5_ASAP7_75t_L g1552 ( 
.A(n_1381),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1382),
.A2(n_741),
.B1(n_742),
.B2(n_740),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_SL g1554 ( 
.A(n_1452),
.B(n_1289),
.Y(n_1554)
);

NAND3xp33_ASAP7_75t_SL g1555 ( 
.A(n_1483),
.B(n_744),
.C(n_743),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_SL g1556 ( 
.A(n_1454),
.B(n_1289),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1413),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1380),
.B(n_1274),
.Y(n_1558)
);

NOR2xp33_ASAP7_75t_R g1559 ( 
.A(n_1432),
.B(n_1239),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1333),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1414),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1406),
.B(n_1396),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1403),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1381),
.B(n_1237),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1372),
.B(n_1283),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1462),
.B(n_1260),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1469),
.B(n_1278),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1442),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1380),
.A2(n_1281),
.B1(n_1287),
.B2(n_1264),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1420),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1459),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1373),
.B(n_1285),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1430),
.B(n_1410),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1363),
.B(n_1278),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1460),
.Y(n_1575)
);

AND2x4_ASAP7_75t_SL g1576 ( 
.A(n_1436),
.B(n_1260),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1361),
.B(n_1288),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1444),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1335),
.A2(n_1281),
.B(n_1264),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1443),
.B(n_1286),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1505),
.A2(n_1281),
.B1(n_1287),
.B2(n_1293),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1449),
.B(n_1298),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_SL g1583 ( 
.A(n_1496),
.B(n_1326),
.Y(n_1583)
);

NOR2x2_ASAP7_75t_L g1584 ( 
.A(n_1445),
.B(n_821),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1480),
.B(n_825),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1408),
.B(n_746),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1494),
.B(n_769),
.C(n_751),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1355),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1491),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1467),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1345),
.B(n_1242),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1378),
.B(n_825),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1383),
.B(n_830),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1472),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_SL g1595 ( 
.A(n_1393),
.B(n_770),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1437),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1404),
.A2(n_773),
.B1(n_837),
.B2(n_830),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1384),
.B(n_837),
.Y(n_1598)
);

INVx3_ASAP7_75t_SL g1599 ( 
.A(n_1457),
.Y(n_1599)
);

AO21x1_ASAP7_75t_L g1600 ( 
.A1(n_1337),
.A2(n_809),
.B(n_839),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1507),
.B(n_2),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1409),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1487),
.Y(n_1603)
);

NOR2x2_ASAP7_75t_L g1604 ( 
.A(n_1456),
.B(n_3),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_SL g1605 ( 
.A(n_1394),
.B(n_3),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1331),
.Y(n_1606)
);

INVx2_ASAP7_75t_SL g1607 ( 
.A(n_1409),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1482),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1415),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1407),
.B(n_4),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1412),
.B(n_1416),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1331),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1347),
.B(n_5),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1415),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1417),
.B(n_5),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1331),
.Y(n_1616)
);

INVx3_ASAP7_75t_L g1617 ( 
.A(n_1379),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1431),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1501),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1379),
.Y(n_1620)
);

INVx2_ASAP7_75t_SL g1621 ( 
.A(n_1422),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1397),
.B(n_6),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1368),
.B(n_8),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1423),
.B(n_9),
.C(n_10),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1464),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1492),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1398),
.B(n_9),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1493),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1399),
.B(n_10),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1395),
.B(n_1486),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1498),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1422),
.Y(n_1632)
);

OR2x6_ASAP7_75t_L g1633 ( 
.A(n_1379),
.B(n_431),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1351),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1428),
.A2(n_14),
.B1(n_11),
.B2(n_12),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1461),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1504),
.B(n_11),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1357),
.Y(n_1638)
);

INVxp67_ASAP7_75t_L g1639 ( 
.A(n_1377),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1400),
.B(n_15),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_L g1641 ( 
.A1(n_1429),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1641)
);

AND2x4_ASAP7_75t_L g1642 ( 
.A(n_1402),
.B(n_432),
.Y(n_1642)
);

BUFx12f_ASAP7_75t_SL g1643 ( 
.A(n_1479),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1360),
.Y(n_1644)
);

O2A1O1Ixp33_ASAP7_75t_L g1645 ( 
.A1(n_1401),
.A2(n_1458),
.B(n_1478),
.C(n_1426),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1350),
.B(n_16),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1367),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_SL g1648 ( 
.A(n_1440),
.B(n_17),
.Y(n_1648)
);

AOI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1419),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_1649)
);

INVx4_ASAP7_75t_L g1650 ( 
.A(n_1424),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1386),
.Y(n_1651)
);

NOR2xp33_ASAP7_75t_L g1652 ( 
.A(n_1450),
.B(n_18),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1365),
.A2(n_22),
.B1(n_19),
.B2(n_21),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1447),
.B(n_1482),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1387),
.B(n_21),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1434),
.B(n_22),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1435),
.Y(n_1657)
);

AOI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1463),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1390),
.B(n_24),
.Y(n_1659)
);

AND2x4_ASAP7_75t_L g1660 ( 
.A(n_1503),
.B(n_433),
.Y(n_1660)
);

CKINVDCx11_ASAP7_75t_R g1661 ( 
.A(n_1424),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1495),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_L g1663 ( 
.A(n_1473),
.B(n_26),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1484),
.Y(n_1664)
);

INVx1_ASAP7_75t_SL g1665 ( 
.A(n_1502),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1371),
.B(n_26),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1474),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1424),
.Y(n_1668)
);

CKINVDCx11_ASAP7_75t_R g1669 ( 
.A(n_1475),
.Y(n_1669)
);

BUFx4f_ASAP7_75t_L g1670 ( 
.A(n_1465),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1465),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1506),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1364),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1488),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1499),
.B(n_27),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_SL g1676 ( 
.A(n_1466),
.B(n_27),
.Y(n_1676)
);

BUFx6f_ASAP7_75t_L g1677 ( 
.A(n_1661),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1512),
.B(n_1497),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1511),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1518),
.B(n_1375),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1578),
.Y(n_1681)
);

A2O1A1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1645),
.A2(n_1476),
.B(n_1477),
.C(n_1359),
.Y(n_1682)
);

AOI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1667),
.A2(n_1374),
.B1(n_1476),
.B2(n_1376),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1523),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1520),
.B(n_1500),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_L g1686 ( 
.A(n_1555),
.B(n_1490),
.C(n_1441),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1588),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1552),
.B(n_1433),
.Y(n_1688)
);

BUFx8_ASAP7_75t_L g1689 ( 
.A(n_1588),
.Y(n_1689)
);

O2A1O1Ixp5_ASAP7_75t_L g1690 ( 
.A1(n_1646),
.A2(n_1600),
.B(n_1648),
.C(n_1583),
.Y(n_1690)
);

CKINVDCx16_ASAP7_75t_R g1691 ( 
.A(n_1614),
.Y(n_1691)
);

OAI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1579),
.A2(n_1349),
.B(n_1348),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1391),
.Y(n_1693)
);

AOI21xp5_ASAP7_75t_L g1694 ( 
.A1(n_1591),
.A2(n_1481),
.B(n_1453),
.Y(n_1694)
);

NAND2x1p5_ASAP7_75t_L g1695 ( 
.A(n_1513),
.B(n_1356),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1520),
.B(n_1438),
.Y(n_1696)
);

AOI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1535),
.A2(n_1405),
.B(n_1470),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1565),
.A2(n_1455),
.B(n_1451),
.Y(n_1698)
);

BUFx6f_ASAP7_75t_L g1699 ( 
.A(n_1588),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_1536),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1552),
.B(n_1362),
.Y(n_1701)
);

A2O1A1Ixp33_ASAP7_75t_L g1702 ( 
.A1(n_1529),
.A2(n_1475),
.B(n_1362),
.C(n_30),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1586),
.A2(n_1362),
.B(n_1475),
.Y(n_1703)
);

AOI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1572),
.A2(n_1567),
.B(n_1577),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1611),
.B(n_28),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1665),
.B(n_1475),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1547),
.A2(n_1475),
.B1(n_1362),
.B2(n_32),
.Y(n_1707)
);

OA22x2_ASAP7_75t_L g1708 ( 
.A1(n_1649),
.A2(n_32),
.B1(n_29),
.B2(n_31),
.Y(n_1708)
);

O2A1O1Ixp33_ASAP7_75t_SL g1709 ( 
.A1(n_1653),
.A2(n_34),
.B(n_31),
.C(n_33),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1562),
.A2(n_33),
.B(n_34),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1665),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1528),
.B(n_41),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1674),
.B(n_42),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1513),
.Y(n_1714)
);

NOR2xp33_ASAP7_75t_L g1715 ( 
.A(n_1573),
.B(n_435),
.Y(n_1715)
);

AO32x2_ASAP7_75t_L g1716 ( 
.A1(n_1553),
.A2(n_45),
.A3(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1526),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1530),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1640),
.A2(n_48),
.B1(n_44),
.B2(n_46),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1660),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1510),
.A2(n_52),
.B1(n_49),
.B2(n_51),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1639),
.A2(n_52),
.B(n_53),
.Y(n_1722)
);

O2A1O1Ixp5_ASAP7_75t_SL g1723 ( 
.A1(n_1522),
.A2(n_56),
.B(n_53),
.C(n_54),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1538),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1625),
.Y(n_1725)
);

OAI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1649),
.A2(n_57),
.B1(n_54),
.B2(n_56),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1566),
.B(n_57),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1549),
.B(n_1568),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1660),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_SL g1730 ( 
.A(n_1510),
.B(n_58),
.C(n_59),
.Y(n_1730)
);

OR2x2_ASAP7_75t_SL g1731 ( 
.A(n_1624),
.B(n_1672),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1544),
.A2(n_438),
.B(n_436),
.Y(n_1732)
);

INVx1_ASAP7_75t_SL g1733 ( 
.A(n_1540),
.Y(n_1733)
);

BUFx12f_ASAP7_75t_L g1734 ( 
.A(n_1534),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1675),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1545),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1549),
.B(n_62),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1568),
.B(n_63),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1673),
.B(n_1514),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1676),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1630),
.B(n_64),
.Y(n_1741)
);

AND2x6_ASAP7_75t_L g1742 ( 
.A(n_1642),
.B(n_441),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1605),
.A2(n_1627),
.B(n_1629),
.C(n_1622),
.Y(n_1743)
);

OR2x6_ASAP7_75t_L g1744 ( 
.A(n_1633),
.B(n_442),
.Y(n_1744)
);

BUFx12f_ASAP7_75t_L g1745 ( 
.A(n_1519),
.Y(n_1745)
);

BUFx3_ASAP7_75t_L g1746 ( 
.A(n_1602),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1531),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1630),
.B(n_65),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1509),
.Y(n_1749)
);

NOR2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1609),
.B(n_444),
.Y(n_1750)
);

BUFx6f_ASAP7_75t_L g1751 ( 
.A(n_1616),
.Y(n_1751)
);

OAI22x1_ASAP7_75t_L g1752 ( 
.A1(n_1624),
.A2(n_1610),
.B1(n_1659),
.B2(n_1652),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_SL g1753 ( 
.A(n_1672),
.B(n_66),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1539),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1582),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1755)
);

NOR3xp33_ASAP7_75t_L g1756 ( 
.A(n_1553),
.B(n_70),
.C(n_71),
.Y(n_1756)
);

BUFx8_ASAP7_75t_L g1757 ( 
.A(n_1546),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1550),
.Y(n_1758)
);

AOI21xp5_ASAP7_75t_L g1759 ( 
.A1(n_1554),
.A2(n_545),
.B(n_448),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1558),
.B(n_70),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1662),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1672),
.A2(n_75),
.B1(n_72),
.B2(n_73),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1525),
.B(n_75),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1556),
.A2(n_449),
.B(n_447),
.Y(n_1764)
);

A2O1A1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1663),
.A2(n_79),
.B(n_76),
.C(n_77),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1592),
.B(n_76),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1545),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1593),
.B(n_77),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1598),
.B(n_79),
.Y(n_1769)
);

AO21x1_ASAP7_75t_L g1770 ( 
.A1(n_1613),
.A2(n_81),
.B(n_82),
.Y(n_1770)
);

AOI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1533),
.A2(n_544),
.B(n_451),
.Y(n_1771)
);

AOI21x1_ASAP7_75t_L g1772 ( 
.A1(n_1623),
.A2(n_452),
.B(n_450),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1548),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_1773)
);

OAI22xp5_ASAP7_75t_L g1774 ( 
.A1(n_1580),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1655),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1666),
.B(n_86),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1580),
.A2(n_89),
.B1(n_87),
.B2(n_88),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1626),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1628),
.B(n_88),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1631),
.B(n_89),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1596),
.B(n_453),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1595),
.B(n_455),
.Y(n_1782)
);

NOR2xp33_ASAP7_75t_L g1783 ( 
.A(n_1615),
.B(n_456),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1654),
.B(n_90),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1601),
.B(n_91),
.Y(n_1785)
);

CKINVDCx10_ASAP7_75t_R g1786 ( 
.A(n_1633),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1585),
.B(n_92),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1551),
.Y(n_1788)
);

O2A1O1Ixp33_ASAP7_75t_SL g1789 ( 
.A1(n_1637),
.A2(n_94),
.B(n_92),
.C(n_93),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1654),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1517),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1642),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_SL g1793 ( 
.A(n_1643),
.B(n_458),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1656),
.A2(n_460),
.B(n_459),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1515),
.Y(n_1795)
);

NAND2x1p5_ASAP7_75t_L g1796 ( 
.A(n_1564),
.B(n_461),
.Y(n_1796)
);

AOI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1670),
.A2(n_464),
.B(n_462),
.Y(n_1797)
);

AO32x1_ASAP7_75t_L g1798 ( 
.A1(n_1671),
.A2(n_99),
.A3(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_1798)
);

BUFx4f_ASAP7_75t_L g1799 ( 
.A(n_1599),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1527),
.A2(n_538),
.B(n_466),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1616),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1516),
.Y(n_1802)
);

NOR2xp67_ASAP7_75t_L g1803 ( 
.A(n_1560),
.B(n_465),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1587),
.B(n_100),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1559),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1634),
.B(n_101),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1537),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1638),
.B(n_101),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1647),
.B(n_102),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1581),
.A2(n_102),
.B(n_103),
.Y(n_1810)
);

O2A1O1Ixp5_ASAP7_75t_L g1811 ( 
.A1(n_1637),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1557),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1542),
.B(n_467),
.Y(n_1813)
);

NOR2xp67_ASAP7_75t_L g1814 ( 
.A(n_1607),
.B(n_1621),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1541),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1561),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1606),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1581),
.A2(n_110),
.B(n_108),
.C(n_109),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1564),
.B(n_109),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1576),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1657),
.B(n_111),
.Y(n_1821)
);

A2O1A1Ixp33_ASAP7_75t_L g1822 ( 
.A1(n_1618),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_1822)
);

AO21x1_ASAP7_75t_L g1823 ( 
.A1(n_1721),
.A2(n_1656),
.B(n_1571),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1679),
.Y(n_1824)
);

NAND2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1799),
.B(n_1563),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1684),
.Y(n_1826)
);

AND3x4_ASAP7_75t_L g1827 ( 
.A(n_1756),
.B(n_1604),
.C(n_1543),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1697),
.A2(n_1682),
.B(n_1698),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1694),
.A2(n_1704),
.B(n_1703),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1690),
.A2(n_1658),
.B(n_1641),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1728),
.B(n_1701),
.Y(n_1831)
);

INVx4_ASAP7_75t_L g1832 ( 
.A(n_1747),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1810),
.A2(n_1574),
.B(n_1569),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1739),
.B(n_1570),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1696),
.B(n_1575),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_SL g1836 ( 
.A1(n_1770),
.A2(n_1635),
.B(n_1594),
.Y(n_1836)
);

CKINVDCx5p33_ASAP7_75t_R g1837 ( 
.A(n_1745),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1683),
.A2(n_1608),
.B1(n_1636),
.B2(n_1603),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1681),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1680),
.A2(n_1619),
.B(n_1590),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1678),
.B(n_1644),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1702),
.A2(n_1532),
.B(n_1669),
.Y(n_1842)
);

INVx4_ASAP7_75t_L g1843 ( 
.A(n_1677),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1717),
.Y(n_1844)
);

BUFx6f_ASAP7_75t_L g1845 ( 
.A(n_1791),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1706),
.A2(n_1589),
.B(n_1651),
.Y(n_1846)
);

AND2x4_ASAP7_75t_L g1847 ( 
.A(n_1701),
.B(n_1632),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1685),
.B(n_1715),
.Y(n_1848)
);

INVx3_ASAP7_75t_L g1849 ( 
.A(n_1751),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_SL g1850 ( 
.A1(n_1710),
.A2(n_1524),
.B(n_1521),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1731),
.A2(n_1543),
.B1(n_1597),
.B2(n_1606),
.Y(n_1851)
);

OAI21x1_ASAP7_75t_L g1852 ( 
.A1(n_1692),
.A2(n_1617),
.B(n_1612),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1744),
.B(n_1612),
.Y(n_1853)
);

AND2x4_ASAP7_75t_L g1854 ( 
.A(n_1744),
.B(n_1650),
.Y(n_1854)
);

CKINVDCx20_ASAP7_75t_R g1855 ( 
.A(n_1691),
.Y(n_1855)
);

NAND3xp33_ASAP7_75t_L g1856 ( 
.A(n_1722),
.B(n_1719),
.C(n_1765),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1705),
.B(n_1616),
.Y(n_1857)
);

OAI21x1_ASAP7_75t_L g1858 ( 
.A1(n_1794),
.A2(n_1650),
.B(n_1620),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1743),
.A2(n_1620),
.B(n_1668),
.C(n_1584),
.Y(n_1859)
);

NAND2x1_ASAP7_75t_L g1860 ( 
.A(n_1742),
.B(n_1620),
.Y(n_1860)
);

OAI22x1_ASAP7_75t_L g1861 ( 
.A1(n_1761),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1861)
);

OAI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1772),
.A2(n_1668),
.B(n_474),
.Y(n_1862)
);

AOI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1797),
.A2(n_1668),
.B(n_475),
.Y(n_1863)
);

AOI21xp5_ASAP7_75t_L g1864 ( 
.A1(n_1752),
.A2(n_476),
.B(n_469),
.Y(n_1864)
);

BUFx4_ASAP7_75t_SL g1865 ( 
.A(n_1788),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1733),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1709),
.A2(n_481),
.B(n_478),
.Y(n_1867)
);

AND2x4_ASAP7_75t_L g1868 ( 
.A(n_1817),
.B(n_482),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1700),
.B(n_483),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1730),
.A2(n_115),
.B(n_116),
.Y(n_1870)
);

OAI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1707),
.A2(n_117),
.B(n_118),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1751),
.Y(n_1872)
);

BUFx6f_ASAP7_75t_L g1873 ( 
.A(n_1751),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1718),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1724),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1686),
.A2(n_117),
.B(n_119),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1749),
.B(n_119),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1785),
.B(n_488),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1801),
.Y(n_1879)
);

CKINVDCx6p67_ASAP7_75t_R g1880 ( 
.A(n_1734),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1677),
.B(n_489),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1688),
.B(n_490),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1776),
.B(n_120),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1695),
.A2(n_493),
.B(n_491),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1725),
.Y(n_1885)
);

NAND2x1p5_ASAP7_75t_L g1886 ( 
.A(n_1677),
.B(n_498),
.Y(n_1886)
);

AND2x2_ASAP7_75t_SL g1887 ( 
.A(n_1793),
.B(n_120),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1801),
.Y(n_1888)
);

OAI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1822),
.A2(n_121),
.B(n_122),
.Y(n_1889)
);

AOI21xp5_ASAP7_75t_L g1890 ( 
.A1(n_1798),
.A2(n_500),
.B(n_499),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1727),
.B(n_121),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1758),
.Y(n_1892)
);

A2O1A1Ixp33_ASAP7_75t_L g1893 ( 
.A1(n_1740),
.A2(n_124),
.B(n_122),
.C(n_123),
.Y(n_1893)
);

A2O1A1Ixp33_ASAP7_75t_L g1894 ( 
.A1(n_1783),
.A2(n_126),
.B(n_123),
.C(n_125),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1720),
.A2(n_128),
.B1(n_126),
.B2(n_127),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1732),
.A2(n_1818),
.B(n_1764),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_SL g1897 ( 
.A(n_1688),
.B(n_508),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1801),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1693),
.B(n_510),
.Y(n_1899)
);

AOI21xp5_ASAP7_75t_SL g1900 ( 
.A1(n_1773),
.A2(n_513),
.B(n_512),
.Y(n_1900)
);

HB1xp67_ASAP7_75t_L g1901 ( 
.A(n_1795),
.Y(n_1901)
);

AOI21xp5_ASAP7_75t_L g1902 ( 
.A1(n_1759),
.A2(n_517),
.B(n_516),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1778),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1757),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_SL g1905 ( 
.A(n_1782),
.B(n_518),
.Y(n_1905)
);

OAI22x1_ASAP7_75t_L g1906 ( 
.A1(n_1729),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1906)
);

AOI21xp5_ASAP7_75t_L g1907 ( 
.A1(n_1800),
.A2(n_520),
.B(n_519),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1802),
.Y(n_1908)
);

AOI21xp33_ASAP7_75t_L g1909 ( 
.A1(n_1726),
.A2(n_130),
.B(n_131),
.Y(n_1909)
);

AOI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1771),
.A2(n_523),
.B(n_521),
.Y(n_1910)
);

AOI31xp33_ASAP7_75t_L g1911 ( 
.A1(n_1792),
.A2(n_134),
.A3(n_131),
.B(n_132),
.Y(n_1911)
);

NAND2x1p5_ASAP7_75t_L g1912 ( 
.A(n_1736),
.B(n_525),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1757),
.Y(n_1913)
);

O2A1O1Ixp33_ASAP7_75t_L g1914 ( 
.A1(n_1735),
.A2(n_136),
.B(n_132),
.C(n_135),
.Y(n_1914)
);

AO21x1_ASAP7_75t_L g1915 ( 
.A1(n_1775),
.A2(n_135),
.B(n_136),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1807),
.B(n_137),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1811),
.A2(n_137),
.B(n_138),
.Y(n_1917)
);

INVx1_ASAP7_75t_SL g1918 ( 
.A(n_1805),
.Y(n_1918)
);

BUFx3_ASAP7_75t_L g1919 ( 
.A(n_1845),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1824),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1824),
.Y(n_1921)
);

CKINVDCx20_ASAP7_75t_R g1922 ( 
.A(n_1855),
.Y(n_1922)
);

INVx6_ASAP7_75t_SL g1923 ( 
.A(n_1881),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1857),
.B(n_1787),
.Y(n_1924)
);

CKINVDCx16_ASAP7_75t_R g1925 ( 
.A(n_1904),
.Y(n_1925)
);

BUFx2_ASAP7_75t_SL g1926 ( 
.A(n_1913),
.Y(n_1926)
);

BUFx3_ASAP7_75t_L g1927 ( 
.A(n_1845),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1826),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1835),
.B(n_1741),
.Y(n_1929)
);

BUFx12f_ASAP7_75t_L g1930 ( 
.A(n_1837),
.Y(n_1930)
);

BUFx6f_ASAP7_75t_L g1931 ( 
.A(n_1845),
.Y(n_1931)
);

BUFx6f_ASAP7_75t_L g1932 ( 
.A(n_1872),
.Y(n_1932)
);

BUFx2_ASAP7_75t_L g1933 ( 
.A(n_1831),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1826),
.Y(n_1934)
);

AOI22xp5_ASAP7_75t_L g1935 ( 
.A1(n_1856),
.A2(n_1742),
.B1(n_1804),
.B2(n_1784),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1831),
.B(n_1748),
.Y(n_1936)
);

OR2x6_ASAP7_75t_L g1937 ( 
.A(n_1828),
.B(n_1796),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1866),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1874),
.Y(n_1939)
);

INVx4_ASAP7_75t_L g1940 ( 
.A(n_1854),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1874),
.Y(n_1941)
);

CKINVDCx16_ASAP7_75t_R g1942 ( 
.A(n_1843),
.Y(n_1942)
);

INVx4_ASAP7_75t_L g1943 ( 
.A(n_1854),
.Y(n_1943)
);

INVx3_ASAP7_75t_L g1944 ( 
.A(n_1872),
.Y(n_1944)
);

BUFx4f_ASAP7_75t_L g1945 ( 
.A(n_1881),
.Y(n_1945)
);

CKINVDCx16_ASAP7_75t_R g1946 ( 
.A(n_1843),
.Y(n_1946)
);

INVx3_ASAP7_75t_SL g1947 ( 
.A(n_1880),
.Y(n_1947)
);

BUFx3_ASAP7_75t_L g1948 ( 
.A(n_1872),
.Y(n_1948)
);

BUFx12f_ASAP7_75t_L g1949 ( 
.A(n_1832),
.Y(n_1949)
);

INVx2_ASAP7_75t_SL g1950 ( 
.A(n_1844),
.Y(n_1950)
);

INVx6_ASAP7_75t_L g1951 ( 
.A(n_1832),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1873),
.Y(n_1952)
);

BUFx6f_ASAP7_75t_L g1953 ( 
.A(n_1873),
.Y(n_1953)
);

INVx4_ASAP7_75t_L g1954 ( 
.A(n_1853),
.Y(n_1954)
);

BUFx3_ASAP7_75t_L g1955 ( 
.A(n_1873),
.Y(n_1955)
);

INVx1_ASAP7_75t_SL g1956 ( 
.A(n_1918),
.Y(n_1956)
);

BUFx3_ASAP7_75t_L g1957 ( 
.A(n_1888),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1888),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1875),
.Y(n_1959)
);

BUFx12f_ASAP7_75t_L g1960 ( 
.A(n_1886),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1888),
.Y(n_1961)
);

BUFx3_ASAP7_75t_L g1962 ( 
.A(n_1849),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1892),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1901),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1908),
.Y(n_1965)
);

CKINVDCx6p67_ASAP7_75t_R g1966 ( 
.A(n_1887),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1853),
.Y(n_1967)
);

BUFx3_ASAP7_75t_L g1968 ( 
.A(n_1849),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1865),
.Y(n_1969)
);

INVx5_ASAP7_75t_L g1970 ( 
.A(n_1879),
.Y(n_1970)
);

BUFx24_ASAP7_75t_L g1971 ( 
.A(n_1868),
.Y(n_1971)
);

AND2x4_ASAP7_75t_L g1972 ( 
.A(n_1852),
.B(n_1858),
.Y(n_1972)
);

INVx5_ASAP7_75t_L g1973 ( 
.A(n_1879),
.Y(n_1973)
);

INVxp67_ASAP7_75t_SL g1974 ( 
.A(n_1829),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1898),
.Y(n_1975)
);

BUFx4f_ASAP7_75t_SL g1976 ( 
.A(n_1847),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1839),
.Y(n_1977)
);

INVx5_ASAP7_75t_L g1978 ( 
.A(n_1898),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1885),
.Y(n_1979)
);

OR2x2_ASAP7_75t_L g1980 ( 
.A(n_1848),
.B(n_1763),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1825),
.Y(n_1981)
);

CKINVDCx20_ASAP7_75t_R g1982 ( 
.A(n_1878),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1903),
.Y(n_1983)
);

BUFx2_ASAP7_75t_SL g1984 ( 
.A(n_1847),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1860),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1868),
.Y(n_1986)
);

INVx4_ASAP7_75t_L g1987 ( 
.A(n_1912),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1928),
.Y(n_1988)
);

A2O1A1Ixp33_ASAP7_75t_L g1989 ( 
.A1(n_1945),
.A2(n_1876),
.B(n_1914),
.C(n_1870),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1928),
.Y(n_1990)
);

AO21x2_ASAP7_75t_L g1991 ( 
.A1(n_1974),
.A2(n_1917),
.B(n_1890),
.Y(n_1991)
);

INVx1_ASAP7_75t_SL g1992 ( 
.A(n_1956),
.Y(n_1992)
);

BUFx2_ASAP7_75t_L g1993 ( 
.A(n_1954),
.Y(n_1993)
);

INVxp67_ASAP7_75t_SL g1994 ( 
.A(n_1974),
.Y(n_1994)
);

AOI21xp33_ASAP7_75t_SL g1995 ( 
.A1(n_1947),
.A2(n_1827),
.B(n_1911),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1965),
.B(n_1840),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1966),
.A2(n_1708),
.B1(n_1889),
.B2(n_1894),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1965),
.B(n_1841),
.Y(n_1998)
);

O2A1O1Ixp33_ASAP7_75t_L g1999 ( 
.A1(n_1980),
.A2(n_1893),
.B(n_1909),
.C(n_1895),
.Y(n_1999)
);

OAI21x1_ASAP7_75t_SL g2000 ( 
.A1(n_1950),
.A2(n_1915),
.B(n_1850),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1950),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1937),
.A2(n_1896),
.B(n_1867),
.Y(n_2002)
);

AOI22xp33_ASAP7_75t_L g2003 ( 
.A1(n_1966),
.A2(n_1871),
.B1(n_1861),
.B2(n_1906),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1967),
.B(n_1899),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1964),
.B(n_1838),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1959),
.B(n_1834),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1963),
.B(n_1823),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1933),
.B(n_1862),
.Y(n_2008)
);

A2O1A1Ixp33_ASAP7_75t_L g2009 ( 
.A1(n_1945),
.A2(n_1864),
.B(n_1830),
.C(n_1863),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1987),
.B(n_1859),
.Y(n_2010)
);

INVx1_ASAP7_75t_SL g2011 ( 
.A(n_1938),
.Y(n_2011)
);

BUFx3_ASAP7_75t_L g2012 ( 
.A(n_1922),
.Y(n_2012)
);

AND2x6_ASAP7_75t_L g2013 ( 
.A(n_1986),
.B(n_1790),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1936),
.B(n_1877),
.Y(n_2014)
);

OAI22xp5_ASAP7_75t_SL g2015 ( 
.A1(n_1922),
.A2(n_1891),
.B1(n_1883),
.B2(n_1711),
.Y(n_2015)
);

INVx2_ASAP7_75t_L g2016 ( 
.A(n_1941),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1935),
.A2(n_1742),
.B1(n_1755),
.B2(n_1774),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1983),
.Y(n_2018)
);

OAI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1923),
.A2(n_1762),
.B1(n_1833),
.B2(n_1777),
.Y(n_2019)
);

A2O1A1Ixp33_ASAP7_75t_L g2020 ( 
.A1(n_1971),
.A2(n_1842),
.B(n_1884),
.C(n_1869),
.Y(n_2020)
);

INVx4_ASAP7_75t_L g2021 ( 
.A(n_1951),
.Y(n_2021)
);

OAI221xp5_ASAP7_75t_L g2022 ( 
.A1(n_1937),
.A2(n_1900),
.B1(n_1754),
.B2(n_1819),
.C(n_1753),
.Y(n_2022)
);

BUFx12f_ASAP7_75t_L g2023 ( 
.A(n_1930),
.Y(n_2023)
);

CKINVDCx5p33_ASAP7_75t_R g2024 ( 
.A(n_1930),
.Y(n_2024)
);

OR2x6_ASAP7_75t_L g2025 ( 
.A(n_1937),
.B(n_1984),
.Y(n_2025)
);

OAI21x1_ASAP7_75t_L g2026 ( 
.A1(n_1977),
.A2(n_1907),
.B(n_1902),
.Y(n_2026)
);

OA21x2_ASAP7_75t_L g2027 ( 
.A1(n_1972),
.A2(n_1846),
.B(n_1836),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1920),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_1972),
.A2(n_1916),
.B(n_1768),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1949),
.Y(n_2030)
);

AO21x1_ASAP7_75t_SL g2031 ( 
.A1(n_2007),
.A2(n_1996),
.B(n_2003),
.Y(n_2031)
);

OR2x2_ASAP7_75t_L g2032 ( 
.A(n_1994),
.B(n_1921),
.Y(n_2032)
);

INVx2_ASAP7_75t_L g2033 ( 
.A(n_1988),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_2021),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1990),
.Y(n_2035)
);

BUFx3_ASAP7_75t_L g2036 ( 
.A(n_2023),
.Y(n_2036)
);

INVx6_ASAP7_75t_L g2037 ( 
.A(n_2021),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_2028),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2016),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_2001),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2007),
.Y(n_2041)
);

NAND2x1p5_ASAP7_75t_L g2042 ( 
.A(n_2027),
.B(n_1972),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1996),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2018),
.Y(n_2044)
);

AO21x2_ASAP7_75t_L g2045 ( 
.A1(n_2002),
.A2(n_1939),
.B(n_1934),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1994),
.Y(n_2046)
);

OR2x6_ASAP7_75t_L g2047 ( 
.A(n_2002),
.B(n_1971),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_2025),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_1993),
.B(n_1929),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1998),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_2014),
.B(n_1924),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2029),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_1989),
.A2(n_1923),
.B1(n_1976),
.B2(n_1982),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1998),
.B(n_2005),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2029),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_2038),
.Y(n_2056)
);

OR2x2_ASAP7_75t_L g2057 ( 
.A(n_2043),
.B(n_2006),
.Y(n_2057)
);

OA21x2_ASAP7_75t_L g2058 ( 
.A1(n_2055),
.A2(n_2052),
.B(n_2041),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2052),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_SL g2060 ( 
.A1(n_2053),
.A2(n_1997),
.B1(n_2015),
.B2(n_2013),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_2054),
.B(n_1995),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_2055),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2033),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2038),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2032),
.Y(n_2065)
);

OR2x2_ASAP7_75t_L g2066 ( 
.A(n_2043),
.B(n_2046),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2032),
.Y(n_2067)
);

HB1xp67_ASAP7_75t_L g2068 ( 
.A(n_2058),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2065),
.B(n_2048),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2058),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2067),
.B(n_2048),
.Y(n_2071)
);

AO21x2_ASAP7_75t_L g2072 ( 
.A1(n_2059),
.A2(n_2041),
.B(n_2046),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2056),
.Y(n_2073)
);

OR2x2_ASAP7_75t_L g2074 ( 
.A(n_2057),
.B(n_2066),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_2058),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2071),
.B(n_2069),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2073),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2068),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2071),
.B(n_2061),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2068),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2074),
.B(n_2061),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2075),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2072),
.B(n_2031),
.Y(n_2083)
);

AND2x2_ASAP7_75t_L g2084 ( 
.A(n_2070),
.B(n_2031),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2070),
.B(n_2034),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_2078),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2080),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2076),
.Y(n_2088)
);

AND2x2_ASAP7_75t_L g2089 ( 
.A(n_2076),
.B(n_2036),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_2084),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2083),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2082),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2081),
.B(n_2060),
.Y(n_2093)
);

INVx3_ASAP7_75t_L g2094 ( 
.A(n_2082),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2077),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2085),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_2088),
.B(n_2079),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_2094),
.A2(n_2084),
.B(n_2085),
.Y(n_2098)
);

OAI21x1_ASAP7_75t_L g2099 ( 
.A1(n_2094),
.A2(n_2075),
.B(n_2062),
.Y(n_2099)
);

AOI21x1_ASAP7_75t_L g2100 ( 
.A1(n_2090),
.A2(n_2062),
.B(n_2059),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_2094),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_2089),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2092),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2092),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2093),
.A2(n_2060),
.B(n_2009),
.Y(n_2105)
);

INVx1_ASAP7_75t_SL g2106 ( 
.A(n_2102),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2102),
.B(n_2089),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2101),
.Y(n_2108)
);

NAND3xp33_ASAP7_75t_L g2109 ( 
.A(n_2105),
.B(n_2091),
.C(n_2087),
.Y(n_2109)
);

NAND3xp33_ASAP7_75t_L g2110 ( 
.A(n_2109),
.B(n_2107),
.C(n_2108),
.Y(n_2110)
);

AOI222xp33_ASAP7_75t_L g2111 ( 
.A1(n_2106),
.A2(n_2086),
.B1(n_2097),
.B2(n_2091),
.C1(n_2095),
.C2(n_2103),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2107),
.B(n_2088),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2106),
.Y(n_2113)
);

INVxp67_ASAP7_75t_L g2114 ( 
.A(n_2112),
.Y(n_2114)
);

OR2x2_ASAP7_75t_L g2115 ( 
.A(n_2113),
.B(n_2110),
.Y(n_2115)
);

AND2x4_ASAP7_75t_SL g2116 ( 
.A(n_2111),
.B(n_1969),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2110),
.A2(n_2098),
.B(n_2097),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2113),
.B(n_2104),
.Y(n_2118)
);

AOI22xp5_ASAP7_75t_L g2119 ( 
.A1(n_2113),
.A2(n_2096),
.B1(n_2101),
.B2(n_1997),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2115),
.Y(n_2120)
);

INVx2_ASAP7_75t_SL g2121 ( 
.A(n_2116),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2118),
.Y(n_2122)
);

INVxp67_ASAP7_75t_L g2123 ( 
.A(n_2117),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2114),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_2119),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2115),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2114),
.B(n_2100),
.Y(n_2127)
);

OR2x2_ASAP7_75t_L g2128 ( 
.A(n_2115),
.B(n_2099),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_2115),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2129),
.B(n_2036),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2128),
.Y(n_2131)
);

NOR2x1_ASAP7_75t_L g2132 ( 
.A(n_2120),
.B(n_1746),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2121),
.B(n_1947),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2126),
.Y(n_2134)
);

AOI22x1_ASAP7_75t_L g2135 ( 
.A1(n_2123),
.A2(n_2024),
.B1(n_1925),
.B2(n_1926),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2125),
.B(n_2011),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2127),
.B(n_1992),
.Y(n_2137)
);

INVx1_ASAP7_75t_SL g2138 ( 
.A(n_2127),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2124),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2122),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2120),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2121),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2142),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2133),
.Y(n_2144)
);

NOR4xp25_ASAP7_75t_SL g2145 ( 
.A(n_2134),
.B(n_2030),
.C(n_2010),
.D(n_1789),
.Y(n_2145)
);

AOI322xp5_ASAP7_75t_L g2146 ( 
.A1(n_2138),
.A2(n_2003),
.A3(n_2019),
.B1(n_2017),
.B2(n_2012),
.C1(n_2020),
.C2(n_2005),
.Y(n_2146)
);

OR2x2_ASAP7_75t_L g2147 ( 
.A(n_2131),
.B(n_2072),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2141),
.B(n_2064),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2135),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2130),
.B(n_1949),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2136),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2137),
.Y(n_2152)
);

AOI21xp5_ASAP7_75t_SL g2153 ( 
.A1(n_2139),
.A2(n_1813),
.B(n_1781),
.Y(n_2153)
);

OAI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_2135),
.A2(n_1951),
.B1(n_1712),
.B2(n_1814),
.C(n_2037),
.Y(n_2154)
);

AOI211x1_ASAP7_75t_L g2155 ( 
.A1(n_2132),
.A2(n_1713),
.B(n_2019),
.C(n_2050),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2140),
.B(n_2050),
.Y(n_2156)
);

OAI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2142),
.A2(n_1923),
.B1(n_1946),
.B2(n_1942),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2144),
.Y(n_2158)
);

AOI32xp33_ASAP7_75t_L g2159 ( 
.A1(n_2143),
.A2(n_1816),
.A3(n_1812),
.B1(n_1786),
.B2(n_2034),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2151),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2157),
.A2(n_1951),
.B1(n_2037),
.B2(n_1689),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2149),
.B(n_2063),
.Y(n_2162)
);

INVxp67_ASAP7_75t_L g2163 ( 
.A(n_2150),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2152),
.A2(n_2037),
.B1(n_1689),
.B2(n_1960),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2148),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2147),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_L g2167 ( 
.A1(n_2154),
.A2(n_2156),
.B1(n_2145),
.B2(n_2153),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2155),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_2146),
.A2(n_1927),
.B(n_1919),
.Y(n_2169)
);

NAND3xp33_ASAP7_75t_L g2170 ( 
.A(n_2149),
.B(n_1699),
.C(n_1687),
.Y(n_2170)
);

INVxp33_ASAP7_75t_L g2171 ( 
.A(n_2150),
.Y(n_2171)
);

AOI222xp33_ASAP7_75t_L g2172 ( 
.A1(n_2169),
.A2(n_1742),
.B1(n_1738),
.B2(n_1803),
.C1(n_2022),
.C2(n_2017),
.Y(n_2172)
);

OR2x2_ASAP7_75t_L g2173 ( 
.A(n_2158),
.B(n_2049),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_2160),
.B(n_2034),
.Y(n_2174)
);

OAI31xp33_ASAP7_75t_SL g2175 ( 
.A1(n_2168),
.A2(n_1716),
.A3(n_2022),
.B(n_2049),
.Y(n_2175)
);

AOI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2171),
.A2(n_2170),
.B1(n_2163),
.B2(n_2165),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_2167),
.B(n_1919),
.Y(n_2177)
);

NOR2x1p5_ASAP7_75t_L g2178 ( 
.A(n_2162),
.B(n_1687),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2166),
.B(n_1927),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2164),
.Y(n_2180)
);

AOI22xp33_ASAP7_75t_L g2181 ( 
.A1(n_2161),
.A2(n_2037),
.B1(n_1960),
.B2(n_1931),
.Y(n_2181)
);

INVx1_ASAP7_75t_SL g2182 ( 
.A(n_2159),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_2158),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_2158),
.Y(n_2184)
);

AOI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2158),
.A2(n_1699),
.B1(n_1687),
.B2(n_1931),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2158),
.B(n_2051),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_2158),
.Y(n_2187)
);

INVx1_ASAP7_75t_SL g2188 ( 
.A(n_2160),
.Y(n_2188)
);

AOI22xp5_ASAP7_75t_L g2189 ( 
.A1(n_2158),
.A2(n_1699),
.B1(n_1931),
.B2(n_1982),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_2158),
.B(n_1931),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2158),
.B(n_2051),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_2158),
.B(n_1767),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2158),
.Y(n_2193)
);

AOI221x1_ASAP7_75t_L g2194 ( 
.A1(n_2184),
.A2(n_1766),
.B1(n_1769),
.B2(n_1737),
.C(n_1760),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2188),
.B(n_139),
.Y(n_2195)
);

NOR2x1_ASAP7_75t_L g2196 ( 
.A(n_2183),
.B(n_1750),
.Y(n_2196)
);

AND3x2_ASAP7_75t_L g2197 ( 
.A(n_2187),
.B(n_139),
.C(n_140),
.Y(n_2197)
);

OAI211xp5_ASAP7_75t_SL g2198 ( 
.A1(n_2176),
.A2(n_1780),
.B(n_1779),
.C(n_1806),
.Y(n_2198)
);

OAI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2177),
.A2(n_1809),
.B(n_1821),
.C(n_1808),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_2193),
.B(n_141),
.C(n_142),
.Y(n_2200)
);

NOR3x1_ASAP7_75t_L g2201 ( 
.A(n_2174),
.B(n_1905),
.C(n_141),
.Y(n_2201)
);

AOI211x1_ASAP7_75t_L g2202 ( 
.A1(n_2190),
.A2(n_1897),
.B(n_1882),
.C(n_2044),
.Y(n_2202)
);

NAND4xp25_ASAP7_75t_L g2203 ( 
.A(n_2180),
.B(n_1999),
.C(n_1981),
.D(n_1820),
.Y(n_2203)
);

AND3x2_ASAP7_75t_L g2204 ( 
.A(n_2192),
.B(n_142),
.C(n_143),
.Y(n_2204)
);

NOR2xp67_ASAP7_75t_L g2205 ( 
.A(n_2173),
.B(n_143),
.Y(n_2205)
);

AOI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_2188),
.A2(n_1999),
.B1(n_1910),
.B2(n_2000),
.C(n_146),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2186),
.B(n_144),
.Y(n_2207)
);

NAND4xp25_ASAP7_75t_L g2208 ( 
.A(n_2182),
.B(n_1981),
.C(n_1714),
.D(n_1987),
.Y(n_2208)
);

NAND4xp25_ASAP7_75t_L g2209 ( 
.A(n_2181),
.B(n_146),
.C(n_144),
.D(n_145),
.Y(n_2209)
);

NAND2x1_ASAP7_75t_L g2210 ( 
.A(n_2191),
.B(n_2047),
.Y(n_2210)
);

NAND3xp33_ASAP7_75t_L g2211 ( 
.A(n_2179),
.B(n_145),
.C(n_147),
.Y(n_2211)
);

NAND4xp25_ASAP7_75t_L g2212 ( 
.A(n_2172),
.B(n_149),
.C(n_147),
.D(n_148),
.Y(n_2212)
);

AOI21xp5_ASAP7_75t_L g2213 ( 
.A1(n_2175),
.A2(n_2189),
.B(n_2185),
.Y(n_2213)
);

NOR5xp2_ASAP7_75t_L g2214 ( 
.A(n_2178),
.B(n_150),
.C(n_148),
.D(n_149),
.E(n_151),
.Y(n_2214)
);

INVxp67_ASAP7_75t_SL g2215 ( 
.A(n_2174),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_SL g2216 ( 
.A(n_2188),
.B(n_1985),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2188),
.B(n_1985),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2173),
.Y(n_2218)
);

XOR2xp5_ASAP7_75t_L g2219 ( 
.A(n_2183),
.B(n_150),
.Y(n_2219)
);

NOR3xp33_ASAP7_75t_L g2220 ( 
.A(n_2180),
.B(n_151),
.C(n_154),
.Y(n_2220)
);

NOR3x1_ASAP7_75t_L g2221 ( 
.A(n_2177),
.B(n_154),
.C(n_155),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2188),
.B(n_1985),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_SL g2223 ( 
.A(n_2188),
.B(n_1976),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2188),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_SL g2225 ( 
.A(n_2188),
.B(n_1985),
.Y(n_2225)
);

NAND3xp33_ASAP7_75t_L g2226 ( 
.A(n_2176),
.B(n_155),
.C(n_156),
.Y(n_2226)
);

NOR2xp67_ASAP7_75t_L g2227 ( 
.A(n_2187),
.B(n_156),
.Y(n_2227)
);

AOI211xp5_ASAP7_75t_L g2228 ( 
.A1(n_2188),
.A2(n_159),
.B(n_157),
.C(n_158),
.Y(n_2228)
);

NAND3xp33_ASAP7_75t_L g2229 ( 
.A(n_2176),
.B(n_157),
.C(n_158),
.Y(n_2229)
);

CKINVDCx5p33_ASAP7_75t_R g2230 ( 
.A(n_2183),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_2197),
.Y(n_2231)
);

OAI211xp5_ASAP7_75t_L g2232 ( 
.A1(n_2209),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_2232)
);

OAI211xp5_ASAP7_75t_L g2233 ( 
.A1(n_2205),
.A2(n_2195),
.B(n_2224),
.C(n_2220),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_2230),
.B(n_161),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2208),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.C(n_165),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2223),
.A2(n_2047),
.B1(n_2042),
.B2(n_2025),
.C(n_1851),
.Y(n_2236)
);

NAND3xp33_ASAP7_75t_L g2237 ( 
.A(n_2226),
.B(n_165),
.C(n_166),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2204),
.B(n_166),
.Y(n_2238)
);

NOR3xp33_ASAP7_75t_L g2239 ( 
.A(n_2218),
.B(n_167),
.C(n_168),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_2207),
.B(n_167),
.Y(n_2240)
);

NAND2x2_ASAP7_75t_L g2241 ( 
.A(n_2212),
.B(n_168),
.Y(n_2241)
);

OA22x2_ASAP7_75t_L g2242 ( 
.A1(n_2216),
.A2(n_2047),
.B1(n_2040),
.B2(n_2025),
.Y(n_2242)
);

NOR3x1_ASAP7_75t_L g2243 ( 
.A(n_2229),
.B(n_170),
.C(n_171),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2219),
.Y(n_2244)
);

NAND4xp25_ASAP7_75t_L g2245 ( 
.A(n_2221),
.B(n_173),
.C(n_170),
.D(n_172),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_2211),
.B(n_172),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2228),
.B(n_174),
.C(n_175),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2227),
.Y(n_2248)
);

NOR2xp67_ASAP7_75t_L g2249 ( 
.A(n_2200),
.B(n_174),
.Y(n_2249)
);

NOR2xp33_ASAP7_75t_L g2250 ( 
.A(n_2225),
.B(n_175),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2217),
.B(n_176),
.Y(n_2251)
);

NAND3xp33_ASAP7_75t_SL g2252 ( 
.A(n_2214),
.B(n_176),
.C(n_177),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2210),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2222),
.B(n_177),
.Y(n_2254)
);

OAI221xp5_ASAP7_75t_L g2255 ( 
.A1(n_2206),
.A2(n_2047),
.B1(n_2042),
.B2(n_180),
.C(n_178),
.Y(n_2255)
);

O2A1O1Ixp5_ASAP7_75t_L g2256 ( 
.A1(n_2213),
.A2(n_180),
.B(n_178),
.C(n_179),
.Y(n_2256)
);

INVx1_ASAP7_75t_SL g2257 ( 
.A(n_2196),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_2215),
.B(n_2042),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2201),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2194),
.Y(n_2260)
);

AOI211xp5_ASAP7_75t_SL g2261 ( 
.A1(n_2199),
.A2(n_182),
.B(n_179),
.C(n_181),
.Y(n_2261)
);

INVx2_ASAP7_75t_L g2262 ( 
.A(n_2202),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2203),
.B(n_2040),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2198),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2224),
.B(n_2004),
.Y(n_2265)
);

NAND3xp33_ASAP7_75t_L g2266 ( 
.A(n_2220),
.B(n_181),
.C(n_182),
.Y(n_2266)
);

NAND3xp33_ASAP7_75t_SL g2267 ( 
.A(n_2224),
.B(n_183),
.C(n_184),
.Y(n_2267)
);

AOI211x1_ASAP7_75t_L g2268 ( 
.A1(n_2216),
.A2(n_2035),
.B(n_185),
.C(n_183),
.Y(n_2268)
);

AOI211xp5_ASAP7_75t_SL g2269 ( 
.A1(n_2233),
.A2(n_186),
.B(n_184),
.C(n_185),
.Y(n_2269)
);

A2O1A1Ixp33_ASAP7_75t_SL g2270 ( 
.A1(n_2244),
.A2(n_189),
.B(n_187),
.C(n_188),
.Y(n_2270)
);

AOI32xp33_ASAP7_75t_L g2271 ( 
.A1(n_2231),
.A2(n_1716),
.A3(n_1948),
.B1(n_1957),
.B2(n_1955),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2234),
.B(n_188),
.Y(n_2272)
);

AOI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_2265),
.A2(n_2013),
.B1(n_1952),
.B2(n_1953),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2252),
.A2(n_2013),
.B1(n_1952),
.B2(n_1953),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_2238),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2231),
.Y(n_2276)
);

AOI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2267),
.A2(n_2013),
.B1(n_1952),
.B2(n_1953),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2241),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2256),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_2243),
.Y(n_2280)
);

AOI321xp33_ASAP7_75t_L g2281 ( 
.A1(n_2253),
.A2(n_1716),
.A3(n_192),
.B1(n_194),
.B2(n_190),
.C(n_191),
.Y(n_2281)
);

AOI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2232),
.A2(n_2240),
.B1(n_2246),
.B2(n_2245),
.Y(n_2282)
);

CKINVDCx5p33_ASAP7_75t_R g2283 ( 
.A(n_2248),
.Y(n_2283)
);

AOI21xp5_ASAP7_75t_SL g2284 ( 
.A1(n_2260),
.A2(n_190),
.B(n_191),
.Y(n_2284)
);

INVx1_ASAP7_75t_SL g2285 ( 
.A(n_2257),
.Y(n_2285)
);

AOI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_2259),
.A2(n_2255),
.B1(n_2249),
.B2(n_2251),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2266),
.Y(n_2287)
);

NOR3xp33_ASAP7_75t_L g2288 ( 
.A(n_2237),
.B(n_192),
.C(n_193),
.Y(n_2288)
);

NAND3xp33_ASAP7_75t_L g2289 ( 
.A(n_2250),
.B(n_193),
.C(n_194),
.Y(n_2289)
);

NOR2x1_ASAP7_75t_L g2290 ( 
.A(n_2247),
.B(n_195),
.Y(n_2290)
);

AOI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2254),
.A2(n_2013),
.B1(n_1952),
.B2(n_1953),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2268),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2239),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_SL g2294 ( 
.A(n_2264),
.B(n_195),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2262),
.Y(n_2295)
);

NOR2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2261),
.B(n_2263),
.Y(n_2296)
);

XOR2xp5_ASAP7_75t_L g2297 ( 
.A(n_2258),
.B(n_196),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2235),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2242),
.B(n_196),
.Y(n_2299)
);

OAI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2236),
.A2(n_1932),
.B1(n_1955),
.B2(n_1948),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_2234),
.B(n_197),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2238),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_L g2303 ( 
.A1(n_2252),
.A2(n_1957),
.B1(n_1932),
.B2(n_1944),
.Y(n_2303)
);

OAI211xp5_ASAP7_75t_L g2304 ( 
.A1(n_2232),
.A2(n_200),
.B(n_198),
.C(n_199),
.Y(n_2304)
);

AOI322xp5_ASAP7_75t_L g2305 ( 
.A1(n_2252),
.A2(n_2008),
.A3(n_2035),
.B1(n_1944),
.B2(n_1958),
.C1(n_1961),
.C2(n_2039),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2234),
.B(n_199),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_2252),
.A2(n_1932),
.B1(n_1961),
.B2(n_1958),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2238),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_2245),
.B(n_200),
.Y(n_2309)
);

NAND2xp33_ASAP7_75t_L g2310 ( 
.A(n_2239),
.B(n_1932),
.Y(n_2310)
);

INVxp67_ASAP7_75t_L g2311 ( 
.A(n_2234),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2231),
.Y(n_2312)
);

OR2x6_ASAP7_75t_L g2313 ( 
.A(n_2248),
.B(n_201),
.Y(n_2313)
);

AOI21xp33_ASAP7_75t_L g2314 ( 
.A1(n_2253),
.A2(n_202),
.B(n_203),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2238),
.Y(n_2315)
);

AOI211x1_ASAP7_75t_L g2316 ( 
.A1(n_2255),
.A2(n_206),
.B(n_204),
.C(n_205),
.Y(n_2316)
);

O2A1O1Ixp33_ASAP7_75t_L g2317 ( 
.A1(n_2267),
.A2(n_208),
.B(n_205),
.C(n_207),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2238),
.Y(n_2318)
);

INVx1_ASAP7_75t_SL g2319 ( 
.A(n_2238),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_2234),
.B(n_208),
.Y(n_2320)
);

A2O1A1Ixp33_ASAP7_75t_L g2321 ( 
.A1(n_2256),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_2321)
);

AOI22xp5_ASAP7_75t_L g2322 ( 
.A1(n_2234),
.A2(n_2008),
.B1(n_2045),
.B2(n_1954),
.Y(n_2322)
);

XNOR2x1_ASAP7_75t_L g2323 ( 
.A(n_2244),
.B(n_209),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2238),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2238),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2238),
.Y(n_2326)
);

AOI22xp33_ASAP7_75t_L g2327 ( 
.A1(n_2252),
.A2(n_2045),
.B1(n_1968),
.B2(n_1975),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2265),
.B(n_1940),
.Y(n_2328)
);

OAI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2256),
.A2(n_1723),
.B(n_2026),
.Y(n_2329)
);

AOI221x1_ASAP7_75t_SL g2330 ( 
.A1(n_2249),
.A2(n_213),
.B1(n_211),
.B2(n_212),
.C(n_214),
.Y(n_2330)
);

AOI22xp33_ASAP7_75t_L g2331 ( 
.A1(n_2312),
.A2(n_2045),
.B1(n_1968),
.B2(n_1975),
.Y(n_2331)
);

NOR4xp25_ASAP7_75t_L g2332 ( 
.A(n_2285),
.B(n_2276),
.C(n_2279),
.D(n_2295),
.Y(n_2332)
);

AOI22xp5_ASAP7_75t_L g2333 ( 
.A1(n_2274),
.A2(n_1940),
.B1(n_1943),
.B2(n_2039),
.Y(n_2333)
);

OR2x2_ASAP7_75t_L g2334 ( 
.A(n_2299),
.B(n_213),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2323),
.Y(n_2335)
);

NOR4xp25_ASAP7_75t_L g2336 ( 
.A(n_2319),
.B(n_2278),
.C(n_2304),
.D(n_2287),
.Y(n_2336)
);

AOI22xp5_ASAP7_75t_L g2337 ( 
.A1(n_2309),
.A2(n_1943),
.B1(n_1962),
.B2(n_2033),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2313),
.Y(n_2338)
);

NOR2x1_ASAP7_75t_L g2339 ( 
.A(n_2284),
.B(n_2313),
.Y(n_2339)
);

NOR2x1_ASAP7_75t_L g2340 ( 
.A(n_2313),
.B(n_215),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_2292),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2297),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2269),
.B(n_215),
.Y(n_2343)
);

NOR4xp25_ASAP7_75t_L g2344 ( 
.A(n_2293),
.B(n_218),
.C(n_216),
.D(n_217),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2330),
.B(n_216),
.Y(n_2345)
);

AOI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_2294),
.A2(n_1962),
.B1(n_1986),
.B2(n_2027),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2317),
.Y(n_2347)
);

AOI221xp5_ASAP7_75t_SL g2348 ( 
.A1(n_2310),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.C(n_223),
.Y(n_2348)
);

OAI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2303),
.A2(n_1970),
.B1(n_1978),
.B2(n_1973),
.Y(n_2349)
);

OAI22xp5_ASAP7_75t_SL g2350 ( 
.A1(n_2316),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2272),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2301),
.Y(n_2352)
);

NOR2x1_ASAP7_75t_L g2353 ( 
.A(n_2289),
.B(n_224),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2306),
.Y(n_2354)
);

AO22x1_ASAP7_75t_L g2355 ( 
.A1(n_2290),
.A2(n_227),
.B1(n_224),
.B2(n_225),
.Y(n_2355)
);

AOI221xp5_ASAP7_75t_L g2356 ( 
.A1(n_2300),
.A2(n_229),
.B1(n_225),
.B2(n_228),
.C(n_231),
.Y(n_2356)
);

AOI221xp5_ASAP7_75t_L g2357 ( 
.A1(n_2327),
.A2(n_232),
.B1(n_228),
.B2(n_231),
.C(n_233),
.Y(n_2357)
);

NOR2x1_ASAP7_75t_L g2358 ( 
.A(n_2320),
.B(n_232),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2305),
.B(n_233),
.Y(n_2359)
);

AOI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2283),
.A2(n_1986),
.B1(n_2006),
.B2(n_1991),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2321),
.Y(n_2361)
);

NOR2x1_ASAP7_75t_L g2362 ( 
.A(n_2280),
.B(n_234),
.Y(n_2362)
);

OA22x2_ASAP7_75t_L g2363 ( 
.A1(n_2277),
.A2(n_237),
.B1(n_234),
.B2(n_236),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2288),
.B(n_237),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2296),
.Y(n_2365)
);

AOI31xp33_ASAP7_75t_L g2366 ( 
.A1(n_2275),
.A2(n_242),
.A3(n_239),
.B(n_240),
.Y(n_2366)
);

NOR2x1_ASAP7_75t_L g2367 ( 
.A(n_2302),
.B(n_239),
.Y(n_2367)
);

NOR4xp25_ASAP7_75t_L g2368 ( 
.A(n_2298),
.B(n_244),
.C(n_242),
.D(n_243),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_SL g2369 ( 
.A(n_2286),
.B(n_245),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2308),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2315),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2307),
.A2(n_1970),
.B1(n_1978),
.B2(n_1973),
.Y(n_2372)
);

NOR2x1_ASAP7_75t_L g2373 ( 
.A(n_2318),
.B(n_245),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2324),
.Y(n_2374)
);

AOI22xp5_ASAP7_75t_L g2375 ( 
.A1(n_2325),
.A2(n_1986),
.B1(n_1991),
.B2(n_1970),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_2282),
.B(n_246),
.Y(n_2376)
);

INVx3_ASAP7_75t_L g2377 ( 
.A(n_2326),
.Y(n_2377)
);

NOR4xp25_ASAP7_75t_L g2378 ( 
.A(n_2311),
.B(n_248),
.C(n_246),
.D(n_247),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2328),
.Y(n_2379)
);

NOR2x1_ASAP7_75t_L g2380 ( 
.A(n_2270),
.B(n_247),
.Y(n_2380)
);

AOI221xp5_ASAP7_75t_L g2381 ( 
.A1(n_2314),
.A2(n_2271),
.B1(n_2329),
.B2(n_2291),
.C(n_2273),
.Y(n_2381)
);

NOR2x1_ASAP7_75t_L g2382 ( 
.A(n_2281),
.B(n_248),
.Y(n_2382)
);

A2O1A1Ixp33_ASAP7_75t_SL g2383 ( 
.A1(n_2322),
.A2(n_251),
.B(n_249),
.C(n_250),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_2274),
.B(n_249),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2269),
.B(n_251),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_2269),
.B(n_252),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_SL g2387 ( 
.A(n_2274),
.B(n_252),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2323),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2323),
.Y(n_2389)
);

OR2x2_ASAP7_75t_L g2390 ( 
.A(n_2299),
.B(n_254),
.Y(n_2390)
);

NOR2x1_ASAP7_75t_L g2391 ( 
.A(n_2284),
.B(n_254),
.Y(n_2391)
);

OAI22x1_ASAP7_75t_L g2392 ( 
.A1(n_2297),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2269),
.B(n_256),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2323),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2323),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_2285),
.A2(n_1970),
.B1(n_1978),
.B2(n_1973),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2313),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2341),
.B(n_257),
.Y(n_2398)
);

AO22x1_ASAP7_75t_L g2399 ( 
.A1(n_2339),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_SL g2400 ( 
.A(n_2378),
.B(n_261),
.Y(n_2400)
);

NOR2x1_ASAP7_75t_L g2401 ( 
.A(n_2340),
.B(n_261),
.Y(n_2401)
);

NAND3xp33_ASAP7_75t_L g2402 ( 
.A(n_2391),
.B(n_262),
.C(n_263),
.Y(n_2402)
);

BUFx12f_ASAP7_75t_L g2403 ( 
.A(n_2334),
.Y(n_2403)
);

NAND2xp5_ASAP7_75t_L g2404 ( 
.A(n_2355),
.B(n_2344),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2397),
.B(n_262),
.Y(n_2405)
);

OAI221xp5_ASAP7_75t_L g2406 ( 
.A1(n_2332),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C(n_267),
.Y(n_2406)
);

NOR3xp33_ASAP7_75t_L g2407 ( 
.A(n_2397),
.B(n_266),
.C(n_267),
.Y(n_2407)
);

NAND3xp33_ASAP7_75t_L g2408 ( 
.A(n_2356),
.B(n_268),
.C(n_269),
.Y(n_2408)
);

NAND4xp25_ASAP7_75t_L g2409 ( 
.A(n_2357),
.B(n_271),
.C(n_269),
.D(n_270),
.Y(n_2409)
);

OAI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2348),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.C(n_273),
.Y(n_2410)
);

NOR2x1_ASAP7_75t_L g2411 ( 
.A(n_2362),
.B(n_272),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2368),
.B(n_273),
.Y(n_2412)
);

NAND3xp33_ASAP7_75t_L g2413 ( 
.A(n_2367),
.B(n_274),
.C(n_275),
.Y(n_2413)
);

NAND3xp33_ASAP7_75t_L g2414 ( 
.A(n_2373),
.B(n_274),
.C(n_275),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2350),
.Y(n_2415)
);

NOR3xp33_ASAP7_75t_L g2416 ( 
.A(n_2365),
.B(n_276),
.C(n_277),
.Y(n_2416)
);

INVx3_ASAP7_75t_L g2417 ( 
.A(n_2338),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2396),
.A2(n_1973),
.B1(n_1978),
.B2(n_1815),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_SL g2419 ( 
.A(n_2380),
.B(n_276),
.Y(n_2419)
);

NOR2x1_ASAP7_75t_L g2420 ( 
.A(n_2358),
.B(n_277),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_2392),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2343),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2385),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2386),
.Y(n_2424)
);

NOR3xp33_ASAP7_75t_L g2425 ( 
.A(n_2377),
.B(n_278),
.C(n_279),
.Y(n_2425)
);

NOR2x1_ASAP7_75t_L g2426 ( 
.A(n_2366),
.B(n_278),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2382),
.B(n_279),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_L g2428 ( 
.A(n_2393),
.B(n_280),
.Y(n_2428)
);

NOR3xp33_ASAP7_75t_SL g2429 ( 
.A(n_2345),
.B(n_280),
.C(n_281),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2363),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_SL g2431 ( 
.A(n_2336),
.B(n_281),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2337),
.A2(n_1979),
.B1(n_1983),
.B2(n_284),
.Y(n_2432)
);

NAND2xp33_ASAP7_75t_L g2433 ( 
.A(n_2353),
.B(n_282),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2390),
.B(n_283),
.Y(n_2434)
);

INVxp67_ASAP7_75t_SL g2435 ( 
.A(n_2376),
.Y(n_2435)
);

NOR2x1_ASAP7_75t_L g2436 ( 
.A(n_2369),
.B(n_284),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2379),
.B(n_285),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2377),
.B(n_285),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2359),
.Y(n_2439)
);

NOR4xp75_ASAP7_75t_L g2440 ( 
.A(n_2364),
.B(n_288),
.C(n_286),
.D(n_287),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2383),
.B(n_2361),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2347),
.B(n_286),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2384),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2370),
.B(n_287),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2371),
.B(n_288),
.Y(n_2445)
);

OAI22xp33_ASAP7_75t_SL g2446 ( 
.A1(n_2387),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2374),
.Y(n_2447)
);

NAND3x1_ASAP7_75t_SL g2448 ( 
.A(n_2381),
.B(n_290),
.C(n_292),
.Y(n_2448)
);

NAND3xp33_ASAP7_75t_L g2449 ( 
.A(n_2335),
.B(n_293),
.C(n_295),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2388),
.B(n_293),
.Y(n_2450)
);

AOI21xp5_ASAP7_75t_L g2451 ( 
.A1(n_2389),
.A2(n_295),
.B(n_296),
.Y(n_2451)
);

AND3x1_ASAP7_75t_L g2452 ( 
.A(n_2395),
.B(n_296),
.C(n_297),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2394),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2342),
.B(n_297),
.Y(n_2454)
);

XNOR2xp5_ASAP7_75t_L g2455 ( 
.A(n_2351),
.B(n_298),
.Y(n_2455)
);

NAND3xp33_ASAP7_75t_L g2456 ( 
.A(n_2352),
.B(n_298),
.C(n_299),
.Y(n_2456)
);

AND3x1_ASAP7_75t_L g2457 ( 
.A(n_2354),
.B(n_299),
.C(n_300),
.Y(n_2457)
);

NOR2xp33_ASAP7_75t_L g2458 ( 
.A(n_2333),
.B(n_300),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2346),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2349),
.A2(n_301),
.B1(n_302),
.B2(n_303),
.Y(n_2460)
);

OAI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2331),
.A2(n_303),
.B(n_304),
.Y(n_2461)
);

NOR4xp25_ASAP7_75t_L g2462 ( 
.A(n_2431),
.B(n_2372),
.C(n_2360),
.D(n_306),
.Y(n_2462)
);

NOR3xp33_ASAP7_75t_L g2463 ( 
.A(n_2417),
.B(n_2375),
.C(n_304),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2401),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2405),
.Y(n_2465)
);

NAND3xp33_ASAP7_75t_SL g2466 ( 
.A(n_2406),
.B(n_305),
.C(n_306),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2438),
.Y(n_2467)
);

NAND4xp25_ASAP7_75t_L g2468 ( 
.A(n_2428),
.B(n_307),
.C(n_308),
.D(n_309),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_L g2469 ( 
.A(n_2399),
.B(n_307),
.Y(n_2469)
);

XNOR2x1_ASAP7_75t_L g2470 ( 
.A(n_2426),
.B(n_308),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2407),
.B(n_309),
.Y(n_2471)
);

NOR2x1p5_ASAP7_75t_L g2472 ( 
.A(n_2412),
.B(n_310),
.Y(n_2472)
);

AND3x2_ASAP7_75t_L g2473 ( 
.A(n_2415),
.B(n_310),
.C(n_311),
.Y(n_2473)
);

NOR3xp33_ASAP7_75t_L g2474 ( 
.A(n_2417),
.B(n_311),
.C(n_312),
.Y(n_2474)
);

NAND4xp25_ASAP7_75t_L g2475 ( 
.A(n_2402),
.B(n_312),
.C(n_314),
.D(n_315),
.Y(n_2475)
);

NAND3xp33_ASAP7_75t_SL g2476 ( 
.A(n_2421),
.B(n_314),
.C(n_315),
.Y(n_2476)
);

NAND4xp25_ASAP7_75t_L g2477 ( 
.A(n_2409),
.B(n_316),
.C(n_317),
.D(n_318),
.Y(n_2477)
);

NAND4xp25_ASAP7_75t_L g2478 ( 
.A(n_2427),
.B(n_2408),
.C(n_2441),
.D(n_2410),
.Y(n_2478)
);

AND2x4_ASAP7_75t_L g2479 ( 
.A(n_2430),
.B(n_316),
.Y(n_2479)
);

OR2x2_ASAP7_75t_L g2480 ( 
.A(n_2434),
.B(n_317),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2442),
.B(n_318),
.Y(n_2481)
);

AND3x2_ASAP7_75t_L g2482 ( 
.A(n_2425),
.B(n_319),
.C(n_320),
.Y(n_2482)
);

OR2x2_ASAP7_75t_L g2483 ( 
.A(n_2404),
.B(n_320),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2452),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2419),
.B(n_321),
.Y(n_2485)
);

OR2x2_ASAP7_75t_L g2486 ( 
.A(n_2400),
.B(n_321),
.Y(n_2486)
);

NAND3x1_ASAP7_75t_L g2487 ( 
.A(n_2411),
.B(n_322),
.C(n_323),
.Y(n_2487)
);

NOR2x1_ASAP7_75t_L g2488 ( 
.A(n_2420),
.B(n_322),
.Y(n_2488)
);

INVxp67_ASAP7_75t_L g2489 ( 
.A(n_2457),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_SL g2490 ( 
.A(n_2440),
.B(n_323),
.C(n_324),
.Y(n_2490)
);

NOR2x1_ASAP7_75t_L g2491 ( 
.A(n_2413),
.B(n_324),
.Y(n_2491)
);

OR2x2_ASAP7_75t_L g2492 ( 
.A(n_2414),
.B(n_325),
.Y(n_2492)
);

NOR3xp33_ASAP7_75t_L g2493 ( 
.A(n_2447),
.B(n_326),
.C(n_327),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2416),
.B(n_2451),
.Y(n_2494)
);

NAND4xp25_ASAP7_75t_L g2495 ( 
.A(n_2453),
.B(n_327),
.C(n_328),
.D(n_329),
.Y(n_2495)
);

NOR3xp33_ASAP7_75t_L g2496 ( 
.A(n_2435),
.B(n_329),
.C(n_330),
.Y(n_2496)
);

NOR2x1_ASAP7_75t_L g2497 ( 
.A(n_2456),
.B(n_330),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2444),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2398),
.B(n_331),
.Y(n_2499)
);

OAI211xp5_ASAP7_75t_L g2500 ( 
.A1(n_2460),
.A2(n_331),
.B(n_332),
.C(n_333),
.Y(n_2500)
);

NAND5xp2_ASAP7_75t_L g2501 ( 
.A(n_2439),
.B(n_2458),
.C(n_2461),
.D(n_2443),
.E(n_2424),
.Y(n_2501)
);

AO211x2_ASAP7_75t_L g2502 ( 
.A1(n_2459),
.A2(n_332),
.B(n_333),
.C(n_334),
.Y(n_2502)
);

NAND3xp33_ASAP7_75t_SL g2503 ( 
.A(n_2429),
.B(n_334),
.C(n_335),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_L g2504 ( 
.A(n_2448),
.B(n_336),
.C(n_337),
.Y(n_2504)
);

OR2x2_ASAP7_75t_L g2505 ( 
.A(n_2449),
.B(n_336),
.Y(n_2505)
);

NAND3xp33_ASAP7_75t_SL g2506 ( 
.A(n_2483),
.B(n_2422),
.C(n_2423),
.Y(n_2506)
);

OAI211xp5_ASAP7_75t_L g2507 ( 
.A1(n_2469),
.A2(n_2436),
.B(n_2445),
.C(n_2450),
.Y(n_2507)
);

NAND4xp75_ASAP7_75t_L g2508 ( 
.A(n_2488),
.B(n_2437),
.C(n_2454),
.D(n_2403),
.Y(n_2508)
);

AOI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2462),
.A2(n_2446),
.B1(n_2433),
.B2(n_2432),
.C(n_2418),
.Y(n_2509)
);

OAI221xp5_ASAP7_75t_SL g2510 ( 
.A1(n_2486),
.A2(n_2504),
.B1(n_2485),
.B2(n_2492),
.C(n_2489),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2479),
.B(n_2455),
.Y(n_2511)
);

NOR3xp33_ASAP7_75t_SL g2512 ( 
.A(n_2478),
.B(n_337),
.C(n_338),
.Y(n_2512)
);

NAND5xp2_ASAP7_75t_L g2513 ( 
.A(n_2484),
.B(n_338),
.C(n_339),
.D(n_340),
.E(n_341),
.Y(n_2513)
);

HB1xp67_ASAP7_75t_L g2514 ( 
.A(n_2502),
.Y(n_2514)
);

AOI21xp5_ASAP7_75t_SL g2515 ( 
.A1(n_2470),
.A2(n_340),
.B(n_341),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2473),
.Y(n_2516)
);

NOR2x1_ASAP7_75t_L g2517 ( 
.A(n_2476),
.B(n_342),
.Y(n_2517)
);

NOR4xp25_ASAP7_75t_L g2518 ( 
.A(n_2487),
.B(n_344),
.C(n_345),
.D(n_346),
.Y(n_2518)
);

NAND4xp75_ASAP7_75t_L g2519 ( 
.A(n_2491),
.B(n_344),
.C(n_345),
.D(n_347),
.Y(n_2519)
);

CKINVDCx16_ASAP7_75t_R g2520 ( 
.A(n_2503),
.Y(n_2520)
);

NAND5xp2_ASAP7_75t_L g2521 ( 
.A(n_2463),
.B(n_347),
.C(n_348),
.D(n_349),
.E(n_350),
.Y(n_2521)
);

NAND4xp75_ASAP7_75t_L g2522 ( 
.A(n_2497),
.B(n_348),
.C(n_349),
.D(n_351),
.Y(n_2522)
);

AOI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2466),
.A2(n_351),
.B1(n_352),
.B2(n_353),
.C(n_354),
.Y(n_2523)
);

NOR2xp67_ASAP7_75t_L g2524 ( 
.A(n_2490),
.B(n_2468),
.Y(n_2524)
);

OR2x2_ASAP7_75t_L g2525 ( 
.A(n_2475),
.B(n_352),
.Y(n_2525)
);

AND2x4_ASAP7_75t_L g2526 ( 
.A(n_2472),
.B(n_353),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2480),
.Y(n_2527)
);

AOI211x1_ASAP7_75t_L g2528 ( 
.A1(n_2500),
.A2(n_354),
.B(n_355),
.C(n_356),
.Y(n_2528)
);

OAI21xp33_ASAP7_75t_L g2529 ( 
.A1(n_2501),
.A2(n_2477),
.B(n_2471),
.Y(n_2529)
);

OAI211xp5_ASAP7_75t_SL g2530 ( 
.A1(n_2494),
.A2(n_356),
.B(n_357),
.C(n_359),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2499),
.B(n_357),
.Y(n_2531)
);

NOR2x1p5_ASAP7_75t_L g2532 ( 
.A(n_2505),
.B(n_360),
.Y(n_2532)
);

OAI22x1_ASAP7_75t_L g2533 ( 
.A1(n_2464),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.Y(n_2533)
);

OR5x1_ASAP7_75t_L g2534 ( 
.A(n_2495),
.B(n_361),
.C(n_362),
.D(n_363),
.E(n_364),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2482),
.Y(n_2535)
);

NAND5xp2_ASAP7_75t_L g2536 ( 
.A(n_2465),
.B(n_363),
.C(n_364),
.D(n_365),
.E(n_366),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2481),
.Y(n_2537)
);

NOR3x1_ASAP7_75t_L g2538 ( 
.A(n_2467),
.B(n_365),
.C(n_367),
.Y(n_2538)
);

NAND3xp33_ASAP7_75t_SL g2539 ( 
.A(n_2496),
.B(n_368),
.C(n_369),
.Y(n_2539)
);

CKINVDCx16_ASAP7_75t_R g2540 ( 
.A(n_2498),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2493),
.Y(n_2541)
);

AOI22xp5_ASAP7_75t_L g2542 ( 
.A1(n_2524),
.A2(n_2474),
.B1(n_370),
.B2(n_371),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_2526),
.B(n_369),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2526),
.B(n_2518),
.Y(n_2544)
);

AND2x4_ASAP7_75t_L g2545 ( 
.A(n_2532),
.B(n_371),
.Y(n_2545)
);

INVx3_ASAP7_75t_L g2546 ( 
.A(n_2516),
.Y(n_2546)
);

NAND2xp33_ASAP7_75t_SL g2547 ( 
.A(n_2512),
.B(n_372),
.Y(n_2547)
);

NOR2xp67_ASAP7_75t_SL g2548 ( 
.A(n_2508),
.B(n_2537),
.Y(n_2548)
);

NAND4xp75_ASAP7_75t_L g2549 ( 
.A(n_2535),
.B(n_372),
.C(n_373),
.D(n_374),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2519),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2527),
.B(n_373),
.Y(n_2551)
);

AND2x4_ASAP7_75t_L g2552 ( 
.A(n_2517),
.B(n_374),
.Y(n_2552)
);

AND2x2_ASAP7_75t_L g2553 ( 
.A(n_2514),
.B(n_375),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2522),
.Y(n_2554)
);

AND2x4_ASAP7_75t_L g2555 ( 
.A(n_2541),
.B(n_375),
.Y(n_2555)
);

AND2x4_ASAP7_75t_L g2556 ( 
.A(n_2538),
.B(n_376),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2511),
.B(n_376),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2531),
.Y(n_2558)
);

AND3x4_ASAP7_75t_L g2559 ( 
.A(n_2534),
.B(n_377),
.C(n_378),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_2533),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2528),
.Y(n_2561)
);

NAND2xp5_ASAP7_75t_L g2562 ( 
.A(n_2523),
.B(n_377),
.Y(n_2562)
);

NAND4xp25_ASAP7_75t_L g2563 ( 
.A(n_2521),
.B(n_2509),
.C(n_2510),
.D(n_2529),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2525),
.Y(n_2564)
);

AND2x2_ASAP7_75t_L g2565 ( 
.A(n_2520),
.B(n_378),
.Y(n_2565)
);

AOI21xp5_ASAP7_75t_L g2566 ( 
.A1(n_2544),
.A2(n_2547),
.B(n_2515),
.Y(n_2566)
);

HB1xp67_ASAP7_75t_L g2567 ( 
.A(n_2549),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2565),
.Y(n_2568)
);

OAI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2542),
.A2(n_2540),
.B1(n_2507),
.B2(n_2530),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2543),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2562),
.A2(n_2506),
.B(n_2539),
.Y(n_2571)
);

AND2x4_ASAP7_75t_L g2572 ( 
.A(n_2545),
.B(n_2513),
.Y(n_2572)
);

AOI22xp5_ASAP7_75t_L g2573 ( 
.A1(n_2553),
.A2(n_2536),
.B1(n_380),
.B2(n_381),
.Y(n_2573)
);

INVx2_ASAP7_75t_SL g2574 ( 
.A(n_2552),
.Y(n_2574)
);

INVxp67_ASAP7_75t_L g2575 ( 
.A(n_2557),
.Y(n_2575)
);

OAI22xp5_ASAP7_75t_L g2576 ( 
.A1(n_2559),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2556),
.Y(n_2577)
);

INVx1_ASAP7_75t_L g2578 ( 
.A(n_2561),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2551),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2560),
.B(n_379),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2563),
.A2(n_382),
.B(n_383),
.Y(n_2581)
);

AO22x2_ASAP7_75t_L g2582 ( 
.A1(n_2550),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_2582)
);

NAND5xp2_ASAP7_75t_L g2583 ( 
.A(n_2554),
.B(n_384),
.C(n_385),
.D(n_386),
.E(n_387),
.Y(n_2583)
);

AO22x1_ASAP7_75t_L g2584 ( 
.A1(n_2567),
.A2(n_2546),
.B1(n_2558),
.B2(n_2564),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2576),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2573),
.B(n_2555),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2572),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2581),
.Y(n_2588)
);

OA22x2_ASAP7_75t_L g2589 ( 
.A1(n_2578),
.A2(n_2548),
.B1(n_389),
.B2(n_390),
.Y(n_2589)
);

AO22x1_ASAP7_75t_L g2590 ( 
.A1(n_2577),
.A2(n_388),
.B1(n_391),
.B2(n_392),
.Y(n_2590)
);

NOR2x1p5_ASAP7_75t_L g2591 ( 
.A(n_2579),
.B(n_391),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2580),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2582),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2582),
.Y(n_2594)
);

XOR2xp5_ASAP7_75t_L g2595 ( 
.A(n_2569),
.B(n_393),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2589),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2591),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2595),
.Y(n_2598)
);

NOR2xp67_ASAP7_75t_SL g2599 ( 
.A(n_2587),
.B(n_2568),
.Y(n_2599)
);

CKINVDCx16_ASAP7_75t_R g2600 ( 
.A(n_2592),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2593),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2585),
.A2(n_2574),
.B1(n_2570),
.B2(n_2588),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2594),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2599),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2597),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2596),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2601),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2603),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2600),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2598),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2604),
.B(n_2566),
.Y(n_2611)
);

AOI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2609),
.A2(n_2575),
.B1(n_2586),
.B2(n_2584),
.Y(n_2612)
);

OAI21xp5_ASAP7_75t_L g2613 ( 
.A1(n_2607),
.A2(n_2571),
.B(n_2602),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2608),
.A2(n_2590),
.B1(n_2583),
.B2(n_395),
.Y(n_2614)
);

OAI22xp33_ASAP7_75t_L g2615 ( 
.A1(n_2606),
.A2(n_393),
.B1(n_394),
.B2(n_395),
.Y(n_2615)
);

AOI21x1_ASAP7_75t_L g2616 ( 
.A1(n_2611),
.A2(n_2605),
.B(n_2610),
.Y(n_2616)
);

OAI21xp5_ASAP7_75t_L g2617 ( 
.A1(n_2612),
.A2(n_396),
.B(n_397),
.Y(n_2617)
);

AOI22xp33_ASAP7_75t_L g2618 ( 
.A1(n_2617),
.A2(n_2613),
.B1(n_2614),
.B2(n_2615),
.Y(n_2618)
);

XOR2xp5_ASAP7_75t_L g2619 ( 
.A(n_2616),
.B(n_396),
.Y(n_2619)
);

OA21x2_ASAP7_75t_L g2620 ( 
.A1(n_2618),
.A2(n_399),
.B(n_400),
.Y(n_2620)
);

AOI21xp33_ASAP7_75t_L g2621 ( 
.A1(n_2619),
.A2(n_401),
.B(n_402),
.Y(n_2621)
);

AOI222xp33_ASAP7_75t_L g2622 ( 
.A1(n_2620),
.A2(n_401),
.B1(n_402),
.B2(n_403),
.C1(n_404),
.C2(n_405),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_SL g2623 ( 
.A1(n_2621),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_2623)
);

OAI21xp5_ASAP7_75t_L g2624 ( 
.A1(n_2623),
.A2(n_406),
.B(n_407),
.Y(n_2624)
);

AOI322xp5_ASAP7_75t_L g2625 ( 
.A1(n_2624),
.A2(n_2622),
.A3(n_408),
.B1(n_409),
.B2(n_411),
.C1(n_412),
.C2(n_413),
.Y(n_2625)
);

AOI221xp5_ASAP7_75t_L g2626 ( 
.A1(n_2625),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.C(n_413),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_SL g2627 ( 
.A1(n_2626),
.A2(n_414),
.B1(n_415),
.B2(n_416),
.Y(n_2627)
);

AOI211xp5_ASAP7_75t_L g2628 ( 
.A1(n_2627),
.A2(n_414),
.B(n_416),
.C(n_417),
.Y(n_2628)
);


endmodule