module fake_jpeg_1536_n_262 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

INVx4_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_47),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_51),
.Y(n_86)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_44),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx6p67_ASAP7_75t_R g95 ( 
.A(n_45),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_7),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_19),
.B(n_23),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_58),
.Y(n_88)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_0),
.Y(n_58)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_19),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_60),
.B(n_61),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_6),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_66),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_20),
.B(n_10),
.Y(n_66)
);

INVx6_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_17),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_74),
.Y(n_98)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_22),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_76),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_39),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_73),
.A2(n_24),
.B1(n_36),
.B2(n_30),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_79),
.A2(n_68),
.B1(n_13),
.B2(n_14),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_50),
.B(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_30),
.B1(n_36),
.B2(n_28),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_54),
.B1(n_76),
.B2(n_53),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_67),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_94),
.B1(n_99),
.B2(n_109),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_39),
.B1(n_32),
.B2(n_31),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_57),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_32),
.B1(n_27),
.B2(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_54),
.B1(n_72),
.B2(n_71),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_66),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_45),
.A2(n_27),
.B1(n_0),
.B2(n_3),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_5),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_110),
.B(n_95),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_113),
.A2(n_96),
.B1(n_84),
.B2(n_80),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_45),
.A2(n_4),
.B1(n_11),
.B2(n_12),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_52),
.B1(n_64),
.B2(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_58),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_119),
.B(n_124),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_120),
.A2(n_146),
.B1(n_151),
.B2(n_93),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_125),
.Y(n_159)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_44),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_41),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_88),
.B(n_49),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_135),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_63),
.C(n_48),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_82),
.C(n_105),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_62),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_143),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_137),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_141),
.B1(n_142),
.B2(n_105),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_68),
.B1(n_59),
.B2(n_14),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_129),
.B1(n_146),
.B2(n_133),
.Y(n_182)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_134),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_82),
.B1(n_120),
.B2(n_121),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_113),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_154),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_94),
.B1(n_91),
.B2(n_99),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_93),
.B1(n_83),
.B2(n_116),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_103),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_117),
.B1(n_83),
.B2(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_147),
.B(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_111),
.B(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_149),
.Y(n_180)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_84),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_114),
.A2(n_109),
.B(n_116),
.C(n_82),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_87),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_152),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_87),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_156),
.A2(n_158),
.B1(n_182),
.B2(n_154),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_118),
.B1(n_115),
.B2(n_80),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_135),
.Y(n_168)
);

XOR2x2_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_171),
.B(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_115),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_177),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_132),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_141),
.A2(n_151),
.B(n_150),
.Y(n_176)
);

NAND2xp33_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_164),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_145),
.B(n_127),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_123),
.B(n_134),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_132),
.B1(n_144),
.B2(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_184),
.A2(n_185),
.B1(n_193),
.B2(n_155),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_132),
.B1(n_121),
.B2(n_136),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_147),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_191),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_201),
.B(n_171),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_165),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_132),
.B1(n_138),
.B2(n_149),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_164),
.Y(n_208)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_180),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_202),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_197),
.B(n_168),
.C(n_177),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_178),
.A2(n_153),
.B(n_156),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_179),
.B(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_175),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_191),
.Y(n_218)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_164),
.A2(n_158),
.B1(n_182),
.B2(n_178),
.Y(n_200)
);

NAND2x1_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_163),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_203),
.B(n_199),
.Y(n_219)
);

A2O1A1O1Ixp25_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_183),
.B(n_188),
.C(n_197),
.D(n_195),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_207),
.B(n_214),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_208),
.A2(n_212),
.B1(n_217),
.B2(n_200),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_210),
.B(n_216),
.Y(n_225)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_197),
.B(n_166),
.C(n_167),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_201),
.A2(n_167),
.B(n_170),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_162),
.B1(n_170),
.B2(n_157),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_218),
.B(n_219),
.Y(n_224)
);

NOR3xp33_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_190),
.C(n_187),
.Y(n_221)
);

NOR3xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_206),
.C(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_205),
.B(n_196),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_229),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_183),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_185),
.B1(n_198),
.B2(n_184),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_208),
.B1(n_200),
.B2(n_194),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_219),
.B(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_210),
.B(n_215),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_233),
.B(n_225),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_236),
.A2(n_230),
.B1(n_223),
.B2(n_207),
.Y(n_244)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_238),
.Y(n_242)
);

XOR2x2_ASAP7_75t_SL g239 ( 
.A(n_227),
.B(n_210),
.Y(n_239)
);

AOI31xp67_ASAP7_75t_L g245 ( 
.A1(n_239),
.A2(n_240),
.A3(n_214),
.B(n_213),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_241),
.A2(n_245),
.B(n_235),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_224),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_234),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_246),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_249),
.B(n_251),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_232),
.B(n_240),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_206),
.B(n_236),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_192),
.Y(n_252)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_250),
.B(n_233),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_250),
.A2(n_226),
.B1(n_239),
.B2(n_221),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_254),
.A2(n_255),
.B(n_188),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_258),
.A2(n_216),
.B(n_217),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g259 ( 
.A(n_256),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_260),
.C(n_257),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_202),
.Y(n_262)
);


endmodule