module real_jpeg_8519_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_285, n_284, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_285;
input n_284;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_211;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_205;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_253;
wire n_273;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_31),
.B1(n_41),
.B2(n_43),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_1),
.A2(n_31),
.B1(n_65),
.B2(n_66),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_19),
.B1(n_20),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_2),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_52),
.B1(n_65),
.B2(n_66),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_41),
.B1(n_43),
.B2(n_52),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_2),
.A2(n_6),
.B(n_66),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_38),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_27),
.B(n_40),
.C(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_29),
.Y(n_151)
);

AOI21xp33_ASAP7_75t_L g172 ( 
.A1(n_2),
.A2(n_3),
.B(n_28),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_3),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_3),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_4),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_6),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_64)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_6),
.A2(n_41),
.B(n_64),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_6),
.B(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_SL g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_9),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_9),
.A2(n_21),
.B1(n_27),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_9),
.A2(n_21),
.B1(n_65),
.B2(n_66),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_9),
.A2(n_21),
.B1(n_41),
.B2(n_43),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_10),
.A2(n_19),
.B1(n_20),
.B2(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_10),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_10),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_10),
.A2(n_41),
.B1(n_43),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_60),
.Y(n_130)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_74),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_73),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_32),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_32),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B1(n_29),
.B2(n_30),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_18),
.A2(n_26),
.B(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_20),
.A2(n_24),
.B(n_52),
.C(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_23),
.B(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_23),
.A2(n_26),
.B1(n_51),
.B2(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_23),
.B(n_26),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_26),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_27),
.A2(n_39),
.B(n_40),
.C(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_40),
.Y(n_47)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_29),
.A2(n_50),
.B(n_59),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_33),
.B(n_281),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_33),
.B(n_281),
.Y(n_282)
);

FAx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_48),
.CI(n_53),
.CON(n_33),
.SN(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_36),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_38),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_37),
.B(n_132),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_45),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_38),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_38),
.A2(n_45),
.B1(n_130),
.B2(n_147),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_39),
.A2(n_259),
.B(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_SL g136 ( 
.A1(n_41),
.A2(n_44),
.B(n_52),
.Y(n_136)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_43),
.A2(n_52),
.B(n_69),
.C(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_46),
.B(n_132),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_51),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_52),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_52),
.B(n_64),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.C(n_61),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_54),
.A2(n_61),
.B1(n_261),
.B2(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_54),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_55),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_56),
.A2(n_57),
.B1(n_146),
.B2(n_152),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_56),
.B(n_146),
.C(n_189),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_56),
.A2(n_57),
.B1(n_129),
.B2(n_133),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_56),
.B(n_129),
.C(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_56),
.A2(n_57),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_61),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_61),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_72),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_63),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_70),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_64),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_64),
.A2(n_70),
.B1(n_95),
.B2(n_98),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_64),
.A2(n_224),
.B(n_225),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_64),
.A2(n_70),
.B1(n_72),
.B2(n_224),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_65),
.B(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_280),
.B(n_282),
.Y(n_74)
);

OAI321xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_253),
.A3(n_273),
.B1(n_278),
.B2(n_279),
.C(n_284),
.Y(n_75)
);

AOI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_208),
.A3(n_228),
.B1(n_247),
.B2(n_252),
.C(n_285),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_177),
.C(n_205),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_157),
.B(n_176),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_142),
.B(n_156),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_124),
.B(n_141),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_113),
.B(n_123),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_103),
.B(n_112),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_84),
.B(n_92),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_84),
.A2(n_105),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_84),
.B(n_146),
.C(n_151),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_87),
.B(n_88),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_87),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_87),
.B(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_87),
.A2(n_139),
.B1(n_184),
.B2(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_88),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_89),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_90),
.A2(n_183),
.B(n_185),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_100),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_102),
.B1(n_129),
.B2(n_133),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_129),
.C(n_140),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_93),
.A2(n_102),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_97),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_98),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_182),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_108),
.B(n_111),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_116),
.B1(n_117),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_118),
.C(n_121),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_122),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_110),
.B(n_170),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_115),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_121),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_120),
.A2(n_121),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_196),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_145),
.C(n_155),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_126),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_134),
.B2(n_140),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_129),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_133),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_163),
.C(n_167),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_138),
.B(n_198),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_144),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_153),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_146),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_152),
.A2(n_234),
.B(n_235),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_152),
.B(n_234),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_154),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_158),
.B(n_159),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_168),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_169),
.C(n_175),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_166),
.B2(n_167),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_166),
.A2(n_167),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_166),
.A2(n_167),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_166),
.A2(n_167),
.B1(n_267),
.B2(n_271),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_166),
.B(n_261),
.C(n_262),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_166),
.B(n_271),
.C(n_272),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_167),
.B(n_200),
.C(n_202),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_169),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_173),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

AOI21xp33_ASAP7_75t_L g248 ( 
.A1(n_178),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_190),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_179),
.B(n_190),
.Y(n_250)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_186),
.CI(n_187),
.CON(n_179),
.SN(n_179)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_204),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_199),
.C(n_204),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_207),
.Y(n_249)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_209),
.A2(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_210),
.B(n_211),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_227),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_220),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_220),
.C(n_227),
.Y(n_229)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_215),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_226),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_222),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_223),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_237),
.B(n_239),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_245),
.B2(n_246),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_236),
.B1(n_243),
.B2(n_244),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_233),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_244),
.C(n_246),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_255),
.C(n_263),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_235),
.B(n_255),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_236),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_239),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_265),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_265),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_258),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_263),
.A2(n_264),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_272),
.Y(n_265)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_267),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);


endmodule