module real_jpeg_18361_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_83;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_1),
.A2(n_14),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_1),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_1),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_1),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_1),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_1),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_1),
.B(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_2),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_2),
.Y(n_161)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_2),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_3),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_3),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_3),
.B(n_319),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_3),
.B(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_4),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_4),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_4),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_4),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_4),
.B(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_4),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_4),
.B(n_157),
.Y(n_387)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_5),
.Y(n_169)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_5),
.Y(n_347)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_5),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_73),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_7),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_7),
.B(n_205),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_7),
.B(n_210),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_7),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_8),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_8),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_8),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_8),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_8),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_8),
.B(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_9),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_10),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_10),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_10),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_10),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_10),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_12),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_13),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_13),
.B(n_233),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_13),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_13),
.B(n_363),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_13),
.B(n_167),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_13),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_13),
.B(n_415),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_14),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_14),
.B(n_163),
.Y(n_221)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_14),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_14),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_14),
.B(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_14),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_14),
.B(n_505),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_15),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_16),
.Y(n_58)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_16),
.Y(n_126)
);

BUFx4f_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_17),
.Y(n_304)
);

BUFx5_ASAP7_75t_L g455 ( 
.A(n_17),
.Y(n_455)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

A2O1A1O1Ixp25_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_438),
.B(n_525),
.C(n_532),
.D(n_534),
.Y(n_22)
);

NAND2x1_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_329),
.Y(n_23)
);

A2O1A1O1Ixp25_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_225),
.B(n_288),
.C(n_289),
.D(n_328),
.Y(n_24)
);

NAND4xp25_ASAP7_75t_L g329 ( 
.A(n_25),
.B(n_289),
.C(n_330),
.D(n_332),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_178),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_26),
.B(n_178),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_102),
.C(n_148),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_27),
.A2(n_28),
.B1(n_103),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_68),
.Y(n_28)
);

INVxp33_ASAP7_75t_SL g180 ( 
.A(n_29),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_43),
.C(n_51),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_30),
.B(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_35),
.C(n_39),
.Y(n_91)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_32),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_32),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_39),
.B2(n_42),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_38),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_39),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_39),
.B(n_209),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_40),
.Y(n_250)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_42),
.B(n_209),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_43),
.A2(n_44),
.B1(n_51),
.B2(n_52),
.Y(n_280)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_44),
.A2(n_242),
.B(n_247),
.Y(n_241)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_50),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.C(n_64),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_53),
.B(n_64),
.Y(n_151)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_58),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_58),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_59),
.B(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_63),
.Y(n_220)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_67),
.Y(n_320)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_67),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_90),
.B1(n_100),
.B2(n_101),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_69),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B(n_75),
.C(n_87),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_70),
.A2(n_72),
.B1(n_88),
.B2(n_89),
.Y(n_177)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_73),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_74),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_75),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_83),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_76),
.A2(n_83),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_76),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_76),
.A2(n_166),
.B1(n_253),
.B2(n_263),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_76),
.B(n_263),
.C(n_463),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_76),
.A2(n_131),
.B1(n_132),
.B2(n_253),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_79),
.B(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g506 ( 
.A(n_81),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_82),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_83),
.B(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_83),
.Y(n_254)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_99),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_94),
.B(n_98),
.C(n_99),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_97),
.A2(n_98),
.B1(n_131),
.B2(n_132),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_97),
.A2(n_98),
.B1(n_204),
.B2(n_521),
.Y(n_520)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_97),
.B(n_452),
.C(n_521),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_98),
.B(n_131),
.C(n_318),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_101),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_103),
.Y(n_286)
);

XNOR2x1_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_116),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_130),
.C(n_146),
.Y(n_186)
);

XNOR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_105),
.B(n_109),
.C(n_113),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_111),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_112),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_113),
.A2(n_448),
.B1(n_449),
.B2(n_450),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_113),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_113),
.B(n_449),
.C(n_452),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_115),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_130),
.B1(n_146),
.B2(n_147),
.Y(n_116)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_118),
.B(n_122),
.C(n_129),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_119),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_119),
.B(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_129),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_122),
.A2(n_123),
.B1(n_154),
.B2(n_155),
.Y(n_264)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_127),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_127),
.A2(n_129),
.B1(n_209),
.B2(n_213),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_127),
.B(n_349),
.Y(n_393)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_128),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_129),
.B(n_204),
.C(n_209),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_129),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_137),
.C(n_142),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_132),
.B1(n_142),
.B2(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_132),
.B(n_253),
.C(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_137),
.A2(n_138),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_137),
.A2(n_138),
.B1(n_322),
.B2(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_138),
.B(n_318),
.C(n_327),
.Y(n_466)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_141),
.Y(n_403)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_142),
.Y(n_174)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_148),
.B(n_285),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_170),
.C(n_175),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_149),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_158),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_150),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_152),
.A2(n_153),
.B1(n_158),
.B2(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_158),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_166),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_159),
.A2(n_166),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_159),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_162),
.B(n_261),
.Y(n_260)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_166),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_166),
.A2(n_209),
.B1(n_213),
.B2(n_263),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_166),
.B(n_213),
.C(n_312),
.Y(n_467)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_171),
.B(n_176),
.Y(n_277)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_179),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.C(n_182),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_202),
.B1(n_223),
.B2(n_224),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_184),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_201),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_185),
.B(n_188),
.C(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_200),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_190),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_199),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_193),
.B(n_196),
.C(n_199),
.Y(n_300)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_196),
.A2(n_197),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_196),
.B(n_479),
.C(n_482),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_197),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_197),
.B(n_307),
.C(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_202),
.B(n_223),
.C(n_291),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_214),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_203),
.B(n_215),
.C(n_216),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.Y(n_203)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_204),
.Y(n_521)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_222),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_218),
.B(n_222),
.C(n_254),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_220),
.Y(n_369)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_221),
.Y(n_222)
);

OAI21x1_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_282),
.B(n_287),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_275),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g331 ( 
.A(n_227),
.B(n_275),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_255),
.C(n_259),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_228),
.B(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_240),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_241),
.C(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.C(n_237),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_230),
.B(n_339),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_339)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_251),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_255),
.A2(n_256),
.B1(n_259),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_259),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.C(n_265),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_260),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_264),
.B(n_265),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_272),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_266),
.B(n_272),
.Y(n_375)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_269),
.B(n_375),
.Y(n_374)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_271),
.Y(n_366)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_274),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_281),
.Y(n_278)
);

NOR2x1_ASAP7_75t_L g330 ( 
.A(n_282),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_292),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_293),
.B(n_296),
.C(n_309),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_309),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_308),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_297),
.B(n_300),
.C(n_301),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

AO22x1_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_302),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_303),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_305),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_315),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_310),
.B(n_316),
.C(n_317),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_313),
.B(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_313),
.B(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_318),
.B(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_322),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_355),
.B(n_437),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_352),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_334),
.B(n_352),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_340),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_335),
.A2(n_336),
.B1(n_377),
.B2(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_338),
.B(n_340),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.C(n_348),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_341),
.Y(n_360)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_346),
.Y(n_425)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_348),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI21x1_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_379),
.B(n_436),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_376),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_357),
.B(n_376),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_374),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_358),
.B(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_361),
.B(n_374),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_367),
.C(n_370),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_370),
.Y(n_384)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI21x1_ASAP7_75t_L g379 ( 
.A1(n_380),
.A2(n_396),
.B(n_435),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_394),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_381),
.B(n_394),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.C(n_392),
.Y(n_381)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_382),
.A2(n_383),
.B1(n_406),
.B2(n_408),
.Y(n_405)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_385),
.A2(n_392),
.B1(n_393),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_386),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_399)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_409),
.B(n_434),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_405),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_398),
.B(n_405),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.C(n_404),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_399),
.B(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_400),
.A2(n_401),
.B1(n_404),
.B2(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_404),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_406),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_410),
.A2(n_420),
.B(n_433),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_417),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_411),
.B(n_417),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_414),
.Y(n_426)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_427),
.B(n_432),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_426),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_422),
.B(n_426),
.Y(n_432)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_494),
.C(n_514),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_490),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g527 ( 
.A1(n_441),
.A2(n_528),
.B(n_529),
.Y(n_527)
);

NOR2xp67_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_484),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_442),
.B(n_484),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_459),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_443),
.B(n_460),
.C(n_468),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.C(n_457),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_444),
.B(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_457),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_447),
.B1(n_452),
.B2(n_456),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_452),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_452),
.A2(n_456),
.B1(n_520),
.B2(n_522),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_454),
.Y(n_453)
);

INVx8_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_458),
.A2(n_518),
.B(n_533),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_468),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_466),
.C(n_467),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_488),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_467),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_477),
.B2(n_478),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_471),
.B(n_472),
.C(n_477),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_476),
.Y(n_472)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_473),
.Y(n_508)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_487),
.C(n_489),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_485),
.B(n_487),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_492),
.Y(n_491)
);

OR2x6_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_493),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_493),
.Y(n_528)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

A2O1A1O1Ixp25_ASAP7_75t_L g526 ( 
.A1(n_495),
.A2(n_515),
.B(n_527),
.C(n_530),
.D(n_531),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_513),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_496),
.B(n_513),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_499),
.C(n_512),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_500),
.B1(n_511),
.B2(n_512),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_499),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_500),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_501),
.B(n_507),
.C(n_509),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_507),
.B1(n_509),
.B2(n_510),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g509 ( 
.A(n_504),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_507),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_524),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_516),
.B(n_524),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_523),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_519),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g522 ( 
.A(n_520),
.Y(n_522)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_533),
.Y(n_532)
);


endmodule