module fake_jpeg_12446_n_604 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_604);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_604;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_12),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g148 ( 
.A(n_61),
.Y(n_148)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_31),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_83),
.Y(n_124)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g190 ( 
.A(n_66),
.Y(n_190)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_19),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_74),
.Y(n_161)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_78),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_24),
.B(n_9),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_86),
.Y(n_186)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

CKINVDCx9p33_ASAP7_75t_R g193 ( 
.A(n_88),
.Y(n_193)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_39),
.B(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_110),
.Y(n_127)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_92),
.Y(n_163)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_93),
.Y(n_179)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_96),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_30),
.Y(n_101)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_37),
.Y(n_103)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_104),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_105),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_106),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_107),
.Y(n_196)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_45),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_111),
.Y(n_173)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_112),
.B(n_113),
.Y(n_178)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_41),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_114),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_41),
.Y(n_115)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_118),
.Y(n_142)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_28),
.Y(n_117)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_26),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_122),
.Y(n_170)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_28),
.Y(n_121)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_83),
.B(n_46),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_129),
.B(n_145),
.Y(n_203)
);

OA22x2_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_43),
.B1(n_26),
.B2(n_39),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_135),
.A2(n_18),
.B(n_80),
.C(n_79),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_42),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_46),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_156),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_43),
.B1(n_56),
.B2(n_32),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_153),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_88),
.B(n_57),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_155),
.B(n_8),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_116),
.B(n_42),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_72),
.B(n_34),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_160),
.B(n_175),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_27),
.B1(n_43),
.B2(n_57),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_168),
.A2(n_177),
.B1(n_180),
.B2(n_23),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_56),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_60),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_176),
.B(n_183),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_115),
.A2(n_27),
.B1(n_52),
.B2(n_51),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_102),
.A2(n_52),
.B1(n_51),
.B2(n_50),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_114),
.B(n_34),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_103),
.A2(n_55),
.B(n_29),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_187),
.B(n_29),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_58),
.B(n_55),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_109),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_73),
.B(n_48),
.C(n_44),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_90),
.C(n_86),
.Y(n_248)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_200),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_204),
.Y(n_278)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_205),
.Y(n_303)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_206),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_148),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_207),
.B(n_222),
.Y(n_294)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_208),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_128),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_209),
.B(n_219),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_135),
.B1(n_143),
.B2(n_157),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_210),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_127),
.A2(n_168),
.B1(n_177),
.B2(n_124),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_211),
.A2(n_234),
.B1(n_244),
.B2(n_268),
.Y(n_279)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_125),
.B(n_0),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_214),
.Y(n_281)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_141),
.Y(n_213)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_148),
.Y(n_215)
);

INVx4_ASAP7_75t_SL g290 ( 
.A(n_215),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_126),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_220),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_221),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_142),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_223),
.A2(n_253),
.B1(n_257),
.B2(n_262),
.Y(n_285)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_190),
.Y(n_224)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_224),
.Y(n_291)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_225),
.Y(n_295)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_226),
.Y(n_300)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_136),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_228),
.B(n_231),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g229 ( 
.A1(n_127),
.A2(n_124),
.A3(n_170),
.B1(n_176),
.B2(n_154),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_229),
.B(n_236),
.Y(n_299)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_230),
.Y(n_297)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

AO22x1_ASAP7_75t_SL g232 ( 
.A1(n_137),
.A2(n_48),
.B1(n_44),
.B2(n_111),
.Y(n_232)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_232),
.A2(n_165),
.B1(n_162),
.B2(n_166),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_233),
.B(n_241),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_74),
.B1(n_107),
.B2(n_106),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_235),
.B(n_239),
.Y(n_314)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_159),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_237),
.B(n_240),
.Y(n_322)
);

INVx3_ASAP7_75t_SL g238 ( 
.A(n_147),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_238),
.B(n_247),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_142),
.B(n_17),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_164),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_170),
.A2(n_17),
.B(n_13),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_242),
.B(n_246),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_131),
.Y(n_243)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_243),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_155),
.A2(n_105),
.B1(n_100),
.B2(n_99),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_245),
.A2(n_199),
.B1(n_133),
.B2(n_18),
.Y(n_315)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_194),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_248),
.B(n_252),
.Y(n_324)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_198),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_249),
.Y(n_274)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_251),
.Y(n_289)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_132),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_255),
.B(n_260),
.Y(n_317)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_132),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g304 ( 
.A1(n_258),
.A2(n_266),
.B(n_268),
.C(n_232),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_184),
.A2(n_85),
.B1(n_78),
.B2(n_18),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_162),
.C(n_161),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_172),
.B(n_10),
.Y(n_260)
);

INVx11_ASAP7_75t_L g261 ( 
.A(n_163),
.Y(n_261)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_261),
.Y(n_286)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_171),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_181),
.B(n_188),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_263),
.B(n_10),
.Y(n_326)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_130),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_264),
.A2(n_265),
.B1(n_267),
.B2(n_269),
.Y(n_308)
);

INVx6_ASAP7_75t_L g265 ( 
.A(n_161),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_138),
.A2(n_18),
.B(n_10),
.Y(n_266)
);

INVx11_ASAP7_75t_L g267 ( 
.A(n_144),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_149),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_211),
.A2(n_167),
.B1(n_189),
.B2(n_152),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_270),
.A2(n_307),
.B1(n_259),
.B2(n_245),
.Y(n_331)
);

CKINVDCx12_ASAP7_75t_R g271 ( 
.A(n_201),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_271),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_293),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_218),
.B(n_123),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_282),
.B(n_296),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_212),
.B(n_186),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_212),
.B(n_186),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_301),
.B(n_305),
.Y(n_360)
);

NOR4xp25_ASAP7_75t_SL g302 ( 
.A(n_214),
.B(n_15),
.C(n_17),
.D(n_16),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_302),
.A2(n_266),
.B(n_281),
.Y(n_329)
);

O2A1O1Ixp33_ASAP7_75t_L g366 ( 
.A1(n_304),
.A2(n_4),
.B(n_1),
.C(n_3),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_229),
.B(n_140),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_221),
.A2(n_140),
.B1(n_166),
.B2(n_165),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g313 ( 
.A(n_250),
.B(n_182),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_319),
.C(n_216),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_325),
.B1(n_215),
.B2(n_238),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g316 ( 
.A(n_203),
.B(n_10),
.CI(n_16),
.CON(n_316),
.SN(n_316)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_316),
.B(n_5),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_217),
.B(n_6),
.C(n_14),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_223),
.A2(n_6),
.B1(n_13),
.B2(n_11),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_320),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_326),
.B(n_17),
.Y(n_350)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_327),
.Y(n_374)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_328),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_329),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_330),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_331),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_299),
.A2(n_235),
.B(n_248),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_363),
.B(n_366),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_305),
.A2(n_258),
.B1(n_232),
.B2(n_269),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_342),
.B1(n_353),
.B2(n_309),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_304),
.A2(n_228),
.B1(n_251),
.B2(n_257),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_334),
.A2(n_355),
.B1(n_365),
.B2(n_289),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_264),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_335),
.B(n_341),
.Y(n_390)
);

AO22x1_ASAP7_75t_SL g336 ( 
.A1(n_279),
.A2(n_267),
.B1(n_261),
.B2(n_265),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_361),
.Y(n_391)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_318),
.Y(n_337)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_318),
.Y(n_338)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_338),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_339),
.B(n_362),
.Y(n_384)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_276),
.Y(n_340)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_262),
.Y(n_341)
);

OAI22x1_ASAP7_75t_SL g342 ( 
.A1(n_279),
.A2(n_249),
.B1(n_231),
.B2(n_247),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_343),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_347),
.Y(n_373)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_323),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_348),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_285),
.A2(n_224),
.B(n_200),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_349),
.A2(n_369),
.B(n_275),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_350),
.B(n_357),
.Y(n_393)
);

NOR2x1_ASAP7_75t_R g351 ( 
.A(n_321),
.B(n_202),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_351),
.A2(n_290),
.B(n_286),
.Y(n_407)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_356),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_324),
.A2(n_253),
.B1(n_243),
.B2(n_204),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_281),
.B(n_256),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_354),
.B(n_358),
.C(n_288),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_277),
.A2(n_282),
.B1(n_313),
.B2(n_325),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_311),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_314),
.B(n_317),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_281),
.B(n_287),
.C(n_301),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_296),
.B(n_230),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_1),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_295),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_364),
.A2(n_368),
.B1(n_283),
.B2(n_300),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_287),
.A2(n_11),
.B1(n_13),
.B2(n_4),
.Y(n_365)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_288),
.A2(n_1),
.B(n_4),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_402),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_372),
.B(n_351),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_319),
.C(n_306),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_379),
.C(n_403),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_306),
.C(n_298),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_360),
.A2(n_293),
.B1(n_312),
.B2(n_316),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_386),
.B1(n_388),
.B2(n_398),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_387),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_360),
.A2(n_293),
.B1(n_312),
.B2(n_302),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_329),
.A2(n_326),
.B(n_288),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_389),
.A2(n_362),
.B(n_366),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_333),
.A2(n_293),
.B1(n_289),
.B2(n_309),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_396),
.A2(n_400),
.B1(n_406),
.B2(n_330),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_355),
.A2(n_308),
.B1(n_311),
.B2(n_274),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_365),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_399),
.B(n_391),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_309),
.B1(n_274),
.B2(n_298),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_359),
.A2(n_283),
.B1(n_291),
.B2(n_284),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_401),
.A2(n_407),
.B(n_408),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_334),
.A2(n_278),
.B1(n_303),
.B2(n_280),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_339),
.B(n_303),
.C(n_310),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_332),
.A2(n_278),
.B1(n_310),
.B2(n_273),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_337),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_359),
.A2(n_273),
.B1(n_291),
.B2(n_284),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_409),
.A2(n_429),
.B(n_407),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_383),
.Y(n_410)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_410),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_347),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_411),
.B(n_421),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_345),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_413),
.C(n_415),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_372),
.B(n_345),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_414),
.A2(n_416),
.B1(n_419),
.B2(n_433),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_340),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_378),
.A2(n_336),
.B1(n_361),
.B2(n_342),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_397),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_417),
.Y(n_445)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_418),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_378),
.A2(n_336),
.B1(n_370),
.B2(n_344),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_373),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_443),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_353),
.Y(n_421)
);

XNOR2x1_ASAP7_75t_L g459 ( 
.A(n_423),
.B(n_377),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_393),
.B(n_373),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_432),
.Y(n_472)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_427),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_381),
.A2(n_370),
.B(n_349),
.Y(n_429)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_275),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_327),
.B1(n_338),
.B2(n_363),
.Y(n_433)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_434),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_346),
.Y(n_435)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

OAI21xp33_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_368),
.B(n_364),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_437),
.A2(n_439),
.B(n_401),
.Y(n_447)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_374),
.Y(n_438)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_367),
.B(n_369),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_379),
.B(n_367),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g469 ( 
.A(n_440),
.B(n_377),
.Y(n_469)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_382),
.Y(n_441)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_441),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_390),
.B(n_328),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_376),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_387),
.A2(n_356),
.B1(n_343),
.B2(n_352),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_435),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_446),
.B(n_460),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_447),
.A2(n_452),
.B(n_430),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_403),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_451),
.B(n_453),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_430),
.A2(n_401),
.B(n_400),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_403),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_465),
.C(n_473),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_420),
.B(n_382),
.Y(n_457)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_427),
.B(n_406),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

XNOR2x1_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_440),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_434),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_415),
.B(n_384),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_418),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_431),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_SL g491 ( 
.A(n_469),
.B(n_475),
.Y(n_491)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_412),
.B(n_389),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_474),
.B(n_376),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g475 ( 
.A(n_413),
.B(n_385),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_441),
.Y(n_476)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_476),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_493),
.Y(n_506)
);

INVx13_ASAP7_75t_L g479 ( 
.A(n_445),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_479),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_463),
.A2(n_424),
.B1(n_426),
.B2(n_422),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_481),
.A2(n_500),
.B1(n_501),
.B2(n_388),
.Y(n_508)
);

AO22x1_ASAP7_75t_L g482 ( 
.A1(n_450),
.A2(n_409),
.B1(n_429),
.B2(n_426),
.Y(n_482)
);

A2O1A1Ixp33_ASAP7_75t_L g520 ( 
.A1(n_482),
.A2(n_480),
.B(n_487),
.C(n_478),
.Y(n_520)
);

OAI21xp33_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_423),
.B(n_422),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_483),
.B(n_498),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_472),
.Y(n_484)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_484),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_456),
.B(n_438),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_485),
.Y(n_524)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_444),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_487),
.B(n_488),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_444),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_454),
.A2(n_426),
.B1(n_414),
.B2(n_458),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_490),
.A2(n_502),
.B1(n_503),
.B2(n_439),
.Y(n_512)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_448),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_492),
.B(n_497),
.Y(n_526)
);

CKINVDCx14_ASAP7_75t_R g509 ( 
.A(n_496),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_449),
.B(n_405),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_499),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_463),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_456),
.A2(n_424),
.B1(n_454),
.B2(n_395),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_452),
.A2(n_386),
.B1(n_443),
.B2(n_419),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_447),
.A2(n_398),
.B1(n_433),
.B2(n_416),
.Y(n_503)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_502),
.A2(n_453),
.B1(n_399),
.B2(n_470),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_507),
.A2(n_512),
.B1(n_481),
.B2(n_480),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_503),
.B1(n_490),
.B2(n_478),
.Y(n_534)
);

BUFx24_ASAP7_75t_SL g510 ( 
.A(n_496),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_510),
.B(n_521),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_449),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_513),
.B(n_516),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_494),
.B(n_451),
.C(n_455),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_525),
.C(n_495),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_494),
.B(n_473),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_500),
.Y(n_517)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_469),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_518),
.B(n_519),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_489),
.B(n_459),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_520),
.B(n_477),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_465),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_482),
.B(n_475),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_482),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_462),
.C(n_467),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_528),
.B(n_541),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_509),
.B(n_501),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_529),
.B(n_543),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_505),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_530),
.B(n_538),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_488),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_531),
.B(n_542),
.Y(n_547)
);

XOR2x1_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_537),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_534),
.A2(n_511),
.B1(n_525),
.B2(n_506),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_545),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_476),
.B1(n_485),
.B2(n_486),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_515),
.B(n_499),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_517),
.A2(n_486),
.B1(n_466),
.B2(n_467),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_523),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_516),
.B(n_445),
.C(n_466),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_544),
.B(n_546),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_506),
.B(n_392),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_526),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g572 ( 
.A1(n_548),
.A2(n_555),
.B1(n_549),
.B2(n_554),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_541),
.B(n_513),
.C(n_518),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_550),
.B(n_551),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_531),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_537),
.A2(n_520),
.B(n_504),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_375),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_531),
.A2(n_514),
.B(n_522),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g564 ( 
.A1(n_555),
.A2(n_557),
.B(n_535),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_533),
.B(n_519),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_SL g571 ( 
.A(n_556),
.B(n_560),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_L g557 ( 
.A1(n_532),
.A2(n_504),
.B(n_527),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_544),
.B(n_461),
.C(n_417),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_558),
.B(n_542),
.C(n_528),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_392),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_558),
.Y(n_563)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_563),
.Y(n_583)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_564),
.A2(n_575),
.B(n_404),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_565),
.B(n_566),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_552),
.A2(n_540),
.B1(n_471),
.B2(n_464),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_559),
.B(n_539),
.C(n_536),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_567),
.B(n_570),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_561),
.A2(n_557),
.B1(n_547),
.B2(n_549),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g585 ( 
.A(n_568),
.B(n_397),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_562),
.B(n_397),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_569),
.B(n_560),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_547),
.A2(n_545),
.B1(n_402),
.B2(n_380),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_572),
.B(n_573),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g573 ( 
.A1(n_548),
.A2(n_380),
.B1(n_371),
.B2(n_479),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_565),
.B(n_550),
.C(n_539),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_577),
.B(n_579),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_574),
.B(n_553),
.C(n_556),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_581),
.B(n_585),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_567),
.A2(n_553),
.B(n_375),
.Y(n_582)
);

AO21x1_ASAP7_75t_L g587 ( 
.A1(n_582),
.A2(n_584),
.B(n_564),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_587),
.B(n_590),
.Y(n_595)
);

OAI21x1_ASAP7_75t_SL g588 ( 
.A1(n_578),
.A2(n_568),
.B(n_575),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_L g593 ( 
.A1(n_588),
.A2(n_589),
.B(n_584),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_SL g589 ( 
.A1(n_577),
.A2(n_571),
.B(n_404),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_576),
.B(n_571),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_404),
.C(n_290),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_592),
.B(n_585),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_593),
.A2(n_594),
.B(n_591),
.Y(n_598)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_586),
.A2(n_583),
.B(n_580),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_596),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_595),
.B(n_591),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_599),
.B(n_597),
.C(n_272),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_272),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_272),
.C(n_286),
.Y(n_602)
);

AND2x4_ASAP7_75t_SL g603 ( 
.A(n_602),
.B(n_272),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_603),
.A2(n_286),
.B(n_4),
.Y(n_604)
);


endmodule