module real_aes_8378_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_725;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g535 ( .A1(n_0), .A2(n_180), .B(n_536), .C(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_1), .B(n_486), .Y(n_540) );
NAND3xp33_ASAP7_75t_SL g108 ( .A(n_2), .B(n_87), .C(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g124 ( .A(n_2), .Y(n_124) );
INVx1_ASAP7_75t_L g192 ( .A(n_3), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_4), .B(n_152), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_5), .A2(n_459), .B(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g488 ( .A1(n_6), .A2(n_172), .B(n_489), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_7), .A2(n_35), .B1(n_146), .B2(n_201), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_8), .B(n_172), .Y(n_181) );
AND2x6_ASAP7_75t_L g164 ( .A(n_9), .B(n_165), .Y(n_164) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_10), .A2(n_164), .B(n_464), .C(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_11), .B(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
INVx1_ASAP7_75t_L g185 ( .A(n_13), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_14), .B(n_150), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_15), .B(n_152), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_16), .B(n_138), .Y(n_256) );
AO32x2_ASAP7_75t_L g198 ( .A1(n_17), .A2(n_137), .A3(n_163), .B1(n_172), .B2(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_18), .B(n_146), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_19), .B(n_138), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_20), .A2(n_50), .B1(n_146), .B2(n_201), .Y(n_202) );
AOI22xp33_ASAP7_75t_SL g240 ( .A1(n_21), .A2(n_77), .B1(n_146), .B2(n_150), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_22), .B(n_146), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_23), .A2(n_163), .B(n_464), .C(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_24), .A2(n_55), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_24), .Y(n_128) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_25), .A2(n_163), .B(n_464), .C(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_26), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_27), .B(n_167), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_28), .A2(n_459), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_29), .B(n_167), .Y(n_215) );
INVx2_ASAP7_75t_L g148 ( .A(n_30), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_31), .A2(n_462), .B(n_472), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g145 ( .A(n_32), .B(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_33), .B(n_167), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_34), .B(n_222), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_36), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_37), .B(n_511), .Y(n_510) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_38), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_39), .B(n_152), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_40), .B(n_459), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g461 ( .A1(n_41), .A2(n_462), .B(n_466), .C(n_472), .Y(n_461) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_42), .B(n_146), .Y(n_175) );
INVx1_ASAP7_75t_L g537 ( .A(n_43), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_44), .A2(n_88), .B1(n_201), .B2(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g467 ( .A(n_45), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_46), .B(n_146), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_47), .B(n_146), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_48), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_49), .B(n_158), .Y(n_179) );
AOI22xp33_ASAP7_75t_SL g254 ( .A1(n_51), .A2(n_56), .B1(n_146), .B2(n_150), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_52), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_53), .B(n_146), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_54), .B(n_146), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_55), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g446 ( .A1(n_55), .A2(n_129), .B1(n_130), .B2(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_57), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g165 ( .A(n_58), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_59), .B(n_459), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_60), .B(n_486), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_61), .A2(n_158), .B(n_188), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_62), .B(n_146), .Y(n_193) );
INVx1_ASAP7_75t_L g141 ( .A(n_63), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_64), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_65), .B(n_152), .Y(n_504) );
AO32x2_ASAP7_75t_L g236 ( .A1(n_66), .A2(n_163), .A3(n_172), .B1(n_237), .B2(n_241), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_67), .B(n_153), .Y(n_550) );
INVx1_ASAP7_75t_L g156 ( .A(n_68), .Y(n_156) );
INVx1_ASAP7_75t_L g210 ( .A(n_69), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g534 ( .A(n_70), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_71), .B(n_469), .Y(n_514) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_72), .A2(n_464), .B(n_472), .C(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_73), .B(n_150), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_74), .Y(n_481) );
INVx1_ASAP7_75t_L g111 ( .A(n_75), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_76), .B(n_468), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g441 ( .A1(n_78), .A2(n_82), .B1(n_442), .B2(n_750), .C1(n_755), .C2(n_756), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_79), .B(n_201), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_80), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_81), .B(n_150), .Y(n_214) );
INVx1_ASAP7_75t_L g755 ( .A(n_82), .Y(n_755) );
INVx2_ASAP7_75t_L g139 ( .A(n_83), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_84), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_85), .B(n_162), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_86), .B(n_150), .Y(n_176) );
OR2x2_ASAP7_75t_L g121 ( .A(n_87), .B(n_122), .Y(n_121) );
OR2x2_ASAP7_75t_L g445 ( .A(n_87), .B(n_123), .Y(n_445) );
INVx2_ASAP7_75t_L g451 ( .A(n_87), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_89), .A2(n_99), .B1(n_150), .B2(n_151), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_90), .B(n_459), .Y(n_500) );
INVx1_ASAP7_75t_L g503 ( .A(n_91), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_92), .A2(n_101), .B1(n_112), .B2(n_757), .Y(n_100) );
INVxp67_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_94), .B(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_95), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g525 ( .A(n_96), .Y(n_525) );
INVx1_ASAP7_75t_L g546 ( .A(n_97), .Y(n_546) );
AND2x2_ASAP7_75t_L g474 ( .A(n_98), .B(n_167), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_104), .Y(n_758) );
CKINVDCx9p33_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
OA211x2_ASAP7_75t_L g112 ( .A1(n_109), .A2(n_113), .B(n_118), .C(n_438), .Y(n_112) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g440 ( .A(n_115), .Y(n_440) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
OAI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_126), .B(n_434), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx2_ASAP7_75t_L g437 ( .A(n_121), .Y(n_437) );
NOR2x2_ASAP7_75t_L g756 ( .A(n_122), .B(n_451), .Y(n_756) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g450 ( .A(n_123), .B(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
XNOR2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_130), .Y(n_126) );
INVx1_ASAP7_75t_SL g447 ( .A(n_130), .Y(n_447) );
OR3x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_362), .C(n_411), .Y(n_130) );
NAND5xp2_ASAP7_75t_L g131 ( .A(n_132), .B(n_277), .C(n_305), .D(n_335), .E(n_349), .Y(n_131) );
AOI221xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_195), .B1(n_227), .B2(n_232), .C(n_243), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_134), .B(n_168), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_134), .B(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g257 ( .A(n_135), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_135), .B(n_171), .Y(n_265) );
AND2x2_ASAP7_75t_L g288 ( .A(n_135), .B(n_170), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_135), .B(n_182), .Y(n_303) );
OR2x2_ASAP7_75t_L g312 ( .A(n_135), .B(n_250), .Y(n_312) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_135), .Y(n_315) );
AND2x2_ASAP7_75t_L g423 ( .A(n_135), .B(n_250), .Y(n_423) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_143), .B(n_166), .Y(n_135) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_136), .A2(n_183), .B(n_194), .Y(n_182) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_137), .B(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_139), .B(n_140), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
OAI21xp5_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_155), .B(n_163), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_145), .A2(n_149), .B(n_152), .Y(n_144) );
INVx3_ASAP7_75t_L g209 ( .A(n_146), .Y(n_209) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_146), .Y(n_527) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
BUFx3_ASAP7_75t_L g239 ( .A(n_147), .Y(n_239) );
AND2x6_ASAP7_75t_L g464 ( .A(n_147), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g151 ( .A(n_148), .Y(n_151) );
INVx1_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx2_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g174 ( .A1(n_152), .A2(n_175), .B(n_176), .Y(n_174) );
INVx2_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
O2A1O1Ixp5_ASAP7_75t_SL g208 ( .A1(n_152), .A2(n_209), .B(n_210), .C(n_211), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_152), .B(n_484), .Y(n_483) );
INVx5_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g237 ( .A1(n_153), .A2(n_162), .B1(n_238), .B2(n_240), .Y(n_237) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_154), .Y(n_162) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_154), .Y(n_190) );
INVx1_ASAP7_75t_L g222 ( .A(n_154), .Y(n_222) );
AND2x2_ASAP7_75t_L g460 ( .A(n_154), .B(n_159), .Y(n_460) );
INVx1_ASAP7_75t_L g465 ( .A(n_154), .Y(n_465) );
O2A1O1Ixp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_157), .B(n_160), .C(n_161), .Y(n_155) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_157), .A2(n_180), .B(n_192), .C(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_157), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_161), .A2(n_224), .B(n_225), .Y(n_223) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_162), .A2(n_180), .B1(n_200), .B2(n_202), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_162), .A2(n_180), .B1(n_253), .B2(n_254), .Y(n_252) );
INVx4_ASAP7_75t_L g538 ( .A(n_162), .Y(n_538) );
NAND3xp33_ASAP7_75t_L g276 ( .A(n_163), .B(n_251), .C(n_252), .Y(n_276) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_164), .A2(n_174), .B(n_177), .Y(n_173) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_164), .A2(n_184), .B(n_191), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_164), .A2(n_208), .B(n_212), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_223), .Y(n_217) );
AND2x4_ASAP7_75t_L g459 ( .A(n_164), .B(n_460), .Y(n_459) );
INVx4_ASAP7_75t_SL g473 ( .A(n_164), .Y(n_473) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_164), .B(n_460), .Y(n_547) );
OA21x2_ASAP7_75t_L g206 ( .A1(n_167), .A2(n_207), .B(n_215), .Y(n_206) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_167), .A2(n_217), .B(n_226), .Y(n_216) );
INVx2_ASAP7_75t_L g241 ( .A(n_167), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_167), .A2(n_458), .B(n_461), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_167), .A2(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_167), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_168), .B(n_315), .Y(n_371) );
INVx2_ASAP7_75t_SL g168 ( .A(n_169), .Y(n_168) );
OAI311xp33_ASAP7_75t_L g313 ( .A1(n_169), .A2(n_314), .A3(n_315), .B1(n_316), .C1(n_331), .Y(n_313) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_182), .Y(n_169) );
AND2x2_ASAP7_75t_L g274 ( .A(n_170), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g281 ( .A(n_170), .Y(n_281) );
AND2x2_ASAP7_75t_L g402 ( .A(n_170), .B(n_231), .Y(n_402) );
INVx3_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_171), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g258 ( .A(n_171), .B(n_182), .Y(n_258) );
AND2x2_ASAP7_75t_L g310 ( .A(n_171), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g324 ( .A(n_171), .B(n_257), .Y(n_324) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_181), .Y(n_171) );
INVx4_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_172), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_172), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_180), .Y(n_177) );
INVx2_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
AND2x2_ASAP7_75t_L g273 ( .A(n_182), .B(n_257), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_186), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_186), .A2(n_550), .B(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_188), .A2(n_525), .B(n_526), .C(n_527), .Y(n_524) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_189), .A2(n_213), .B(n_214), .Y(n_212) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g469 ( .A(n_190), .Y(n_469) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_203), .Y(n_195) );
OR2x2_ASAP7_75t_L g368 ( .A(n_196), .B(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_196), .B(n_374), .Y(n_385) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_197), .B(n_381), .Y(n_380) );
BUFx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
AND2x2_ASAP7_75t_L g309 ( .A(n_198), .B(n_236), .Y(n_309) );
AND2x2_ASAP7_75t_L g320 ( .A(n_198), .B(n_216), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_198), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_203), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_203), .B(n_270), .Y(n_314) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g301 ( .A(n_204), .B(n_260), .Y(n_301) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_216), .Y(n_204) );
INVx2_ASAP7_75t_L g234 ( .A(n_205), .Y(n_234) );
AND2x2_ASAP7_75t_L g328 ( .A(n_205), .B(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
OR2x2_ASAP7_75t_L g345 ( .A(n_206), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_206), .Y(n_408) );
AND2x2_ASAP7_75t_L g247 ( .A(n_216), .B(n_242), .Y(n_247) );
INVx1_ASAP7_75t_L g268 ( .A(n_216), .Y(n_268) );
AND2x2_ASAP7_75t_L g289 ( .A(n_216), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g330 ( .A(n_216), .Y(n_330) );
INVx1_ASAP7_75t_L g346 ( .A(n_216), .Y(n_346) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_216), .Y(n_421) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_221), .Y(n_218) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVxp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_229), .B(n_334), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_229), .A2(n_319), .B1(n_368), .B2(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
OAI211xp5_ASAP7_75t_SL g411 ( .A1(n_230), .A2(n_412), .B(n_414), .C(n_432), .Y(n_411) );
INVx2_ASAP7_75t_L g264 ( .A(n_231), .Y(n_264) );
AND2x2_ASAP7_75t_L g322 ( .A(n_231), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g333 ( .A(n_231), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_232), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_235), .Y(n_232) );
AND2x2_ASAP7_75t_L g306 ( .A(n_233), .B(n_270), .Y(n_306) );
BUFx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g338 ( .A(n_234), .B(n_329), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_234), .B(n_271), .Y(n_357) );
AND2x4_ASAP7_75t_L g293 ( .A(n_235), .B(n_267), .Y(n_293) );
AND2x2_ASAP7_75t_L g431 ( .A(n_235), .B(n_407), .Y(n_431) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_242), .Y(n_235) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_236), .Y(n_260) );
INVx1_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
INVx1_ASAP7_75t_L g370 ( .A(n_236), .Y(n_370) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_239), .Y(n_471) );
INVx2_ASAP7_75t_L g539 ( .A(n_239), .Y(n_539) );
INVx1_ASAP7_75t_L g516 ( .A(n_241), .Y(n_516) );
OR2x2_ASAP7_75t_L g261 ( .A(n_242), .B(n_246), .Y(n_261) );
AND2x2_ASAP7_75t_L g270 ( .A(n_242), .B(n_271), .Y(n_270) );
NOR2xp67_ASAP7_75t_L g290 ( .A(n_242), .B(n_291), .Y(n_290) );
OAI221xp5_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .B1(n_259), .B2(n_262), .C(n_266), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_245), .A2(n_267), .B(n_269), .C(n_272), .Y(n_266) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_246), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_SL g374 ( .A(n_246), .B(n_268), .Y(n_374) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_246), .Y(n_381) );
AND2x2_ASAP7_75t_L g299 ( .A(n_247), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g336 ( .A(n_247), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_258), .Y(n_248) );
INVx2_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
AOI222xp33_ASAP7_75t_L g376 ( .A1(n_249), .A2(n_260), .B1(n_377), .B2(n_379), .C1(n_380), .C2(n_382), .Y(n_376) );
AND2x2_ASAP7_75t_L g433 ( .A(n_249), .B(n_402), .Y(n_433) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_257), .Y(n_249) );
INVx1_ASAP7_75t_L g323 ( .A(n_250), .Y(n_323) );
AO21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_255), .Y(n_250) );
INVx3_ASAP7_75t_L g486 ( .A(n_251), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_251), .B(n_506), .Y(n_505) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_251), .A2(n_522), .B(n_529), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_251), .B(n_530), .Y(n_529) );
AO21x2_ASAP7_75t_L g544 ( .A1(n_251), .A2(n_545), .B(n_552), .Y(n_544) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x4_ASAP7_75t_L g275 ( .A(n_256), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g361 ( .A(n_258), .B(n_295), .Y(n_361) );
AOI21xp33_ASAP7_75t_L g372 ( .A1(n_259), .A2(n_373), .B(n_375), .Y(n_372) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g300 ( .A(n_260), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_260), .B(n_267), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_260), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
INVx3_ASAP7_75t_L g326 ( .A(n_264), .Y(n_326) );
OR2x2_ASAP7_75t_L g378 ( .A(n_264), .B(n_300), .Y(n_378) );
AND2x2_ASAP7_75t_L g294 ( .A(n_265), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g332 ( .A(n_265), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_265), .B(n_326), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_265), .B(n_322), .Y(n_348) );
AND2x2_ASAP7_75t_L g352 ( .A(n_265), .B(n_334), .Y(n_352) );
INVxp67_ASAP7_75t_L g284 ( .A(n_267), .Y(n_284) );
BUFx3_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_269), .A2(n_342), .B1(n_347), .B2(n_348), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_269), .B(n_374), .Y(n_404) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g390 ( .A(n_270), .B(n_381), .Y(n_390) );
AND2x2_ASAP7_75t_L g419 ( .A(n_270), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g424 ( .A(n_270), .B(n_374), .Y(n_424) );
INVx1_ASAP7_75t_L g337 ( .A(n_271), .Y(n_337) );
BUFx2_ASAP7_75t_L g343 ( .A(n_271), .Y(n_343) );
INVx1_ASAP7_75t_L g428 ( .A(n_272), .Y(n_428) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_273), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g304 ( .A(n_274), .Y(n_304) );
NOR2x1_ASAP7_75t_L g280 ( .A(n_275), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_275), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
INVx3_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
OR2x2_ASAP7_75t_L g400 ( .A(n_275), .B(n_401), .Y(n_400) );
AOI211xp5_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_282), .B(n_285), .C(n_297), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_278), .A2(n_415), .B1(n_422), .B2(n_424), .C(n_425), .Y(n_414) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_286), .B(n_292), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_289), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_288), .B(n_326), .Y(n_340) );
AND2x2_ASAP7_75t_L g382 ( .A(n_288), .B(n_322), .Y(n_382) );
INVx1_ASAP7_75t_SL g395 ( .A(n_289), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_289), .B(n_343), .Y(n_398) );
INVx1_ASAP7_75t_L g416 ( .A(n_290), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
AOI221xp5_ASAP7_75t_L g383 ( .A1(n_294), .A2(n_384), .B1(n_386), .B2(n_390), .C(n_391), .Y(n_383) );
AND2x2_ASAP7_75t_L g410 ( .A(n_295), .B(n_402), .Y(n_410) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g394 ( .A(n_296), .Y(n_394) );
AOI21xp33_ASAP7_75t_SL g297 ( .A1(n_298), .A2(n_301), .B(n_302), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g365 ( .A(n_300), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g351 ( .A(n_301), .Y(n_351) );
INVx1_ASAP7_75t_L g379 ( .A(n_302), .Y(n_379) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
O2A1O1Ixp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_310), .C(n_313), .Y(n_305) );
OAI31xp33_ASAP7_75t_L g432 ( .A1(n_306), .A2(n_344), .A3(n_431), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g406 ( .A(n_309), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_SL g427 ( .A(n_309), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_311), .B(n_326), .Y(n_354) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g429 ( .A(n_312), .B(n_326), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_321), .B1(n_325), .B2(n_328), .Y(n_316) );
NAND2xp33_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_320), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g359 ( .A(n_320), .B(n_343), .Y(n_359) );
AND2x2_ASAP7_75t_L g413 ( .A(n_320), .B(n_408), .Y(n_413) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_324), .Y(n_321) );
INVx1_ASAP7_75t_L g388 ( .A(n_324), .Y(n_388) );
NOR2xp67_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI32xp33_ASAP7_75t_L g391 ( .A1(n_326), .A2(n_360), .A3(n_392), .B1(n_394), .B2(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g366 ( .A(n_329), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_329), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g389 ( .A(n_333), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_338), .B(n_339), .C(n_341), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_337), .B(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g349 ( .A1(n_338), .A2(n_350), .B1(n_351), .B2(n_352), .C(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g350 ( .A(n_348), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_355), .B1(n_358), .B2(n_360), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_SL g415 ( .A(n_358), .B(n_416), .C(n_417), .D(n_418), .Y(n_415) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NAND4xp25_ASAP7_75t_SL g362 ( .A(n_363), .B(n_376), .C(n_383), .D(n_396), .Y(n_362) );
O2A1O1Ixp33_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_367), .B(n_371), .C(n_372), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_SL g393 ( .A(n_369), .Y(n_393) );
INVx2_ASAP7_75t_L g417 ( .A(n_374), .Y(n_417) );
OR2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_397), .A2(n_399), .B(n_403), .Y(n_396) );
INVxp67_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g422 ( .A(n_402), .B(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_SL g403 ( .A1(n_404), .A2(n_405), .B(n_409), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
CKINVDCx16_ASAP7_75t_R g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_425) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND3xp33_ASAP7_75t_SL g438 ( .A(n_434), .B(n_439), .C(n_441), .Y(n_438) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVxp67_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_446), .B1(n_448), .B2(n_452), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g751 ( .A(n_444), .Y(n_751) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g752 ( .A(n_446), .Y(n_752) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g753 ( .A(n_449), .Y(n_753) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g754 ( .A(n_452), .Y(n_754) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
OR5x1_ASAP7_75t_L g453 ( .A(n_454), .B(n_623), .C(n_701), .D(n_725), .E(n_742), .Y(n_453) );
OAI211xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_495), .B(n_541), .C(n_600), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_475), .Y(n_455) );
AND2x2_ASAP7_75t_L g554 ( .A(n_456), .B(n_477), .Y(n_554) );
INVx5_ASAP7_75t_SL g582 ( .A(n_456), .Y(n_582) );
AND2x2_ASAP7_75t_L g618 ( .A(n_456), .B(n_603), .Y(n_618) );
OR2x2_ASAP7_75t_L g657 ( .A(n_456), .B(n_476), .Y(n_657) );
OR2x2_ASAP7_75t_L g688 ( .A(n_456), .B(n_579), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g724 ( .A(n_456), .B(n_592), .Y(n_724) );
AND2x2_ASAP7_75t_L g736 ( .A(n_456), .B(n_579), .Y(n_736) );
OR2x6_ASAP7_75t_L g456 ( .A(n_457), .B(n_474), .Y(n_456) );
BUFx2_ASAP7_75t_L g511 ( .A(n_459), .Y(n_511) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_463), .A2(n_473), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_463), .A2(n_473), .B(n_534), .C(n_535), .Y(n_533) );
INVx5_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B(n_470), .C(n_471), .Y(n_466) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_468), .A2(n_471), .B(n_503), .C(n_504), .Y(n_502) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g735 ( .A(n_475), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_L g598 ( .A(n_476), .B(n_599), .Y(n_598) );
OR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_487), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_477), .B(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_477), .Y(n_591) );
INVx3_ASAP7_75t_L g606 ( .A(n_477), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_477), .B(n_487), .Y(n_630) );
OR2x2_ASAP7_75t_L g639 ( .A(n_477), .B(n_582), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_477), .B(n_603), .Y(n_643) );
AND2x2_ASAP7_75t_L g649 ( .A(n_477), .B(n_650), .Y(n_649) );
INVxp67_ASAP7_75t_L g686 ( .A(n_477), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_477), .B(n_544), .Y(n_700) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_485), .Y(n_477) );
OA21x2_ASAP7_75t_L g531 ( .A1(n_486), .A2(n_532), .B(n_540), .Y(n_531) );
OR2x2_ASAP7_75t_L g592 ( .A(n_487), .B(n_544), .Y(n_592) );
AND2x2_ASAP7_75t_L g603 ( .A(n_487), .B(n_579), .Y(n_603) );
AND2x2_ASAP7_75t_L g615 ( .A(n_487), .B(n_606), .Y(n_615) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_487), .B(n_544), .Y(n_638) );
INVx1_ASAP7_75t_SL g650 ( .A(n_487), .Y(n_650) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g543 ( .A(n_488), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_488), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_507), .Y(n_496) );
AND2x2_ASAP7_75t_L g563 ( .A(n_497), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_497), .B(n_520), .Y(n_567) );
AND2x2_ASAP7_75t_L g570 ( .A(n_497), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_497), .B(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g595 ( .A(n_497), .B(n_586), .Y(n_595) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_497), .Y(n_614) );
AND2x2_ASAP7_75t_L g635 ( .A(n_497), .B(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g645 ( .A(n_497), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g691 ( .A(n_497), .B(n_574), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_497), .B(n_597), .Y(n_718) );
INVx5_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g588 ( .A(n_498), .Y(n_588) );
AND2x2_ASAP7_75t_L g654 ( .A(n_498), .B(n_586), .Y(n_654) );
AND2x2_ASAP7_75t_L g738 ( .A(n_498), .B(n_606), .Y(n_738) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_507), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_507), .Y(n_727) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_520), .Y(n_507) );
AND2x2_ASAP7_75t_L g557 ( .A(n_508), .B(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g566 ( .A(n_508), .B(n_564), .Y(n_566) );
INVx5_ASAP7_75t_L g574 ( .A(n_508), .Y(n_574) );
AND2x2_ASAP7_75t_L g597 ( .A(n_508), .B(n_531), .Y(n_597) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_508), .Y(n_634) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AOI21xp5_ASAP7_75t_SL g509 ( .A1(n_510), .A2(n_512), .B(n_516), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
INVx1_ASAP7_75t_L g675 ( .A(n_520), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_520), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g708 ( .A(n_520), .B(n_574), .Y(n_708) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_520), .A2(n_631), .B(n_738), .C(n_739), .Y(n_737) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_531), .Y(n_520) );
BUFx2_ASAP7_75t_L g558 ( .A(n_521), .Y(n_558) );
INVx2_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_528), .Y(n_522) );
INVx2_ASAP7_75t_L g564 ( .A(n_531), .Y(n_564) );
AND2x2_ASAP7_75t_L g571 ( .A(n_531), .B(n_562), .Y(n_571) );
AND2x2_ASAP7_75t_L g662 ( .A(n_531), .B(n_574), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
AOI211x1_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_555), .B(n_568), .C(n_593), .Y(n_541) );
INVx1_ASAP7_75t_L g659 ( .A(n_542), .Y(n_659) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_554), .Y(n_542) );
INVx5_ASAP7_75t_SL g579 ( .A(n_544), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_544), .B(n_649), .Y(n_648) );
AOI311xp33_ASAP7_75t_L g667 ( .A1(n_544), .A2(n_668), .A3(n_670), .B(n_671), .C(n_677), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_544), .A2(n_615), .B(n_703), .C(n_706), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
INVxp67_ASAP7_75t_L g622 ( .A(n_554), .Y(n_622) );
NAND4xp25_ASAP7_75t_SL g555 ( .A(n_556), .B(n_559), .C(n_565), .D(n_567), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_556), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g613 ( .A(n_557), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_563), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_560), .B(n_566), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_560), .B(n_573), .Y(n_693) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_561), .B(n_574), .Y(n_711) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g586 ( .A(n_562), .Y(n_586) );
INVxp67_ASAP7_75t_L g621 ( .A(n_563), .Y(n_621) );
AND2x4_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g647 ( .A(n_564), .B(n_586), .Y(n_647) );
INVx1_ASAP7_75t_L g674 ( .A(n_564), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_564), .B(n_661), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_565), .B(n_635), .Y(n_655) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_566), .B(n_588), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_566), .B(n_635), .Y(n_734) );
INVx1_ASAP7_75t_L g745 ( .A(n_567), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .B(n_575), .C(n_583), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g587 ( .A(n_571), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g625 ( .A(n_571), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g607 ( .A(n_572), .Y(n_607) );
AND2x2_ASAP7_75t_L g584 ( .A(n_573), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_573), .B(n_635), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_573), .B(n_654), .Y(n_678) );
OR2x2_ASAP7_75t_L g594 ( .A(n_574), .B(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g626 ( .A(n_574), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_574), .B(n_586), .Y(n_641) );
AND2x2_ASAP7_75t_L g698 ( .A(n_574), .B(n_654), .Y(n_698) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_574), .Y(n_705) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g709 ( .A1(n_576), .A2(n_588), .B1(n_710), .B2(n_712), .C(n_715), .Y(n_709) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g599 ( .A(n_579), .B(n_582), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_579), .B(n_649), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_579), .B(n_606), .Y(n_714) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g699 ( .A(n_581), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g713 ( .A(n_581), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_582), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_582), .B(n_603), .Y(n_610) );
AND2x2_ASAP7_75t_L g680 ( .A(n_582), .B(n_681), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_582), .B(n_629), .Y(n_726) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_582), .B(n_730), .Y(n_729) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_587), .B(n_589), .Y(n_583) );
INVx2_ASAP7_75t_L g616 ( .A(n_584), .Y(n_616) );
HB1xp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g636 ( .A(n_586), .Y(n_636) );
OR2x2_ASAP7_75t_L g640 ( .A(n_588), .B(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g743 ( .A(n_588), .B(n_711), .Y(n_743) );
INVx1_ASAP7_75t_SL g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AOI21xp33_ASAP7_75t_SL g593 ( .A1(n_594), .A2(n_596), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g747 ( .A(n_594), .Y(n_747) );
INVx2_ASAP7_75t_SL g661 ( .A(n_595), .Y(n_661) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
A2O1A1Ixp33_ASAP7_75t_L g742 ( .A1(n_598), .A2(n_679), .B(n_743), .C(n_744), .Y(n_742) );
OAI322xp33_ASAP7_75t_SL g611 ( .A1(n_599), .A2(n_612), .A3(n_615), .B1(n_616), .B2(n_617), .C1(n_619), .C2(n_622), .Y(n_611) );
INVx2_ASAP7_75t_L g631 ( .A(n_599), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_607), .B1(n_608), .B2(n_610), .C(n_611), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
OAI22xp33_ASAP7_75t_SL g677 ( .A1(n_602), .A2(n_678), .B1(n_679), .B2(n_682), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_603), .B(n_606), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_603), .B(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g676 ( .A(n_605), .B(n_638), .Y(n_676) );
INVx1_ASAP7_75t_L g666 ( .A(n_606), .Y(n_666) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_610), .A2(n_720), .B(n_722), .Y(n_719) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_612), .A2(n_645), .B(n_648), .Y(n_644) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp67_ASAP7_75t_SL g673 ( .A(n_614), .B(n_674), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_614), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g730 ( .A(n_615), .Y(n_730) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_624), .B(n_651), .C(n_667), .D(n_683), .Y(n_623) );
AOI211xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_627), .B(n_632), .C(n_644), .Y(n_624) );
INVx1_ASAP7_75t_L g716 ( .A(n_625), .Y(n_716) );
AND2x2_ASAP7_75t_L g664 ( .A(n_626), .B(n_647), .Y(n_664) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_631), .B(n_666), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_640), .B2(n_642), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_634), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g682 ( .A(n_635), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g696 ( .A1(n_635), .A2(n_674), .B(n_697), .C(n_699), .Y(n_696) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g681 ( .A(n_638), .Y(n_681) );
INVx1_ASAP7_75t_L g741 ( .A(n_639), .Y(n_741) );
NAND2xp33_ASAP7_75t_SL g731 ( .A(n_640), .B(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g670 ( .A(n_649), .Y(n_670) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_655), .B(n_656), .C(n_658), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_660), .B1(n_663), .B2(n_665), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_661), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_666), .B(n_687), .Y(n_749) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_SL g671 ( .A1(n_672), .A2(n_675), .B(n_676), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_689), .B1(n_692), .B2(n_694), .C(n_696), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVxp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_699), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g701 ( .A(n_702), .B(n_709), .C(n_719), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx16_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B(n_728), .C(n_737), .Y(n_725) );
INVx1_ASAP7_75t_L g746 ( .A(n_726), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_733), .B2(n_735), .Y(n_728) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g744 ( .A1(n_745), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
OAI22x1_ASAP7_75t_SL g750 ( .A1(n_751), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_758), .Y(n_757) );
endmodule