module fake_jpeg_26865_n_129 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_129);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx4f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_5),
.B(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_64),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_41),
.B1(n_47),
.B2(n_52),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_69),
.B1(n_57),
.B2(n_53),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_63),
.A2(n_59),
.B1(n_49),
.B2(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_75),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_77),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_43),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_0),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_54),
.C(n_51),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_5),
.C(n_6),
.Y(n_96)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_1),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_1),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_91),
.B1(n_93),
.B2(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_2),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_90),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_3),
.C(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_4),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_29),
.B1(n_39),
.B2(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_102),
.B1(n_104),
.B2(n_92),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_23),
.B1(n_37),
.B2(n_36),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_106),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_86),
.C(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_86),
.Y(n_107)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_112),
.B(n_101),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_98),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_115),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_101),
.A3(n_96),
.B1(n_16),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AOI322xp5_ASAP7_75t_L g122 ( 
.A1(n_120),
.A2(n_121),
.A3(n_113),
.B1(n_108),
.B2(n_112),
.C1(n_117),
.C2(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_122),
.A2(n_119),
.B(n_118),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_124),
.B(n_13),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_30),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_40),
.C(n_7),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_6),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_8),
.Y(n_129)
);


endmodule