module real_jpeg_32661_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx3_ASAP7_75t_L g119 ( 
.A(n_0),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_0),
.Y(n_185)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_0),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_1),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_1),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_1),
.A2(n_141),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_1),
.A2(n_141),
.B1(n_517),
.B2(n_519),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_2),
.A2(n_121),
.B1(n_122),
.B2(n_127),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_2),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_2),
.A2(n_121),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

AO22x1_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_177),
.B1(n_179),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_3),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_4),
.A2(n_237),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_4),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_4),
.A2(n_240),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_4),
.A2(n_240),
.B1(n_312),
.B2(n_315),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_6),
.Y(n_86)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_7),
.Y(n_178)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_7),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_8),
.A2(n_60),
.B1(n_291),
.B2(n_295),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_8),
.A2(n_60),
.B1(n_381),
.B2(n_383),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_8),
.A2(n_60),
.B1(n_435),
.B2(n_439),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_9),
.B(n_36),
.Y(n_158)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_9),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_9),
.B(n_67),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_9),
.A2(n_284),
.B1(n_402),
.B2(n_405),
.Y(n_401)
);

OAI32xp33_ASAP7_75t_L g409 ( 
.A1(n_9),
.A2(n_341),
.A3(n_410),
.B1(n_413),
.B2(n_420),
.Y(n_409)
);

OAI21xp33_ASAP7_75t_L g450 ( 
.A1(n_9),
.A2(n_174),
.B(n_370),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_10),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_10),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_10),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_12),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_13),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_13),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_14),
.A2(n_169),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_14),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_14),
.A2(n_173),
.B1(n_395),
.B2(n_506),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_15),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_15),
.A2(n_76),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_15),
.A2(n_76),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_15),
.A2(n_76),
.B1(n_395),
.B2(n_398),
.Y(n_394)
);

OAI22x1_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_16),
.A2(n_52),
.B1(n_110),
.B2(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_16),
.A2(n_52),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_16),
.A2(n_52),
.B1(n_373),
.B2(n_374),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_491),
.Y(n_17)
);

OAI21x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_323),
.B(n_487),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI21xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_260),
.B(n_300),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_21),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_165),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_22),
.B(n_166),
.C(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_68),
.C(n_115),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_23),
.A2(n_24),
.B1(n_69),
.B2(n_70),
.Y(n_264)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_58),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_49),
.Y(n_25)
);

AO22x1_ASAP7_75t_L g253 ( 
.A1(n_26),
.A2(n_59),
.B1(n_67),
.B2(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_26),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_26),
.B(n_254),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

AOI22x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_27)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_28),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_31),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_31),
.Y(n_164)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_34),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_40),
.B1(n_43),
.B2(n_47),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_49),
.B(n_67),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_57),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_57),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_66),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_79),
.B(n_106),
.Y(n_70)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_71),
.Y(n_288)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_75),
.Y(n_294)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g245 ( 
.A1(n_79),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_245)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_79),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g400 ( 
.A1(n_79),
.A2(n_106),
.B(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_80),
.B(n_109),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_80),
.A2(n_107),
.B1(n_249),
.B2(n_516),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_93),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_87),
.B2(n_91),
.Y(n_81)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_87),
.B1(n_91),
.B2(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_83),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_83),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_83),
.Y(n_397)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_83),
.Y(n_508)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_86),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_90),
.Y(n_217)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_97),
.B1(n_100),
.B2(n_105),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_96),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_96),
.Y(n_299)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.Y(n_106)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_107),
.Y(n_247)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_109),
.Y(n_246)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_112),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g519 ( 
.A(n_112),
.Y(n_519)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_113),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_115),
.A2(n_116),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_144),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_117),
.A2(n_144),
.B1(n_145),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_117),
.Y(n_307)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_131),
.B2(n_136),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_118),
.A2(n_131),
.B1(n_433),
.B2(n_441),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_120),
.Y(n_230)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_125),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_126),
.Y(n_140)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_126),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_126),
.Y(n_376)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_130),
.Y(n_317)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_131),
.B(n_372),
.Y(n_428)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_131),
.A2(n_176),
.B(n_503),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g427 ( 
.A(n_135),
.Y(n_427)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_137),
.A2(n_174),
.B1(n_231),
.B2(n_311),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_140),
.Y(n_458)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

AOI32xp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_149),
.A3(n_154),
.B1(n_158),
.B2(n_159),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_158),
.Y(n_285)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_227),
.Y(n_165)
);

XOR2x2_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_186),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_167),
.B(n_187),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_174),
.B1(n_175),
.B2(n_183),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_174),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_169),
.Y(n_344)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_174),
.A2(n_362),
.B(n_370),
.Y(n_361)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_178),
.Y(n_205)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_178),
.Y(n_334)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g371 ( 
.A(n_183),
.Y(n_371)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_185),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_211),
.B1(n_218),
.B2(n_225),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_188),
.A2(n_211),
.B1(n_225),
.B2(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g270 ( 
.A(n_188),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g393 ( 
.A1(n_188),
.A2(n_225),
.B1(n_380),
.B2(n_394),
.Y(n_393)
);

OAI21xp33_ASAP7_75t_SL g470 ( 
.A1(n_188),
.A2(n_353),
.B(n_394),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_188),
.A2(n_218),
.B1(n_225),
.B2(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_203),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_192),
.B1(n_196),
.B2(n_199),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

OAI22x1_ASAP7_75t_L g203 ( 
.A1(n_196),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_202),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_217),
.Y(n_382)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_223),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_224),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_224),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_225),
.A2(n_380),
.B(n_385),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_225),
.B(n_284),
.Y(n_445)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_226),
.A2(n_270),
.B1(n_271),
.B2(n_277),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_226),
.B(n_271),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_227),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_244),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_228),
.B(n_245),
.C(n_253),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_229),
.B(n_235),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx2_ASAP7_75t_R g503 ( 
.A(n_234),
.Y(n_503)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_239),
.Y(n_276)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_253),
.Y(n_244)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_247),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_247),
.B(n_284),
.Y(n_378)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_261),
.B(n_489),
.C(n_490),
.Y(n_488)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_262),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_302)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_278),
.C(n_286),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_286),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_270),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_270),
.B(n_271),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_279),
.B(n_514),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_282),
.A2(n_284),
.B(n_285),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_284),
.B(n_341),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g355 ( 
.A1(n_284),
.A2(n_340),
.B(n_356),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_284),
.B(n_421),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_284),
.B(n_453),
.Y(n_452)
);

AOI22x1_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_290),
.Y(n_321)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_298),
.Y(n_412)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_301),
.B(n_303),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_308),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_304),
.B(n_481),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_306),
.A2(n_308),
.B1(n_309),
.B2(n_482),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_306),
.Y(n_482)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_318),
.C(n_320),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_310),
.A2(n_318),
.B1(n_319),
.B2(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_310),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_311),
.A2(n_425),
.B(n_428),
.Y(n_424)
);

BUFx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_317),
.Y(n_440)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_320),
.B(n_466),
.Y(n_465)
);

AOI31xp67_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_474),
.A3(n_483),
.B(n_484),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

AOI211x1_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_429),
.B(n_461),
.C(n_463),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_386),
.B(n_387),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_327),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_360),
.Y(n_327)
);

NOR2x1_ASAP7_75t_SL g386 ( 
.A(n_328),
.B(n_360),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_352),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_329),
.B(n_352),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_339),
.B1(n_343),
.B2(n_345),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_331),
.Y(n_363)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_338),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g423 ( 
.A(n_342),
.Y(n_423)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_349),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_377),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_361),
.B(n_389),
.C(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx6_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_391),
.Y(n_387)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_388),
.B(n_391),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_408),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_393),
.B(n_408),
.C(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_400),
.Y(n_473)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx5_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_409),
.B(n_424),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_409),
.B(n_424),
.Y(n_471)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx2_ASAP7_75t_SL g411 ( 
.A(n_412),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_416),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_SL g421 ( 
.A(n_422),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_426),
.Y(n_425)
);

INVx5_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_428),
.A2(n_434),
.B(n_447),
.Y(n_446)
);

AOI21xp33_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_443),
.B(n_460),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_442),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_442),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

BUFx2_ASAP7_75t_SL g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_449),
.B(n_459),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_445),
.B(n_446),
.Y(n_459)
);

INVx8_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx5_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_472),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_464),
.B(n_472),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_465),
.B(n_469),
.C(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_471),
.Y(n_479)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_480),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_478),
.B(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_480),
.Y(n_486)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_488),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_523),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_496),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_494),
.B(n_496),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_500),
.B1(n_510),
.B2(n_522),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_502),
.B1(n_504),
.B2(n_509),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_504),
.Y(n_509)
);

BUFx4f_ASAP7_75t_SL g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_515),
.B1(n_520),
.B2(n_521),
.Y(n_512)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_513),
.Y(n_521)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_515),
.Y(n_520)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);


endmodule