module fake_jpeg_19715_n_326 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_326);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_41),
.Y(n_57)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_24),
.B1(n_21),
.B2(n_29),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_58),
.B1(n_32),
.B2(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_49),
.B(n_25),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_23),
.C(n_20),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_51),
.B(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_21),
.B1(n_29),
.B2(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_43),
.B(n_20),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_36),
.Y(n_78)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_33),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_29),
.B1(n_19),
.B2(n_38),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_74),
.B1(n_50),
.B2(n_31),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_76),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_56),
.A2(n_19),
.B1(n_39),
.B2(n_33),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_27),
.B1(n_25),
.B2(n_32),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_75),
.B1(n_83),
.B2(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_89),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_45),
.A2(n_19),
.B1(n_30),
.B2(n_28),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_51),
.B(n_43),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_78),
.B(n_48),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_45),
.A2(n_36),
.B1(n_31),
.B2(n_28),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_48),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_61),
.A2(n_27),
.B(n_31),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_88),
.B1(n_95),
.B2(n_63),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_52),
.A2(n_31),
.B1(n_16),
.B2(n_18),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_46),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_91),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_92),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_20),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_71),
.B(n_60),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_107),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_101),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_59),
.B1(n_50),
.B2(n_17),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_110),
.B1(n_114),
.B2(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_48),
.C(n_62),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_85),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_113),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_17),
.B1(n_20),
.B2(n_18),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_18),
.B1(n_15),
.B2(n_12),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_66),
.B1(n_73),
.B2(n_81),
.Y(n_134)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_22),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_74),
.A2(n_22),
.B1(n_62),
.B2(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_119),
.B(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_135),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_136),
.Y(n_159)
);

INVxp67_ASAP7_75t_SL g129 ( 
.A(n_124),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_78),
.B(n_90),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_130),
.A2(n_140),
.B(n_145),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_134),
.A2(n_144),
.B1(n_154),
.B2(n_122),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_104),
.B(n_81),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_113),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_124),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_143),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_89),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_91),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_92),
.B1(n_94),
.B2(n_87),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_75),
.B(n_82),
.C(n_68),
.D(n_69),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_69),
.B1(n_79),
.B2(n_87),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_79),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_149),
.Y(n_169)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_150),
.Y(n_170)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_153),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_79),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_112),
.A2(n_95),
.B1(n_93),
.B2(n_22),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_95),
.B1(n_15),
.B2(n_12),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_115),
.B1(n_123),
.B2(n_108),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_105),
.B(n_102),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_157),
.A2(n_176),
.B1(n_179),
.B2(n_187),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_120),
.B(n_114),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_175),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_109),
.C(n_121),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_146),
.C(n_155),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_123),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_166),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_140),
.A2(n_120),
.B(n_103),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_171),
.B(n_174),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_165),
.A2(n_185),
.B1(n_153),
.B2(n_151),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_132),
.Y(n_166)
);

AO22x1_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_120),
.B1(n_106),
.B2(n_123),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_178),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_117),
.B(n_108),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_137),
.A2(n_118),
.B1(n_15),
.B2(n_12),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_97),
.B1(n_11),
.B2(n_10),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_145),
.B(n_126),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_11),
.B1(n_10),
.B2(n_2),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_62),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_11),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_6),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_150),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_131),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_0),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_131),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_125),
.A2(n_139),
.B1(n_142),
.B2(n_136),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_189),
.A2(n_148),
.B1(n_3),
.B2(n_4),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_125),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_6),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_201),
.C(n_213),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_192),
.A2(n_208),
.B1(n_187),
.B2(n_176),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_196),
.A2(n_156),
.B(n_188),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_162),
.B(n_148),
.C(n_3),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_185),
.B1(n_165),
.B2(n_182),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_159),
.Y(n_207)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_169),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_9),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_7),
.C(n_170),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_4),
.C(n_5),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_214),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_216),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_6),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_6),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_166),
.B(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_7),
.C(n_161),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_167),
.C(n_178),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_230),
.B(n_194),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_221),
.A2(n_239),
.B1(n_205),
.B2(n_206),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_225),
.B1(n_217),
.B2(n_215),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_188),
.B1(n_178),
.B2(n_167),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_229),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_161),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_236),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_198),
.A2(n_164),
.B(n_171),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_178),
.C(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_233),
.C(n_235),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_7),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_219),
.C(n_196),
.Y(n_233)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_160),
.C(n_182),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_192),
.A2(n_183),
.B1(n_172),
.B2(n_175),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_170),
.C(n_177),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_195),
.C(n_206),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_257),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_249),
.A2(n_235),
.B(n_233),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_197),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_262),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_238),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_237),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_253),
.C(n_256),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_218),
.C(n_210),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_205),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_202),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_199),
.C(n_200),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_223),
.A2(n_211),
.B1(n_194),
.B2(n_199),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_234),
.A2(n_200),
.B1(n_213),
.B2(n_214),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_260),
.B(n_244),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_228),
.B1(n_243),
.B2(n_225),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_7),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_261),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_236),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_220),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_268),
.B(n_256),
.Y(n_281)
);

INVx13_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_272),
.B(n_247),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_268),
.B(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_278),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_248),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g279 ( 
.A(n_253),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_292),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_267),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_294),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_285),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_284),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_263),
.B(n_264),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_291),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_271),
.A2(n_246),
.B(n_262),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_289),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_246),
.C(n_247),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_250),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_293),
.A2(n_265),
.B(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_222),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_265),
.B1(n_272),
.B2(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_295),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_270),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_269),
.B1(n_222),
.B2(n_266),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_291),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_305),
.B(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_312),
.Y(n_318)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_296),
.A2(n_288),
.B(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_313),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_288),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_303),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_304),
.C(n_299),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_303),
.Y(n_315)
);

AOI21x1_ASAP7_75t_SL g313 ( 
.A1(n_302),
.A2(n_298),
.B(n_297),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_318),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_316),
.B(n_308),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_320),
.B(n_321),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_314),
.A2(n_311),
.B(n_313),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_322),
.Y(n_323)
);

OAI21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_317),
.B(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_317),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_318),
.Y(n_326)
);


endmodule