module fake_jpeg_5355_n_252 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_252);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_252;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_18),
.B(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_21),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_24),
.B1(n_29),
.B2(n_26),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_18),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_49),
.B(n_60),
.Y(n_69)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_32),
.A2(n_30),
.B1(n_19),
.B2(n_28),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_47),
.A2(n_55),
.B1(n_61),
.B2(n_21),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_25),
.B1(n_29),
.B2(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_32),
.A2(n_19),
.B1(n_28),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_84)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_23),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_16),
.B1(n_29),
.B2(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_40),
.B(n_42),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_70),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_45),
.B1(n_60),
.B2(n_49),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_40),
.B1(n_24),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_75),
.B1(n_79),
.B2(n_83),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_31),
.B1(n_16),
.B2(n_15),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_63),
.B1(n_50),
.B2(n_44),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_37),
.B1(n_21),
.B2(n_16),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_62),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_22),
.B1(n_30),
.B2(n_28),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_53),
.B1(n_43),
.B2(n_54),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_67),
.B(n_46),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_89),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g87 ( 
.A1(n_68),
.A2(n_43),
.B1(n_60),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_82),
.B1(n_72),
.B2(n_3),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_66),
.B(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_30),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_46),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_90),
.A2(n_95),
.B1(n_100),
.B2(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_80),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_71),
.A2(n_64),
.B1(n_57),
.B2(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_3),
.B1(n_77),
.B2(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_70),
.B(n_65),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_84),
.A2(n_19),
.B1(n_22),
.B2(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_65),
.B(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_0),
.Y(n_104)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_76),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_4),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_36),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_81),
.B(n_82),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_73),
.B(n_81),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_109),
.B(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_106),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_116),
.B1(n_118),
.B2(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_1),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_117),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_77),
.C(n_82),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_87),
.C(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_93),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_103),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_87),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_2),
.B1(n_3),
.B2(n_77),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_98),
.B(n_101),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_92),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_86),
.B1(n_95),
.B2(n_100),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_113),
.B(n_125),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_131),
.A2(n_142),
.B(n_145),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_117),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_132),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_116),
.C(n_123),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_141),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_139),
.A2(n_110),
.B(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_89),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_106),
.B(n_104),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_146),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_114),
.A2(n_106),
.B(n_85),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_85),
.B1(n_92),
.B2(n_9),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_112),
.B(n_4),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_148),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_8),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_110),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_107),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_167),
.C(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_133),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_118),
.C(n_122),
.D(n_124),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_160),
.B(n_149),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_109),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_139),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_164),
.A2(n_171),
.B(n_154),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_147),
.B(n_119),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_128),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_121),
.B(n_119),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_121),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_135),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_170),
.A2(n_141),
.B1(n_144),
.B2(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_173),
.A2(n_176),
.B1(n_182),
.B2(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_174),
.B(n_157),
.C(n_168),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_146),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_175),
.B(n_179),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_144),
.B1(n_146),
.B2(n_131),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_165),
.B(n_136),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_142),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_184),
.B(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_158),
.B(n_143),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_165),
.C(n_172),
.D(n_163),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_167),
.A2(n_131),
.B1(n_138),
.B2(n_149),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_149),
.B1(n_129),
.B2(n_130),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_185),
.A2(n_159),
.B1(n_160),
.B2(n_157),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_148),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_166),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_193),
.B(n_174),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_171),
.B1(n_168),
.B2(n_172),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_196),
.A2(n_200),
.B1(n_126),
.B2(n_10),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_202),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_161),
.C(n_154),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_10),
.C(n_12),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_203),
.A2(n_9),
.B(n_10),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_206),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_155),
.B(n_126),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_189),
.B(n_175),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_92),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_205),
.A2(n_182),
.B1(n_180),
.B2(n_191),
.Y(n_207)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_207),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_201),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_218),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_190),
.B(n_179),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_209),
.A2(n_211),
.B(n_215),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_213),
.B(n_202),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_219),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_13),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_194),
.B(n_14),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_12),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_200),
.A2(n_12),
.B(n_13),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_229),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_219),
.B(n_198),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_222),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_192),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_192),
.Y(n_224)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_225),
.A2(n_13),
.B(n_14),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_234),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_231),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_213),
.B1(n_211),
.B2(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_195),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_228),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_212),
.B(n_218),
.C(n_228),
.D(n_236),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_227),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_208),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_242),
.B(n_212),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_243),
.A2(n_238),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_239),
.Y(n_245)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_245),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_248),
.B(n_244),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_233),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_249),
.Y(n_252)
);


endmodule