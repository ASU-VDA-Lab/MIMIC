module fake_jpeg_11173_n_519 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_519);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_519;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx5p33_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_59),
.Y(n_172)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_61),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_16),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_63),
.B(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_64),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_24),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_0),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_71),
.Y(n_128)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_24),
.B(n_12),
.CON(n_73),
.SN(n_73)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_73),
.B(n_38),
.Y(n_153)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_75),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_76),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_20),
.B(n_12),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_80),
.B(n_81),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_36),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_83),
.Y(n_147)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_84),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_22),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_85),
.B(n_88),
.Y(n_152)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_20),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_22),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_25),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_100),
.B(n_104),
.Y(n_166)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_35),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_103),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_23),
.B(n_1),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_48),
.Y(n_105)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_28),
.Y(n_107)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_108),
.Y(n_165)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_25),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_110),
.B(n_117),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_33),
.Y(n_111)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_33),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g141 ( 
.A(n_112),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_33),
.Y(n_113)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_38),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_39),
.Y(n_115)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_115),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_26),
.B(n_8),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_47),
.Y(n_118)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_47),
.Y(n_119)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_104),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_123),
.B(n_145),
.Y(n_239)
);

BUFx4f_ASAP7_75t_SL g129 ( 
.A(n_96),
.Y(n_129)
);

CKINVDCx9p33_ASAP7_75t_R g217 ( 
.A(n_129),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_85),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_144),
.B(n_151),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_80),
.B(n_26),
.Y(n_145)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_68),
.Y(n_150)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

NAND2xp33_ASAP7_75t_SL g209 ( 
.A(n_153),
.B(n_50),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_70),
.B(n_29),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_158),
.B(n_181),
.Y(n_253)
);

INVx11_ASAP7_75t_L g160 ( 
.A(n_74),
.Y(n_160)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_160),
.Y(n_226)
);

BUFx4f_ASAP7_75t_SL g168 ( 
.A(n_63),
.Y(n_168)
);

INVx13_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_31),
.B1(n_34),
.B2(n_19),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_170),
.B(n_56),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_92),
.B(n_29),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_56),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_75),
.A2(n_45),
.B1(n_31),
.B2(n_53),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_51),
.B1(n_53),
.B2(n_87),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_99),
.B(n_37),
.Y(n_181)
);

INVx11_ASAP7_75t_L g185 ( 
.A(n_76),
.Y(n_185)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_62),
.B(n_55),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_186),
.B(n_2),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_193),
.B(n_219),
.Y(n_284)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

INVx4_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_195),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_196),
.Y(n_268)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_143),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_197),
.Y(n_281)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_198),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_147),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_199),
.B(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_201),
.Y(n_259)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_203),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_206),
.A2(n_141),
.B1(n_213),
.B2(n_124),
.Y(n_275)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_207),
.Y(n_276)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_208),
.Y(n_282)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_209),
.A2(n_223),
.B(n_242),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_140),
.Y(n_210)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_210),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_211),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_186),
.A2(n_66),
.B1(n_64),
.B2(n_112),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g213 ( 
.A1(n_180),
.A2(n_113),
.B1(n_111),
.B2(n_45),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_162),
.A2(n_171),
.B1(n_179),
.B2(n_190),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_216),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_121),
.A2(n_48),
.B1(n_34),
.B2(n_19),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_218),
.A2(n_236),
.B1(n_245),
.B2(n_256),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_55),
.Y(n_219)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_220),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_142),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_221),
.B(n_227),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_155),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_235),
.Y(n_262)
);

OR2x4_ASAP7_75t_L g223 ( 
.A(n_152),
.B(n_166),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_224),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_142),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_169),
.B(n_50),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_228),
.B(n_240),
.Y(n_296)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_234),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_232),
.A2(n_175),
.B1(n_141),
.B2(n_137),
.Y(n_264)
);

CKINVDCx12_ASAP7_75t_R g233 ( 
.A(n_129),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_233),
.Y(n_269)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_188),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_148),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_49),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_133),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_241),
.B(n_247),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_49),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_250),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_154),
.A2(n_18),
.B1(n_37),
.B2(n_5),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g287 ( 
.A1(n_246),
.A2(n_131),
.B1(n_120),
.B2(n_146),
.Y(n_287)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_148),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_254),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_126),
.B(n_18),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_251),
.B(n_252),
.Y(n_288)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_132),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_126),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_255),
.B(n_132),
.Y(n_300)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_189),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_217),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_263),
.B(n_302),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_264),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_136),
.B1(n_164),
.B2(n_135),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_270),
.A2(n_275),
.B1(n_286),
.B2(n_304),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_166),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_278),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_152),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_191),
.B(n_172),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_279),
.A2(n_280),
.B(n_294),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_139),
.B(n_128),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_212),
.A2(n_163),
.B1(n_146),
.B2(n_122),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_287),
.B(n_295),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_242),
.A2(n_138),
.B(n_161),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_222),
.B(n_161),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_246),
.B(n_122),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_256),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_300),
.B(n_127),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_215),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_203),
.A2(n_163),
.B1(n_167),
.B2(n_7),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_225),
.B(n_11),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_305),
.B(n_200),
.Y(n_311)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_238),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_309),
.B(n_311),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_291),
.A2(n_234),
.B1(n_208),
.B2(n_205),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_310),
.A2(n_326),
.B1(n_265),
.B2(n_282),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_SL g349 ( 
.A1(n_312),
.A2(n_301),
.B(n_290),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_278),
.B(n_200),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_313),
.B(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_259),
.Y(n_314)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

AND2x6_ASAP7_75t_L g315 ( 
.A(n_261),
.B(n_127),
.Y(n_315)
);

AND2x6_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_294),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_316),
.B(n_320),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_285),
.B(n_196),
.C(n_210),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_319),
.C(n_334),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_236),
.C(n_211),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_260),
.B(n_231),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_226),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_321),
.Y(n_368)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_259),
.Y(n_322)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_274),
.B(n_231),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_324),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_271),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_329),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_291),
.A2(n_194),
.B1(n_245),
.B2(n_247),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_285),
.B(n_2),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_226),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_330),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_272),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_335),
.Y(n_355)
);

INVx13_ASAP7_75t_L g332 ( 
.A(n_269),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_266),
.B(n_235),
.C(n_249),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_295),
.Y(n_335)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_272),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_339),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_298),
.B(n_4),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_340),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_220),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_342),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_276),
.B(n_4),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_275),
.A2(n_7),
.B1(n_286),
.B2(n_299),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_343),
.A2(n_306),
.B1(n_290),
.B2(n_303),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_336),
.A2(n_280),
.B(n_279),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_346),
.A2(n_351),
.B(n_360),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_298),
.C(n_306),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_362),
.C(n_335),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_371),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_374),
.B1(n_327),
.B2(n_328),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_336),
.A2(n_264),
.B(n_301),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_287),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_354),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_333),
.A2(n_290),
.B1(n_268),
.B2(n_281),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_307),
.B(n_283),
.C(n_257),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_343),
.A2(n_287),
.B1(n_272),
.B2(n_281),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_370),
.Y(n_384)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_314),
.Y(n_369)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_337),
.A2(n_268),
.B1(n_283),
.B2(n_292),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_327),
.A2(n_287),
.B1(n_297),
.B2(n_292),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g372 ( 
.A1(n_316),
.A2(n_288),
.A3(n_267),
.B1(n_289),
.B2(n_265),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_327),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_355),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_376),
.B(n_377),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_325),
.Y(n_377)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_378),
.Y(n_420)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_344),
.Y(n_379)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_379),
.Y(n_406)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_381),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_362),
.B(n_347),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_387),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_324),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_385),
.B(n_389),
.Y(n_405)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_353),
.Y(n_386)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_318),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_273),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_365),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_390),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_391),
.B(n_394),
.Y(n_415)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_398),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_345),
.B(n_319),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_329),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_399),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_396),
.A2(n_350),
.B(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_369),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_332),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_355),
.B(n_334),
.C(n_338),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_402),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_351),
.A2(n_308),
.B(n_309),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_364),
.B(n_326),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_273),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_375),
.B(n_308),
.C(n_322),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_366),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_378),
.A2(n_371),
.B1(n_346),
.B2(n_373),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_424),
.B1(n_386),
.B2(n_381),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_359),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_409),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_374),
.B1(n_354),
.B2(n_328),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_410),
.A2(n_414),
.B1(n_419),
.B2(n_384),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_354),
.B1(n_372),
.B2(n_366),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_383),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g417 ( 
.A1(n_382),
.A2(n_367),
.B(n_359),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_417),
.Y(n_430)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_418),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_382),
.A2(n_312),
.B1(n_348),
.B2(n_361),
.Y(n_419)
);

AOI21xp33_ASAP7_75t_L g421 ( 
.A1(n_380),
.A2(n_315),
.B(n_339),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_421),
.A2(n_422),
.B(n_392),
.Y(n_442)
);

NOR3xp33_ASAP7_75t_SL g423 ( 
.A(n_401),
.B(n_340),
.C(n_364),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g443 ( 
.A(n_423),
.Y(n_443)
);

OAI22x1_ASAP7_75t_SL g424 ( 
.A1(n_384),
.A2(n_310),
.B1(n_356),
.B2(n_358),
.Y(n_424)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_412),
.B(n_394),
.C(n_387),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_435),
.C(n_438),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_425),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_434),
.A2(n_424),
.B1(n_414),
.B2(n_410),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_415),
.C(n_391),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_437),
.B(n_442),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_400),
.C(n_403),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_395),
.C(n_380),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_446),
.C(n_449),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_409),
.A2(n_398),
.B(n_379),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_441),
.B(n_358),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_407),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_445),
.B1(n_408),
.B2(n_413),
.Y(n_454)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_397),
.B1(n_390),
.B2(n_388),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_426),
.C(n_404),
.Y(n_446)
);

INVx13_ASAP7_75t_L g447 ( 
.A(n_408),
.Y(n_447)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_447),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_448),
.A2(n_427),
.B1(n_413),
.B2(n_411),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_262),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_430),
.A2(n_422),
.B(n_418),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_450),
.A2(n_442),
.B(n_429),
.Y(n_469)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_441),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_466),
.Y(n_479)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_454),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_457),
.A2(n_464),
.B1(n_448),
.B2(n_430),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_432),
.B(n_409),
.C(n_407),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_458),
.B(n_462),
.C(n_456),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_435),
.B(n_419),
.C(n_427),
.Y(n_462)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_463),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_434),
.A2(n_405),
.B1(n_411),
.B2(n_423),
.Y(n_464)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_465),
.Y(n_478)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_431),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_468),
.A2(n_457),
.B1(n_464),
.B2(n_449),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_471),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_470),
.B(n_472),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_465),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_438),
.C(n_437),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_458),
.B(n_439),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_473),
.B(n_461),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_460),
.B(n_462),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_474),
.B(n_451),
.C(n_456),
.Y(n_481)
);

BUFx12_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_475),
.Y(n_488)
);

BUFx12_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_477),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_468),
.A2(n_440),
.B1(n_446),
.B2(n_405),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_484),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_485),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_463),
.B1(n_443),
.B2(n_461),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_460),
.C(n_466),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_490),
.C(n_474),
.Y(n_496)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_487),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_455),
.C(n_453),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_483),
.A2(n_479),
.B(n_477),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_492),
.B(n_497),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_489),
.A2(n_469),
.B(n_476),
.Y(n_493)
);

OAI21x1_ASAP7_75t_L g504 ( 
.A1(n_493),
.A2(n_477),
.B(n_475),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_488),
.A2(n_478),
.B1(n_475),
.B2(n_436),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_496),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_473),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_455),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_453),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_496),
.B(n_481),
.C(n_482),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_501),
.B(n_505),
.Y(n_507)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_SL g510 ( 
.A1(n_504),
.A2(n_493),
.B(n_499),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_497),
.B(n_356),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_495),
.B(n_485),
.C(n_447),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_506),
.B(n_491),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_508),
.B(n_510),
.Y(n_512)
);

NOR3xp33_ASAP7_75t_SL g511 ( 
.A(n_509),
.B(n_500),
.C(n_502),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_262),
.Y(n_514)
);

AOI322xp5_ASAP7_75t_L g513 ( 
.A1(n_512),
.A2(n_500),
.A3(n_507),
.B1(n_495),
.B2(n_303),
.C1(n_282),
.C2(n_289),
.Y(n_513)
);

AO21x1_ASAP7_75t_L g515 ( 
.A1(n_513),
.A2(n_514),
.B(n_262),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_515),
.A2(n_295),
.B(n_257),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_516),
.B(n_7),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_267),
.B(n_7),
.Y(n_519)
);


endmodule