module real_jpeg_23754_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_88, n_11, n_14, n_90, n_7, n_3, n_5, n_4, n_1, n_89, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_88;
input n_11;
input n_14;
input n_90;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_89;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B1(n_53),
.B2(n_54),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_0),
.A2(n_53),
.B1(n_73),
.B2(n_80),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_1),
.A2(n_56),
.B1(n_58),
.B2(n_69),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_3),
.B(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_17),
.B1(n_23),
.B2(n_24),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_6),
.B(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_7),
.B(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_7),
.B(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_88),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_8),
.B(n_90),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_10),
.B(n_11),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_12),
.B(n_89),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_13),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_15),
.A2(n_17),
.B1(n_23),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_16),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_17),
.A2(n_23),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_17),
.A2(n_48),
.B(n_49),
.Y(n_47)
);

AOI221xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_55),
.B1(n_72),
.B2(n_81),
.C(n_85),
.Y(n_18)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_50),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_22),
.B(n_75),
.Y(n_74)
);

NOR3xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_32),
.C(n_40),
.Y(n_39)
);

OAI211xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_35),
.B(n_38),
.C(n_47),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_32),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_27),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_28),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_32),
.A2(n_36),
.B(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_36),
.A2(n_39),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_44),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_42),
.Y(n_40)
);

NAND3xp33_ASAP7_75t_SL g75 ( 
.A(n_47),
.B(n_76),
.C(n_79),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_60),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B(n_68),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);


endmodule