module fake_jpeg_10945_n_289 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_289);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_43),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_46),
.B(n_61),
.Y(n_104)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_47),
.Y(n_97)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_24),
.B(n_1),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_68),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g69 ( 
.A(n_40),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_26),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_77),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_74),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_41),
.B1(n_28),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_92),
.B1(n_94),
.B2(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_41),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_83),
.B(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_51),
.B1(n_67),
.B2(n_59),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_84),
.A2(n_93),
.B1(n_106),
.B2(n_2),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_25),
.B1(n_28),
.B2(n_38),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_89),
.B1(n_91),
.B2(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_36),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_47),
.A2(n_25),
.B1(n_38),
.B2(n_24),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_38),
.B1(n_35),
.B2(n_37),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_56),
.A2(n_42),
.B1(n_37),
.B2(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_30),
.B1(n_39),
.B2(n_26),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_60),
.A2(n_26),
.B1(n_21),
.B2(n_39),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_26),
.B1(n_21),
.B2(n_30),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_65),
.A2(n_42),
.B1(n_30),
.B2(n_33),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_15),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_12),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_43),
.A2(n_69),
.B1(n_4),
.B2(n_5),
.Y(n_106)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_122),
.Y(n_147)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_111),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_SL g116 ( 
.A(n_70),
.B(n_77),
.C(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_139),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_136),
.B(n_95),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_80),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_120),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_124),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_11),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_125),
.Y(n_148)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_128),
.B(n_130),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_2),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_131),
.A2(n_94),
.B1(n_90),
.B2(n_108),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_85),
.B(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_132),
.B(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_79),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_84),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_137),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_78),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_8),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_96),
.Y(n_164)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_80),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_97),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_142),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_162),
.B1(n_100),
.B2(n_96),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_108),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_134),
.C(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_135),
.C(n_9),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_160),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g160 ( 
.A(n_110),
.B(n_112),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_131),
.A2(n_107),
.B1(n_95),
.B2(n_100),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_107),
.B1(n_81),
.B2(n_85),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_163),
.A2(n_126),
.B1(n_142),
.B2(n_111),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_120),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_81),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_168),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_172),
.B(n_186),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_152),
.B(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_119),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_126),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_192),
.C(n_166),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_197),
.B1(n_166),
.B2(n_143),
.Y(n_211)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_181),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_109),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_183),
.B(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_117),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_141),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_161),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_188),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_113),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_189),
.B(n_143),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_193),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_123),
.B(n_118),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_191),
.A2(n_171),
.B(n_165),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_194),
.A2(n_196),
.B(n_169),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_144),
.A2(n_125),
.B1(n_10),
.B2(n_11),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_148),
.B1(n_169),
.B2(n_159),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_161),
.A2(n_164),
.B(n_154),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_163),
.B1(n_162),
.B2(n_158),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_165),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_177),
.A2(n_158),
.B1(n_146),
.B2(n_171),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_216),
.B1(n_217),
.B2(n_178),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_179),
.B(n_153),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_210),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_205),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_218),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_211),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_203),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_174),
.A2(n_173),
.B1(n_172),
.B2(n_176),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_185),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_220),
.Y(n_235)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_200),
.A2(n_180),
.B(n_197),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_232),
.B(n_211),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_237),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_182),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_238),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_209),
.B1(n_217),
.B2(n_218),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_226),
.A2(n_233),
.B1(n_228),
.B2(n_221),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_214),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_230),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_173),
.B(n_191),
.C(n_196),
.D(n_194),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_206),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_192),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_244),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_190),
.B(n_195),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_228),
.A2(n_219),
.B1(n_205),
.B2(n_188),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_242),
.A2(n_222),
.B1(n_216),
.B2(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_229),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_231),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_225),
.C(n_233),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_235),
.A2(n_220),
.B(n_204),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_249),
.A2(n_232),
.B(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_181),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_251),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_255),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_241),
.B1(n_242),
.B2(n_247),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_222),
.C(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.C(n_255),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_215),
.C(n_208),
.Y(n_259)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_243),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_184),
.Y(n_267)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_261),
.A2(n_249),
.B(n_245),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_268),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_240),
.B1(n_208),
.B2(n_237),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_269),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_239),
.C(n_193),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_259),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_269),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_263),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_274),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_268),
.B(n_257),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_253),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_279),
.B(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_254),
.C(n_252),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_280),
.B(n_254),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_281),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_278),
.A2(n_275),
.B(n_276),
.Y(n_282)
);

AOI322xp5_ASAP7_75t_L g285 ( 
.A1(n_282),
.A2(n_283),
.A3(n_237),
.B1(n_260),
.B2(n_253),
.C1(n_256),
.C2(n_267),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_261),
.B(n_260),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_284),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_198),
.C(n_159),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_288),
.Y(n_289)
);


endmodule