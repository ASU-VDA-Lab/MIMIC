module fake_jpeg_18048_n_257 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_257);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_53),
.A2(n_55),
.B1(n_46),
.B2(n_42),
.Y(n_79)
);

O2A1O1Ixp33_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_14),
.B(n_13),
.C(n_24),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_54),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_51),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_63),
.B(n_13),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_70),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g61 ( 
.A(n_47),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_70),
.B1(n_71),
.B2(n_50),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_49),
.A2(n_35),
.B1(n_34),
.B2(n_28),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_48),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_20),
.B(n_21),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_68),
.Y(n_72)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_38),
.A2(n_18),
.B1(n_22),
.B2(n_20),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_18),
.B1(n_13),
.B2(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_22),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_24),
.B1(n_14),
.B2(n_23),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_84),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_80),
.B1(n_55),
.B2(n_69),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_15),
.B1(n_21),
.B2(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_50),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_44),
.Y(n_111)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_64),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_48),
.Y(n_106)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_99),
.B(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_72),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_101),
.Y(n_119)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_72),
.B(n_54),
.CI(n_55),
.CON(n_100),
.SN(n_100)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_100),
.B(n_15),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_62),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_86),
.A2(n_62),
.B1(n_71),
.B2(n_29),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_104),
.A2(n_92),
.B1(n_91),
.B2(n_73),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_91),
.B1(n_92),
.B2(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_82),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_110),
.B(n_77),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_64),
.B(n_85),
.Y(n_129)
);

CKINVDCx6p67_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_114),
.A2(n_94),
.B1(n_108),
.B2(n_107),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_131),
.B(n_134),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_127),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_91),
.B1(n_75),
.B2(n_78),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_122),
.B1(n_130),
.B2(n_132),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_76),
.C(n_82),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_124),
.C(n_45),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_76),
.B1(n_89),
.B2(n_85),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_33),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_96),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_133),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_106),
.A2(n_85),
.B1(n_60),
.B2(n_40),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_14),
.B(n_25),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_95),
.A2(n_60),
.B1(n_15),
.B2(n_25),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_0),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_105),
.B1(n_104),
.B2(n_100),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_103),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_141),
.B(n_142),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_110),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_147),
.B(n_157),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_131),
.B1(n_112),
.B2(n_31),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_133),
.A2(n_98),
.B(n_102),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_93),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_142),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_98),
.Y(n_150)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_0),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_21),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_126),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_117),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_114),
.A2(n_23),
.B1(n_112),
.B2(n_17),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_155),
.A2(n_17),
.B1(n_26),
.B2(n_33),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_132),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_115),
.A2(n_43),
.B(n_112),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_144),
.A2(n_123),
.B1(n_117),
.B2(n_126),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_158),
.A2(n_178),
.B1(n_159),
.B2(n_170),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_120),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_161),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_152),
.Y(n_162)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_156),
.C(n_143),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_175),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_145),
.B1(n_139),
.B2(n_149),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_138),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_7),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_137),
.B(n_90),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_90),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_177),
.Y(n_188)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_182),
.C(n_185),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_166),
.B(n_140),
.C(n_136),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_174),
.A2(n_145),
.B1(n_157),
.B2(n_155),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_161),
.A2(n_140),
.B1(n_146),
.B2(n_135),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_177),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_173),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_191),
.B(n_185),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_176),
.B1(n_165),
.B2(n_173),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_143),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_193),
.B(n_160),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_160),
.A2(n_135),
.B1(n_2),
.B2(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_195),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_172),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_203),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_162),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.C(n_184),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_191),
.B(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_178),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_202),
.B(n_209),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_208),
.A2(n_187),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_159),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_199),
.A2(n_188),
.B1(n_180),
.B2(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_213),
.Y(n_224)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_186),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_198),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_207),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_17),
.C(n_26),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_203),
.C(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_208),
.Y(n_220)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_222),
.B(n_228),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_26),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_10),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_8),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_217),
.A2(n_10),
.B1(n_12),
.B2(n_6),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_231),
.B(n_220),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_215),
.C(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_234),
.C(n_6),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_235),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_218),
.C(n_219),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_225),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_237),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_238),
.B(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_230),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_240),
.B(n_241),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_10),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_245),
.B(n_7),
.Y(n_247)
);

XNOR2x2_ASAP7_75t_SL g246 ( 
.A(n_243),
.B(n_7),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_249),
.B(n_4),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_11),
.B(n_12),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_248),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_251),
.B(n_5),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_4),
.C(n_5),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_4),
.C(n_26),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_255),
.B(n_26),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_256),
.A2(n_26),
.B(n_243),
.Y(n_257)
);


endmodule