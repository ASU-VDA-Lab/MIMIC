module real_jpeg_7319_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_1),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_1),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_70),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_1),
.B(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_1),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_1),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_1),
.B(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_2),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_2),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_2),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_2),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_3),
.B(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_3),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_79),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_3),
.B(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_3),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_4),
.Y(n_200)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_4),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_5),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_5),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_5),
.B(n_364),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_5),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_5),
.B(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_5),
.B(n_397),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_5),
.B(n_438),
.Y(n_437)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_7),
.B(n_14),
.Y(n_344)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_8),
.Y(n_280)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_10),
.B(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_10),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_10),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_10),
.B(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_10),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_10),
.B(n_390),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_10),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_10),
.B(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_11),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_11),
.Y(n_156)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_11),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_12),
.B(n_22),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_12),
.B(n_26),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_12),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_12),
.B(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_12),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_12),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_12),
.B(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_13),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_13),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_14),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_14),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_14),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_14),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_14),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_15),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_15),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_15),
.B(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_15),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_110),
.B(n_125),
.C(n_497),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_19),
.B(n_101),
.CI(n_102),
.CON(n_100),
.SN(n_100)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.C(n_29),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_20),
.A2(n_21),
.B1(n_29),
.B2(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_20),
.A2(n_21),
.B1(n_105),
.B2(n_108),
.Y(n_104)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_20),
.B(n_46),
.C(n_105),
.Y(n_497)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_21),
.B(n_183),
.C(n_186),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_21),
.B(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_24),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_25),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_25),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_25),
.A2(n_88),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_137),
.C(n_141),
.Y(n_166)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_29),
.A2(n_41),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_29),
.B(n_233),
.C(n_237),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_29),
.A2(n_76),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_34),
.Y(n_374)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_35),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_100),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_83),
.C(n_84),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_38),
.B(n_495),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_62),
.C(n_73),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_39),
.B(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_54),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_40),
.B(n_58),
.C(n_60),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.C(n_49),
.Y(n_40)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_41),
.B(n_76),
.C(n_82),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_41),
.A2(n_77),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_41),
.A2(n_77),
.B1(n_257),
.B2(n_258),
.Y(n_297)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_44),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_44),
.Y(n_300)
);

INVx6_ASAP7_75t_L g371 ( 
.A(n_44),
.Y(n_371)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_45),
.Y(n_130)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_45),
.Y(n_240)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_45),
.Y(n_394)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_45),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_46),
.A2(n_103),
.B1(n_104),
.B2(n_109),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_46),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_46),
.A2(n_49),
.B1(n_50),
.B2(n_109),
.Y(n_165)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_49),
.A2(n_50),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_120),
.C(n_126),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_49),
.A2(n_50),
.B1(n_301),
.B2(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_50),
.B(n_299),
.C(n_301),
.Y(n_298)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_52),
.Y(n_420)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_52),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_58),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_62),
.B(n_73),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.C(n_69),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_66),
.B1(n_67),
.B2(n_145),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_63),
.Y(n_145)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_66),
.A2(n_67),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_67),
.B(n_150),
.C(n_197),
.Y(n_196)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_69),
.B(n_144),
.Y(n_143)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_72),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_72),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_82),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_77),
.B(n_257),
.C(n_262),
.Y(n_256)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_126),
.C(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_78),
.A2(n_82),
.B1(n_128),
.B2(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_83),
.B(n_84),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_99),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_93),
.C(n_99),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g499 ( 
.A(n_100),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_105),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_105),
.B(n_196),
.C(n_201),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_105),
.A2(n_108),
.B1(n_157),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_105),
.A2(n_108),
.B1(n_201),
.B2(n_245),
.Y(n_244)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_148),
.C(n_157),
.Y(n_147)
);

AO21x1_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_492),
.B(n_496),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_247),
.B(n_489),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_211),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_SL g489 ( 
.A1(n_113),
.A2(n_490),
.B(n_491),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_170),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_114),
.B(n_170),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_161),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_115),
.B(n_162),
.C(n_168),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_143),
.C(n_146),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_116),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_127),
.C(n_131),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_117),
.B(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_122),
.B1(n_125),
.B2(n_126),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_122),
.A2(n_126),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_122),
.B(n_234),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_122),
.A2(n_126),
.B1(n_233),
.B2(n_234),
.Y(n_456)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_123),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_124),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_127),
.B(n_131),
.Y(n_216)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_137),
.B1(n_141),
.B2(n_142),
.Y(n_133)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_137),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_137),
.B(n_225),
.Y(n_255)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_142),
.B(n_224),
.C(n_226),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_143),
.A2(n_146),
.B1(n_147),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g207 ( 
.A1(n_148),
.A2(n_149),
.B1(n_208),
.B2(n_210),
.Y(n_207)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_150),
.A2(n_155),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_150),
.A2(n_191),
.B1(n_197),
.B2(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_150),
.A2(n_191),
.B1(n_410),
.B2(n_415),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_150),
.B(n_415),
.Y(n_457)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_152),
.Y(n_408)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_152),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_153),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_153),
.B(n_271),
.C(n_274),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_153),
.A2(n_193),
.B1(n_271),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_157),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_160),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_160),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_167),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_176),
.Y(n_170)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_171),
.B(n_174),
.CI(n_176),
.CON(n_246),
.SN(n_246)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_195),
.C(n_207),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_189),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_178),
.B(n_182),
.Y(n_318)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_186),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_185),
.Y(n_287)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_189),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_207),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_196),
.B(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_197),
.B(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_197),
.A2(n_222),
.B1(n_305),
.B2(n_306),
.Y(n_376)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_199),
.Y(n_414)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_205),
.Y(n_302)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_206),
.Y(n_400)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_246),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_212),
.B(n_246),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_217),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_213),
.B(n_215),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_217),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_231),
.C(n_243),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_218),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_223),
.C(n_229),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_219),
.B(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_223),
.B(n_229),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_243),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_239),
.C(n_241),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_232),
.B(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_233),
.A2(n_234),
.B1(n_237),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_237),
.Y(n_312)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_238),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_239),
.A2(n_241),
.B1(n_242),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_239),
.Y(n_291)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g500 ( 
.A(n_246),
.Y(n_500)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_382),
.B1(n_482),
.B2(n_487),
.C(n_488),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_322),
.C(n_326),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_249),
.A2(n_483),
.B(n_486),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_315),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_250),
.B(n_315),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_292),
.C(n_294),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_251),
.B(n_292),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_277),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_252),
.B(n_278),
.C(n_289),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_269),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_254),
.B(n_270),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_256),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_262),
.B(n_297),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_333),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_289),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_285),
.C(n_288),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_279),
.A2(n_281),
.B(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_288),
.Y(n_314)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_352),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_309),
.C(n_313),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_298),
.C(n_303),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_378),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_298),
.A2(n_303),
.B1(n_304),
.B2(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_298),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_299),
.B(n_359),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_301),
.Y(n_360)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_313),
.Y(n_330)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_321),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_319),
.C(n_321),
.Y(n_323)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_322),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_323),
.B(n_324),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_353),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_327),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_351),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_328),
.B(n_351),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_331),
.C(n_349),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_329),
.B(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_331),
.B(n_349),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.C(n_340),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_335),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_337),
.B(n_419),
.Y(n_418)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_340),
.B(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.C(n_345),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_341),
.A2(n_342),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_343),
.A2(n_344),
.B1(n_345),
.B2(n_346),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_380),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_354),
.B(n_380),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_357),
.C(n_377),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_355),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_357),
.B(n_377),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.C(n_375),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_358),
.B(n_473),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_361),
.A2(n_375),
.B1(n_376),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_361),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_367),
.C(n_372),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_362),
.A2(n_363),
.B1(n_372),
.B2(n_373),
.Y(n_461)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_367),
.B(n_461),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_404),
.Y(n_403)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_383),
.A2(n_477),
.B(n_481),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_463),
.B(n_476),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_450),
.B(n_462),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_426),
.B(n_449),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_416),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_387),
.B(n_416),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_401),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_402),
.C(n_409),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_395),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_389),
.B(n_396),
.C(n_398),
.Y(n_459)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_409),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_406),
.Y(n_417)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_404),
.Y(n_438)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_410),
.Y(n_415)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_418),
.C(n_421),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_417),
.B(n_446),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_418),
.A2(n_421),
.B1(n_422),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_418),
.Y(n_447)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_443),
.B(n_448),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_436),
.B(n_442),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_435),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_435),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_433),
.Y(n_444)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_434),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_445),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_451),
.B(n_452),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_459),
.C(n_460),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g498 ( 
.A(n_453),
.Y(n_498)
);

FAx1_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_456),
.CI(n_457),
.CON(n_453),
.SN(n_453)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_454),
.B(n_456),
.C(n_457),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_475),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_475),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_472),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_466),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_466),
.B(n_469),
.C(n_472),
.Y(n_478)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_470),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_479),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_493),
.B(n_494),
.Y(n_496)
);


endmodule