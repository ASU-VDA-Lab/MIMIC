module real_aes_7682_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_725;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g272 ( .A1(n_0), .A2(n_273), .B(n_274), .C(n_277), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_1), .B(n_261), .Y(n_278) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_3), .B(n_189), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_4), .A2(n_150), .B(n_153), .C(n_533), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_5), .A2(n_145), .B(n_557), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_6), .A2(n_104), .B1(n_115), .B2(n_759), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_7), .A2(n_145), .B(n_255), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_8), .B(n_261), .Y(n_563) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_9), .A2(n_180), .B(n_217), .Y(n_216) );
AND2x6_ASAP7_75t_L g150 ( .A(n_10), .B(n_151), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g233 ( .A1(n_11), .A2(n_150), .B(n_153), .C(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g501 ( .A(n_12), .Y(n_501) );
INVx1_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_13), .B(n_41), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_14), .B(n_237), .Y(n_535) );
INVx1_ASAP7_75t_L g171 ( .A(n_15), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_16), .B(n_189), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_17), .A2(n_190), .B(n_519), .C(n_521), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_18), .B(n_261), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_19), .B(n_165), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g152 ( .A1(n_20), .A2(n_153), .B(n_156), .C(n_164), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_21), .A2(n_225), .B(n_276), .C(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_22), .B(n_237), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_23), .A2(n_55), .B1(n_755), .B2(n_756), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_23), .Y(n_755) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_24), .B(n_237), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g548 ( .A(n_25), .Y(n_548) );
INVx1_ASAP7_75t_L g473 ( .A(n_26), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_27), .A2(n_153), .B(n_164), .C(n_220), .Y(n_219) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_28), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_29), .Y(n_531) );
INVx1_ASAP7_75t_L g489 ( .A(n_30), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_31), .A2(n_145), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g148 ( .A(n_32), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_33), .A2(n_193), .B(n_202), .C(n_204), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_34), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_35), .A2(n_276), .B(n_560), .C(n_562), .Y(n_559) );
INVxp67_ASAP7_75t_L g490 ( .A(n_36), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_37), .B(n_222), .Y(n_221) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_38), .A2(n_153), .B(n_164), .C(n_472), .Y(n_471) );
CKINVDCx14_ASAP7_75t_R g558 ( .A(n_39), .Y(n_558) );
AOI222xp33_ASAP7_75t_SL g127 ( .A1(n_40), .A2(n_128), .B1(n_134), .B2(n_739), .C1(n_740), .C2(n_744), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_42), .A2(n_277), .B(n_499), .C(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_43), .B(n_144), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g239 ( .A(n_44), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_45), .B(n_189), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_46), .B(n_145), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_47), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_48), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_49), .A2(n_193), .B(n_202), .C(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g275 ( .A(n_50), .Y(n_275) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_51), .A2(n_753), .B1(n_754), .B2(n_757), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g757 ( .A(n_51), .Y(n_757) );
INVx1_ASAP7_75t_L g247 ( .A(n_52), .Y(n_247) );
INVx1_ASAP7_75t_L g507 ( .A(n_53), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_54), .B(n_145), .Y(n_244) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_55), .Y(n_756) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_56), .Y(n_173) );
CKINVDCx14_ASAP7_75t_R g497 ( .A(n_57), .Y(n_497) );
INVx1_ASAP7_75t_L g151 ( .A(n_58), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_59), .B(n_145), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_60), .B(n_261), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_61), .A2(n_163), .B(n_186), .C(n_258), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_62), .Y(n_126) );
INVx1_ASAP7_75t_L g170 ( .A(n_63), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_64), .A2(n_102), .B1(n_130), .B2(n_131), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_64), .Y(n_131) );
INVx1_ASAP7_75t_SL g561 ( .A(n_65), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_66), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_67), .B(n_189), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_68), .B(n_261), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_69), .B(n_190), .Y(n_235) );
INVx1_ASAP7_75t_L g551 ( .A(n_70), .Y(n_551) );
CKINVDCx16_ASAP7_75t_R g271 ( .A(n_71), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_72), .B(n_158), .Y(n_157) );
A2O1A1Ixp33_ASAP7_75t_L g183 ( .A1(n_73), .A2(n_153), .B(n_184), .C(n_193), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_74), .Y(n_256) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_76), .A2(n_145), .B(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g554 ( .A(n_77), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_78), .A2(n_145), .B(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_79), .A2(n_144), .B(n_485), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_80), .Y(n_470) );
INVx1_ASAP7_75t_L g517 ( .A(n_81), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_82), .B(n_161), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_83), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_84), .A2(n_145), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g520 ( .A(n_85), .Y(n_520) );
INVx2_ASAP7_75t_L g168 ( .A(n_86), .Y(n_168) );
INVx1_ASAP7_75t_L g534 ( .A(n_87), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_88), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_89), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g122 ( .A(n_90), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g462 ( .A(n_90), .B(n_124), .Y(n_462) );
OAI22xp5_ASAP7_75t_SL g128 ( .A1(n_91), .A2(n_129), .B1(n_132), .B2(n_133), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_91), .Y(n_133) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_92), .A2(n_153), .B(n_193), .C(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_93), .B(n_145), .Y(n_200) );
INVx1_ASAP7_75t_L g205 ( .A(n_94), .Y(n_205) );
INVxp67_ASAP7_75t_L g259 ( .A(n_95), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_96), .B(n_180), .Y(n_502) );
INVx2_ASAP7_75t_L g510 ( .A(n_97), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g185 ( .A(n_99), .Y(n_185) );
INVx1_ASAP7_75t_L g231 ( .A(n_100), .Y(n_231) );
AND2x2_ASAP7_75t_L g249 ( .A(n_101), .B(n_167), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_102), .Y(n_130) );
INVx1_ASAP7_75t_SL g759 ( .A(n_104), .Y(n_759) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g124 ( .A(n_110), .B(n_125), .Y(n_124) );
OR2x2_ASAP7_75t_L g738 ( .A(n_111), .B(n_124), .Y(n_738) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_111), .B(n_123), .Y(n_746) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_127), .B1(n_747), .B2(n_749), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g748 ( .A(n_119), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_120), .A2(n_750), .B(n_758), .Y(n_749) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_126), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g758 ( .A(n_122), .Y(n_758) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx1_ASAP7_75t_L g739 ( .A(n_128), .Y(n_739) );
INVx1_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
OAI22xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_460), .B1(n_463), .B2(n_736), .Y(n_134) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_135), .A2(n_742), .B1(n_751), .B2(n_752), .Y(n_750) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx2_ASAP7_75t_L g742 ( .A(n_136), .Y(n_742) );
AND3x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_364), .C(n_421), .Y(n_136) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_309), .C(n_345), .Y(n_137) );
OAI211xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_211), .B(n_263), .C(n_296), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_175), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x4_ASAP7_75t_L g266 ( .A(n_141), .B(n_267), .Y(n_266) );
INVx5_ASAP7_75t_L g295 ( .A(n_141), .Y(n_295) );
AND2x2_ASAP7_75t_L g368 ( .A(n_141), .B(n_284), .Y(n_368) );
AND2x2_ASAP7_75t_L g406 ( .A(n_141), .B(n_312), .Y(n_406) );
AND2x2_ASAP7_75t_L g426 ( .A(n_141), .B(n_268), .Y(n_426) );
OR2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_172), .Y(n_141) );
AOI21xp5_ASAP7_75t_SL g142 ( .A1(n_143), .A2(n_152), .B(n_165), .Y(n_142) );
BUFx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g232 ( .A(n_146), .B(n_150), .Y(n_232) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g163 ( .A(n_147), .Y(n_163) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g154 ( .A(n_148), .Y(n_154) );
INVx1_ASAP7_75t_L g226 ( .A(n_148), .Y(n_226) );
INVx1_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g190 ( .A(n_149), .Y(n_190) );
INVx1_ASAP7_75t_L g222 ( .A(n_149), .Y(n_222) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_149), .Y(n_237) );
BUFx3_ASAP7_75t_L g164 ( .A(n_150), .Y(n_164) );
INVx4_ASAP7_75t_SL g194 ( .A(n_150), .Y(n_194) );
INVx5_ASAP7_75t_L g203 ( .A(n_153), .Y(n_203) );
AND2x6_ASAP7_75t_L g153 ( .A(n_154), .B(n_155), .Y(n_153) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
BUFx3_ASAP7_75t_L g208 ( .A(n_154), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_160), .B(n_162), .Y(n_156) );
INVx2_ASAP7_75t_L g161 ( .A(n_158), .Y(n_161) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_161), .A2(n_205), .B(n_206), .C(n_207), .Y(n_204) );
O2A1O1Ixp33_ASAP7_75t_L g246 ( .A1(n_161), .A2(n_207), .B(n_247), .C(n_248), .Y(n_246) );
O2A1O1Ixp5_ASAP7_75t_L g533 ( .A1(n_161), .A2(n_534), .B(n_535), .C(n_536), .Y(n_533) );
O2A1O1Ixp33_ASAP7_75t_L g550 ( .A1(n_161), .A2(n_536), .B(n_551), .C(n_552), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_162), .A2(n_189), .B(n_473), .C(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_163), .B(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_166), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g174 ( .A(n_167), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_167), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_167), .A2(n_244), .B(n_245), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_167), .A2(n_232), .B(n_470), .C(n_471), .Y(n_469) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_167), .A2(n_495), .B(n_502), .Y(n_494) );
AND2x2_ASAP7_75t_SL g167 ( .A(n_168), .B(n_169), .Y(n_167) );
AND2x2_ASAP7_75t_L g181 ( .A(n_168), .B(n_169), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_170), .B(n_171), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_173), .B(n_174), .Y(n_172) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_174), .A2(n_530), .B(n_537), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_175), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_198), .Y(n_175) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_176), .Y(n_307) );
AND2x2_ASAP7_75t_L g321 ( .A(n_176), .B(n_267), .Y(n_321) );
INVx1_ASAP7_75t_L g344 ( .A(n_176), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_176), .B(n_295), .Y(n_383) );
OR2x2_ASAP7_75t_L g420 ( .A(n_176), .B(n_265), .Y(n_420) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_177), .Y(n_356) );
AND2x2_ASAP7_75t_L g363 ( .A(n_177), .B(n_268), .Y(n_363) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g284 ( .A(n_178), .B(n_268), .Y(n_284) );
BUFx2_ASAP7_75t_L g312 ( .A(n_178), .Y(n_312) );
AO21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_182), .B(n_196), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_179), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_179), .B(n_210), .Y(n_209) );
AO21x2_ASAP7_75t_L g229 ( .A1(n_179), .A2(n_230), .B(n_238), .Y(n_229) );
INVx3_ASAP7_75t_L g261 ( .A(n_179), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_179), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_179), .B(n_538), .Y(n_537) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_179), .A2(n_547), .B(n_553), .Y(n_546) );
INVx4_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_180), .A2(n_218), .B(n_219), .Y(n_217) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_180), .Y(n_253) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g240 ( .A(n_181), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_195), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_188), .C(n_191), .Y(n_184) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_187), .A2(n_189), .B1(n_489), .B2(n_490), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_187), .B(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_187), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_189), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g273 ( .A(n_189), .Y(n_273) );
INVx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_190), .B(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g562 ( .A(n_192), .Y(n_562) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g255 ( .A1(n_194), .A2(n_203), .B(n_256), .C(n_257), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_194), .A2(n_203), .B(n_271), .C(n_272), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_194), .A2(n_203), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_194), .A2(n_203), .B(n_497), .C(n_498), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_SL g506 ( .A1(n_194), .A2(n_203), .B(n_507), .C(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_194), .A2(n_203), .B(n_517), .C(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g557 ( .A1(n_194), .A2(n_203), .B(n_558), .C(n_559), .Y(n_557) );
INVx5_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
BUFx2_ASAP7_75t_L g288 ( .A(n_198), .Y(n_288) );
AND2x2_ASAP7_75t_L g445 ( .A(n_198), .B(n_299), .Y(n_445) );
OR2x6_ASAP7_75t_L g198 ( .A(n_199), .B(n_209), .Y(n_198) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
INVx1_ASAP7_75t_L g521 ( .A(n_208), .Y(n_521) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
NAND2xp33_ASAP7_75t_L g212 ( .A(n_213), .B(n_250), .Y(n_212) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_213), .A2(n_346), .B1(n_353), .B2(n_354), .C(n_357), .Y(n_345) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_227), .Y(n_213) );
AND2x2_ASAP7_75t_L g251 ( .A(n_214), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_214), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g280 ( .A(n_215), .B(n_228), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g290 ( .A(n_215), .B(n_229), .Y(n_290) );
OR2x2_ASAP7_75t_L g301 ( .A(n_215), .B(n_252), .Y(n_301) );
AND2x2_ASAP7_75t_L g304 ( .A(n_215), .B(n_292), .Y(n_304) );
AND2x2_ASAP7_75t_L g320 ( .A(n_215), .B(n_241), .Y(n_320) );
OR2x2_ASAP7_75t_L g336 ( .A(n_215), .B(n_229), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_215), .B(n_252), .Y(n_398) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_216), .B(n_241), .Y(n_390) );
AND2x2_ASAP7_75t_L g393 ( .A(n_216), .B(n_229), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_223), .B(n_224), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_224), .A2(n_235), .B(n_236), .Y(n_234) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g314 ( .A(n_227), .B(n_301), .Y(n_314) );
INVx2_ASAP7_75t_L g340 ( .A(n_227), .Y(n_340) );
OR2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_241), .Y(n_227) );
AND2x2_ASAP7_75t_L g262 ( .A(n_228), .B(n_242), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_228), .B(n_252), .Y(n_319) );
OR2x2_ASAP7_75t_L g330 ( .A(n_228), .B(n_242), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_228), .B(n_292), .Y(n_389) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_228), .A2(n_423), .B1(n_425), .B2(n_427), .C(n_430), .Y(n_422) );
INVx5_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_229), .B(n_252), .Y(n_361) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_232), .B(n_233), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_232), .A2(n_531), .B(n_532), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g547 ( .A1(n_232), .A2(n_548), .B(n_549), .Y(n_547) );
INVx4_ASAP7_75t_L g276 ( .A(n_237), .Y(n_276) );
INVx2_ASAP7_75t_L g499 ( .A(n_237), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx2_ASAP7_75t_L g482 ( .A(n_240), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_241), .B(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_241), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g308 ( .A(n_241), .B(n_280), .Y(n_308) );
OR2x2_ASAP7_75t_L g352 ( .A(n_241), .B(n_252), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_241), .B(n_304), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_241), .B(n_397), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_241), .B(n_418), .Y(n_417) );
INVx5_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_SL g281 ( .A(n_242), .B(n_251), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_SL g285 ( .A1(n_242), .A2(n_286), .B(n_289), .C(n_293), .Y(n_285) );
OR2x2_ASAP7_75t_L g323 ( .A(n_242), .B(n_319), .Y(n_323) );
OR2x2_ASAP7_75t_L g359 ( .A(n_242), .B(n_301), .Y(n_359) );
OAI311xp33_ASAP7_75t_L g365 ( .A1(n_242), .A2(n_304), .A3(n_366), .B1(n_369), .C1(n_376), .Y(n_365) );
AND2x2_ASAP7_75t_L g416 ( .A(n_242), .B(n_252), .Y(n_416) );
AND2x2_ASAP7_75t_L g424 ( .A(n_242), .B(n_279), .Y(n_424) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_242), .Y(n_442) );
AND2x2_ASAP7_75t_L g459 ( .A(n_242), .B(n_280), .Y(n_459) );
OR2x6_ASAP7_75t_L g242 ( .A(n_243), .B(n_249), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_262), .Y(n_250) );
AND2x2_ASAP7_75t_L g287 ( .A(n_251), .B(n_288), .Y(n_287) );
INVx2_ASAP7_75t_L g443 ( .A(n_251), .Y(n_443) );
AND2x2_ASAP7_75t_L g279 ( .A(n_252), .B(n_280), .Y(n_279) );
INVx3_ASAP7_75t_L g292 ( .A(n_252), .Y(n_292) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_252), .Y(n_335) );
INVxp67_ASAP7_75t_L g374 ( .A(n_252), .Y(n_374) );
OA21x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_260), .Y(n_252) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_253), .A2(n_505), .B(n_511), .Y(n_504) );
OA21x2_ASAP7_75t_L g514 ( .A1(n_253), .A2(n_515), .B(n_522), .Y(n_514) );
OA21x2_ASAP7_75t_L g555 ( .A1(n_253), .A2(n_556), .B(n_563), .Y(n_555) );
OA21x2_ASAP7_75t_L g268 ( .A1(n_261), .A2(n_269), .B(n_278), .Y(n_268) );
AND2x2_ASAP7_75t_L g452 ( .A(n_262), .B(n_300), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_279), .B1(n_281), .B2(n_282), .C(n_285), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_265), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g305 ( .A(n_265), .B(n_295), .Y(n_305) );
AND2x2_ASAP7_75t_L g313 ( .A(n_265), .B(n_267), .Y(n_313) );
OR2x2_ASAP7_75t_L g325 ( .A(n_265), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g343 ( .A(n_265), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g367 ( .A(n_265), .B(n_368), .Y(n_367) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_265), .Y(n_387) );
AND2x2_ASAP7_75t_L g439 ( .A(n_265), .B(n_363), .Y(n_439) );
OAI31xp33_ASAP7_75t_L g447 ( .A1(n_265), .A2(n_316), .A3(n_415), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_266), .B(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g411 ( .A(n_266), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_266), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g299 ( .A(n_267), .B(n_295), .Y(n_299) );
INVx1_ASAP7_75t_L g386 ( .A(n_267), .Y(n_386) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g436 ( .A(n_268), .B(n_295), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_276), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g536 ( .A(n_277), .Y(n_536) );
INVx1_ASAP7_75t_SL g446 ( .A(n_279), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_280), .B(n_351), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g430 ( .A1(n_281), .A2(n_393), .B1(n_431), .B2(n_434), .Y(n_430) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g294 ( .A(n_284), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_284), .B(n_305), .Y(n_458) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g428 ( .A(n_287), .B(n_429), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_288), .A2(n_347), .B(n_349), .Y(n_346) );
OR2x2_ASAP7_75t_L g354 ( .A(n_288), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g375 ( .A(n_288), .B(n_363), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_288), .B(n_386), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_288), .B(n_426), .Y(n_425) );
OAI221xp5_ASAP7_75t_SL g402 ( .A1(n_289), .A2(n_403), .B1(n_408), .B2(n_411), .C(n_412), .Y(n_402) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
OR2x2_ASAP7_75t_L g379 ( .A(n_290), .B(n_352), .Y(n_379) );
INVx1_ASAP7_75t_L g418 ( .A(n_290), .Y(n_418) );
INVx2_ASAP7_75t_L g394 ( .A(n_291), .Y(n_394) );
INVx1_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
INVx1_ASAP7_75t_SL g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_295), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g362 ( .A(n_295), .B(n_363), .Y(n_362) );
OR2x2_ASAP7_75t_L g450 ( .A(n_295), .B(n_420), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_302), .B2(n_305), .C1(n_306), .C2(n_308), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g306 ( .A(n_299), .B(n_307), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_299), .A2(n_349), .B1(n_377), .B2(n_378), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_299), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OAI21xp33_ASAP7_75t_SL g337 ( .A1(n_308), .A2(n_338), .B(n_341), .Y(n_337) );
OAI211xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_314), .B(n_315), .C(n_337), .Y(n_309) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g315 ( .A1(n_313), .A2(n_316), .B1(n_321), .B2(n_322), .C(n_324), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_313), .B(n_401), .Y(n_400) );
INVxp67_ASAP7_75t_L g407 ( .A(n_313), .Y(n_407) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g409 ( .A(n_318), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g326 ( .A(n_321), .Y(n_326) );
AND2x2_ASAP7_75t_L g332 ( .A(n_321), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_331), .B2(n_334), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_328), .B(n_340), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_329), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g429 ( .A(n_333), .Y(n_429) );
AND2x2_ASAP7_75t_L g448 ( .A(n_333), .B(n_363), .Y(n_448) );
OR2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_340), .B(n_397), .Y(n_456) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_343), .B(n_411), .Y(n_454) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g377 ( .A(n_355), .Y(n_377) );
BUFx2_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
OAI21xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_360), .B(n_362), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_380), .C(n_402), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_372), .B(n_375), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
A2O1A1Ixp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_384), .B(n_388), .C(n_391), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_381), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp67_ASAP7_75t_SL g385 ( .A(n_386), .B(n_387), .Y(n_385) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_SL g410 ( .A(n_390), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B(n_399), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x2_ASAP7_75t_L g415 ( .A(n_393), .B(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_415), .B1(n_417), .B2(n_419), .Y(n_412) );
INVx2_ASAP7_75t_SL g433 ( .A(n_420), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_437), .C(n_449), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_433), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B1(n_444), .B2(n_446), .C(n_447), .Y(n_437) );
A2O1A1Ixp33_ASAP7_75t_L g449 ( .A1(n_438), .A2(n_450), .B(n_451), .C(n_453), .Y(n_449) );
INVx1_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B1(n_457), .B2(n_459), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g741 ( .A(n_461), .Y(n_741) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g743 ( .A(n_463), .Y(n_743) );
OR5x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_630), .C(n_694), .D(n_710), .E(n_725), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_465), .B(n_564), .C(n_591), .D(n_614), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_512), .B(n_523), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_477), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_SL g543 ( .A(n_468), .Y(n_543) );
AND2x4_ASAP7_75t_L g577 ( .A(n_468), .B(n_566), .Y(n_577) );
OR2x2_ASAP7_75t_L g587 ( .A(n_468), .B(n_545), .Y(n_587) );
OR2x2_ASAP7_75t_L g633 ( .A(n_468), .B(n_480), .Y(n_633) );
AND2x2_ASAP7_75t_L g647 ( .A(n_468), .B(n_544), .Y(n_647) );
AND2x2_ASAP7_75t_L g690 ( .A(n_468), .B(n_580), .Y(n_690) );
AND2x2_ASAP7_75t_L g697 ( .A(n_468), .B(n_555), .Y(n_697) );
AND2x2_ASAP7_75t_L g716 ( .A(n_468), .B(n_606), .Y(n_716) );
AND2x2_ASAP7_75t_L g734 ( .A(n_468), .B(n_576), .Y(n_734) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
INVx1_ASAP7_75t_L g699 ( .A(n_477), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_493), .Y(n_477) );
AND2x2_ASAP7_75t_L g609 ( .A(n_478), .B(n_544), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_478), .B(n_629), .Y(n_628) );
AOI32xp33_ASAP7_75t_L g642 ( .A1(n_478), .A2(n_643), .A3(n_646), .B1(n_648), .B2(n_652), .Y(n_642) );
AND2x2_ASAP7_75t_L g712 ( .A(n_478), .B(n_606), .Y(n_712) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g576 ( .A(n_480), .B(n_545), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_480), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g618 ( .A(n_480), .B(n_565), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_480), .B(n_697), .Y(n_696) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_483), .B(n_491), .Y(n_480) );
INVx1_ASAP7_75t_L g581 ( .A(n_481), .Y(n_581) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_484), .A2(n_492), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g583 ( .A(n_493), .B(n_527), .Y(n_583) );
AND2x2_ASAP7_75t_L g659 ( .A(n_493), .B(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g731 ( .A(n_493), .Y(n_731) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
OR2x2_ASAP7_75t_L g526 ( .A(n_494), .B(n_504), .Y(n_526) );
AND2x2_ASAP7_75t_L g540 ( .A(n_494), .B(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_494), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g590 ( .A(n_494), .Y(n_590) );
AND2x2_ASAP7_75t_L g617 ( .A(n_494), .B(n_504), .Y(n_617) );
BUFx3_ASAP7_75t_L g620 ( .A(n_494), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_494), .B(n_595), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_494), .B(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g571 ( .A(n_503), .Y(n_571) );
AND2x2_ASAP7_75t_L g589 ( .A(n_503), .B(n_569), .Y(n_589) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g600 ( .A(n_504), .B(n_514), .Y(n_600) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_504), .Y(n_613) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_513), .B(n_620), .Y(n_670) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_SL g541 ( .A(n_514), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_514), .B(n_589), .C(n_590), .Y(n_588) );
OR2x2_ASAP7_75t_L g596 ( .A(n_514), .B(n_569), .Y(n_596) );
AND2x2_ASAP7_75t_L g616 ( .A(n_514), .B(n_569), .Y(n_616) );
AND2x2_ASAP7_75t_L g660 ( .A(n_514), .B(n_529), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_539), .B(n_542), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND2x2_ASAP7_75t_L g735 ( .A(n_525), .B(n_660), .Y(n_735) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_526), .A2(n_633), .B1(n_675), .B2(n_677), .Y(n_674) );
OR2x2_ASAP7_75t_L g681 ( .A(n_526), .B(n_596), .Y(n_681) );
OR2x2_ASAP7_75t_L g705 ( .A(n_526), .B(n_706), .Y(n_705) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_526), .B(n_625), .Y(n_718) );
AND2x2_ASAP7_75t_L g611 ( .A(n_527), .B(n_612), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_527), .A2(n_684), .B(n_699), .Y(n_698) );
AOI32xp33_ASAP7_75t_L g719 ( .A1(n_527), .A2(n_609), .A3(n_720), .B1(n_722), .B2(n_723), .Y(n_719) );
OR2x2_ASAP7_75t_L g730 ( .A(n_527), .B(n_731), .Y(n_730) );
CKINVDCx16_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g598 ( .A(n_528), .B(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_528), .B(n_612), .Y(n_677) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
AND2x2_ASAP7_75t_L g635 ( .A(n_529), .B(n_600), .Y(n_635) );
AND3x2_ASAP7_75t_L g644 ( .A(n_529), .B(n_540), .C(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g570 ( .A(n_541), .B(n_571), .Y(n_570) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_541), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_541), .B(n_569), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
AND2x2_ASAP7_75t_L g565 ( .A(n_543), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g605 ( .A(n_543), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g623 ( .A(n_543), .B(n_555), .Y(n_623) );
AND2x2_ASAP7_75t_L g641 ( .A(n_543), .B(n_545), .Y(n_641) );
OR2x2_ASAP7_75t_L g655 ( .A(n_543), .B(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g701 ( .A(n_543), .B(n_629), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_544), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_555), .Y(n_544) );
AND2x2_ASAP7_75t_L g602 ( .A(n_545), .B(n_580), .Y(n_602) );
OR2x2_ASAP7_75t_L g656 ( .A(n_545), .B(n_580), .Y(n_656) );
AND2x2_ASAP7_75t_L g709 ( .A(n_545), .B(n_566), .Y(n_709) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g607 ( .A(n_546), .Y(n_607) );
AND2x2_ASAP7_75t_L g629 ( .A(n_546), .B(n_555), .Y(n_629) );
INVx2_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
INVx1_ASAP7_75t_L g586 ( .A(n_555), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_567), .B(n_572), .C(n_584), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_565), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g728 ( .A(n_565), .Y(n_728) );
AND2x2_ASAP7_75t_L g606 ( .A(n_566), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_569), .B(n_570), .Y(n_578) );
INVx1_ASAP7_75t_L g663 ( .A(n_569), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_569), .B(n_590), .Y(n_687) );
AND2x2_ASAP7_75t_L g703 ( .A(n_569), .B(n_617), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_570), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g594 ( .A(n_571), .Y(n_594) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_578), .B1(n_579), .B2(n_582), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_575), .B(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_576), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g601 ( .A(n_577), .B(n_602), .Y(n_601) );
AOI221xp5_ASAP7_75t_SL g666 ( .A1(n_577), .A2(n_619), .B1(n_667), .B2(n_672), .C(n_674), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_577), .B(n_640), .Y(n_673) );
INVx1_ASAP7_75t_L g733 ( .A(n_579), .Y(n_733) );
BUFx3_ASAP7_75t_L g640 ( .A(n_580), .Y(n_640) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI21xp33_ASAP7_75t_SL g584 ( .A1(n_585), .A2(n_587), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_L g649 ( .A(n_586), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_586), .B(n_640), .Y(n_693) );
INVx1_ASAP7_75t_L g650 ( .A(n_587), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_587), .B(n_640), .Y(n_651) );
INVxp67_ASAP7_75t_L g671 ( .A(n_589), .Y(n_671) );
AND2x2_ASAP7_75t_L g612 ( .A(n_590), .B(n_613), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_597), .B(n_601), .C(n_603), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
INVx1_ASAP7_75t_SL g626 ( .A(n_594), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_595), .B(n_626), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_595), .B(n_617), .Y(n_668) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_598), .A2(n_604), .B1(n_608), .B2(n_610), .Y(n_603) );
INVx1_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g619 ( .A(n_600), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g664 ( .A(n_600), .B(n_665), .Y(n_664) );
OAI21xp33_ASAP7_75t_L g667 ( .A1(n_602), .A2(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_606), .A2(n_615), .B1(n_618), .B2(n_619), .C(n_621), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_606), .B(n_640), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_606), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g722 ( .A(n_612), .Y(n_722) );
INVxp67_ASAP7_75t_L g645 ( .A(n_613), .Y(n_645) );
INVx1_ASAP7_75t_L g652 ( .A(n_615), .Y(n_652) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g691 ( .A(n_616), .B(n_620), .Y(n_691) );
INVx1_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_620), .B(n_635), .Y(n_695) );
OAI32xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_624), .A3(n_626), .B1(n_627), .B2(n_628), .Y(n_621) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx2_ASAP7_75t_SL g634 ( .A(n_629), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_629), .B(n_661), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_629), .B(n_690), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g729 ( .A(n_629), .B(n_640), .Y(n_729) );
NAND5xp2_ASAP7_75t_L g630 ( .A(n_631), .B(n_653), .C(n_666), .D(n_678), .E(n_679), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_635), .B1(n_636), .B2(n_638), .C(n_642), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_637), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_640), .B(n_709), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_641), .A2(n_654), .B1(n_657), .B2(n_661), .Y(n_653) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_644), .A2(n_649), .B(n_650), .C(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g676 ( .A(n_656), .Y(n_676) );
INVx1_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_665), .B(n_714), .Y(n_724) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI222xp33_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_682), .B1(n_684), .B2(n_688), .C1(n_691), .C2(n_692), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_698), .B2(n_700), .C(n_702), .Y(n_694) );
INVx1_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B(n_707), .Y(n_702) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g714 ( .A(n_706), .Y(n_714) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g710 ( .A1(n_711), .A2(n_713), .B1(n_715), .B2(n_717), .C(n_719), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_729), .B(n_730), .C(n_732), .Y(n_725) );
INVxp67_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_735), .Y(n_732) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_738), .A2(n_741), .B1(n_742), .B2(n_743), .Y(n_740) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
endmodule