module fake_netlist_6_502_n_3131 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_3131);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_3131;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_1923;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_2977;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2672;
wire n_3030;
wire n_2291;
wire n_830;
wire n_2299;
wire n_461;
wire n_873;
wire n_1371;
wire n_2886;
wire n_2974;
wire n_1285;
wire n_1985;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_2982;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_544;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_836;
wire n_2074;
wire n_2447;
wire n_522;
wire n_2919;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_2739;
wire n_3023;
wire n_822;
wire n_693;
wire n_1313;
wire n_2791;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_3048;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3063;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_2703;
wire n_491;
wire n_2786;
wire n_1591;
wire n_772;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_2730;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_538;
wire n_3028;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3077;
wire n_1345;
wire n_1820;
wire n_2873;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_2880;
wire n_2394;
wire n_2108;
wire n_454;
wire n_1421;
wire n_2836;
wire n_1936;
wire n_1404;
wire n_638;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_3047;
wire n_1280;
wire n_713;
wire n_2655;
wire n_1400;
wire n_2625;
wire n_2843;
wire n_1467;
wire n_976;
wire n_3067;
wire n_2155;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2996;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_451;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_2907;
wire n_577;
wire n_2735;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_2850;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1309;
wire n_1123;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2633;
wire n_483;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_2073;
wire n_2273;
wire n_433;
wire n_2546;
wire n_792;
wire n_2522;
wire n_476;
wire n_2792;
wire n_1328;
wire n_1957;
wire n_2917;
wire n_2616;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_2811;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_2674;
wire n_2832;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_2831;
wire n_2998;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_2692;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_2908;
wire n_764;
wire n_2751;
wire n_2764;
wire n_1663;
wire n_2895;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_2922;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_2821;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_2459;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_715;
wire n_2678;
wire n_1251;
wire n_1265;
wire n_2711;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_674;
wire n_871;
wire n_3069;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_612;
wire n_2641;
wire n_3022;
wire n_3052;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2749;
wire n_2192;
wire n_2345;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_780;
wire n_675;
wire n_2624;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_2193;
wire n_2676;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2347;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_2916;
wire n_1063;
wire n_1588;
wire n_2963;
wire n_2947;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_2980;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_2733;
wire n_2824;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2812;
wire n_484;
wire n_2644;
wire n_2036;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_2687;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_2075;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_2763;
wire n_2762;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_3073;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_2078;
wire n_1634;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_2712;
wire n_2684;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_2691;
wire n_840;
wire n_2913;
wire n_874;
wire n_1756;
wire n_2493;
wire n_1128;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_2646;
wire n_1932;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_2631;
wire n_1364;
wire n_3078;
wire n_2436;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_2693;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_639;
wire n_963;
wire n_794;
wire n_2767;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_2707;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3037;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_2537;
wire n_2897;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_2747;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_2517;
wire n_2713;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_1788;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3018;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_3104;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_2717;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_425;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_3119;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_3129;
wire n_1849;
wire n_2848;
wire n_919;
wire n_2868;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_2857;
wire n_446;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_2896;
wire n_526;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2959;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_458;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_552;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3006;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_2424;
wire n_1604;
wire n_2296;
wire n_1284;
wire n_1142;
wire n_2849;
wire n_1475;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1398;
wire n_716;
wire n_884;
wire n_2354;
wire n_2682;
wire n_1201;
wire n_3032;
wire n_3103;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_474;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_2545;
wire n_889;
wire n_2432;
wire n_2710;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2788;
wire n_477;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2892;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_2748;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2475;
wire n_537;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_444;
wire n_3033;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_511;
wire n_2990;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1286;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_453;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_426;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_2502;
wire n_2801;
wire n_497;
wire n_2920;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_2306;
wire n_1614;
wire n_1892;
wire n_1459;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_2889;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_1243;
wire n_848;
wire n_2732;
wire n_2928;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_3109;
wire n_2023;
wire n_427;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_2863;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_2627;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_2993;
wire n_3016;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3004;
wire n_2830;
wire n_2781;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_1869;
wire n_664;
wire n_2911;
wire n_1764;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_2942;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_2851;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2841;
wire n_2420;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2656;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_2756;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_1549;
wire n_485;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_3120;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_2755;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_466;
wire n_2526;
wire n_3041;
wire n_2423;
wire n_1057;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_2636;
wire n_1818;
wire n_1108;
wire n_710;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_2740;
wire n_746;
wire n_1601;
wire n_609;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_1686;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_2716;
wire n_1320;
wire n_3081;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3010;
wire n_2499;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_2902;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_2988;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_2790;
wire n_2037;
wire n_2808;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_3040;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_2964;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2904;
wire n_2244;
wire n_3013;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_1642;
wire n_711;
wire n_1352;
wire n_579;
wire n_2789;
wire n_3105;
wire n_2872;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_456;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_2882;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_2782;
wire n_1974;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_2871;
wire n_420;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_3075;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_1343;
wire n_1522;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_799;
wire n_1548;
wire n_3044;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_2629;
wire n_1633;
wire n_2195;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_550;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2759;
wire n_2945;
wire n_3061;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2960;
wire n_3005;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_1706;
wire n_1498;
wire n_2653;
wire n_2417;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_502;
wire n_2668;
wire n_672;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_2840;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_3091;
wire n_834;
wire n_2695;
wire n_743;
wire n_766;
wire n_3124;
wire n_430;
wire n_1746;
wire n_1741;
wire n_1002;
wire n_1325;
wire n_1949;
wire n_545;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2888;
wire n_2793;
wire n_2715;
wire n_2885;
wire n_1804;
wire n_2923;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1600;
wire n_2833;
wire n_1113;
wire n_2253;
wire n_2758;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2978;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_2827;
wire n_1177;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1076;
wire n_1118;
wire n_2949;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_1377;
wire n_591;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_2587;
wire n_2931;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_2752;
wire n_1976;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2796;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2186;
wire n_2163;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3034;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_3083;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_2935;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_2702;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_1689;
wire n_2180;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_2117;
wire n_2234;
wire n_2779;
wire n_2685;
wire n_1083;
wire n_445;
wire n_1561;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_752;
wire n_908;
wire n_2649;
wire n_2721;
wire n_944;
wire n_2034;
wire n_1028;
wire n_576;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_2032;
wire n_2744;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_2743;
wire n_1973;
wire n_708;
wire n_2267;
wire n_3035;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_1266;
wire n_709;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_2934;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_2999;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_1582;
wire n_492;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_2950;
wire n_1972;
wire n_719;
wire n_3060;
wire n_2592;
wire n_1525;
wire n_3098;
wire n_2594;
wire n_455;
wire n_2666;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_3123;
wire n_2600;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_3130;
wire n_985;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_980;
wire n_2681;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_2047;
wire n_2651;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2799;
wire n_436;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_2742;
wire n_2640;
wire n_1051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_1996;
wire n_2367;
wire n_2867;
wire n_1039;
wire n_1442;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3116;
wire n_753;
wire n_1753;
wire n_3095;
wire n_2795;
wire n_2471;
wire n_467;
wire n_2540;
wire n_973;
wire n_2807;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_2968;
wire n_633;
wire n_1170;
wire n_1629;
wire n_665;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1632;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3001;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_2927;
wire n_1836;
wire n_2774;
wire n_3039;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_1322;
wire n_640;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_422;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_3079;
wire n_2098;
wire n_3085;
wire n_540;
wire n_2813;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_3070;
wire n_2223;
wire n_2091;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_2912;
wire n_2659;
wire n_2930;
wire n_1025;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_1259;
wire n_3054;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_84),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_310),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_154),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_33),
.Y(n_423)
);

BUFx10_ASAP7_75t_L g424 ( 
.A(n_138),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_79),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_316),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_107),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_169),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_28),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_109),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_399),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_342),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_93),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_144),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_292),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_364),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_25),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_23),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_155),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_303),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_414),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_59),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_5),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_38),
.Y(n_444)
);

BUFx2_ASAP7_75t_L g445 ( 
.A(n_37),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_282),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_107),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_220),
.Y(n_448)
);

BUFx10_ASAP7_75t_L g449 ( 
.A(n_289),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_243),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_223),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_346),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_249),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_251),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_367),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_197),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_184),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_57),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_75),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_31),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_180),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_253),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_106),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_403),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_55),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_10),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_190),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_283),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_276),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_53),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_311),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_325),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_103),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_275),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_397),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_213),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_308),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_49),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_301),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_157),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_321),
.Y(n_483)
);

INVx1_ASAP7_75t_SL g484 ( 
.A(n_383),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_216),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_262),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_235),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_109),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_158),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_56),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_354),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_417),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_214),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_400),
.Y(n_494)
);

BUFx5_ASAP7_75t_L g495 ( 
.A(n_349),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_168),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_11),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_96),
.Y(n_498)
);

INVx2_ASAP7_75t_SL g499 ( 
.A(n_211),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_322),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_73),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_84),
.Y(n_502)
);

BUFx10_ASAP7_75t_L g503 ( 
.A(n_208),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_183),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_304),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_336),
.Y(n_506)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_167),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_67),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_188),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_38),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_290),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_221),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_279),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_121),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_319),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_294),
.Y(n_516)
);

BUFx10_ASAP7_75t_L g517 ( 
.A(n_401),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_185),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_418),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_97),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_247),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_411),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_35),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_281),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_124),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_160),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_233),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_82),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_88),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_102),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_80),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_390),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_25),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_74),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_309),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_259),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_340),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_395),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_131),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_24),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_23),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_234),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_22),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_402),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_207),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_407),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_119),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_205),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_146),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_405),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_185),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_284),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_143),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_327),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_344),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_237),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_248),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_114),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_181),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_419),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_370),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_416),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_317),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_330),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_89),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_100),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_217),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_199),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_45),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_218),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_74),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_320),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_226),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_111),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_246),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_170),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_396),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_298),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_134),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_339),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_348),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_229),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_356),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_271),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_160),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_98),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_141),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_134),
.Y(n_588)
);

BUFx2_ASAP7_75t_R g589 ( 
.A(n_73),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_90),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_28),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_274),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_186),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_203),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_77),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_184),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_183),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_347),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_33),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_124),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_362),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_166),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_338),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_258),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_100),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_116),
.Y(n_606)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_337),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_355),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_57),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_34),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_187),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_149),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_17),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_369),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_102),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_94),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_192),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_68),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_195),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_156),
.Y(n_620)
);

CKINVDCx16_ASAP7_75t_R g621 ( 
.A(n_291),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_105),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_138),
.Y(n_623)
);

CKINVDCx14_ASAP7_75t_R g624 ( 
.A(n_412),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_263),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_231),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_384),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_410),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_269),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_288),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_97),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_191),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_225),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_328),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_161),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_191),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_215),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_55),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_324),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_227),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_4),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_368),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_60),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_238),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_93),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_270),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_190),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_114),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_164),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_106),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_111),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_168),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_228),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_267),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_131),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_105),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_94),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_273),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_104),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_118),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_122),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_165),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_155),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_157),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_127),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_314),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_76),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_61),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_76),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_37),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_296),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_56),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_198),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_239),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_126),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_252),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_103),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_256),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_389),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_312),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_358),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_171),
.Y(n_682)
);

CKINVDCx20_ASAP7_75t_R g683 ( 
.A(n_387),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_194),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_148),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_302),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_27),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_137),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_135),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_112),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_141),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_386),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_29),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_140),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_132),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_19),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_83),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_41),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_153),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_108),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_115),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_48),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_2),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_35),
.Y(n_704)
);

BUFx10_ASAP7_75t_L g705 ( 
.A(n_49),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_350),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_209),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_334),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_2),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_318),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_286),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_326),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_385),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_17),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_332),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_224),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_22),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_158),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_232),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_40),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_261),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_177),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_187),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_152),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_31),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_52),
.Y(n_726)
);

CKINVDCx16_ASAP7_75t_R g727 ( 
.A(n_431),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_695),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_446),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_695),
.Y(n_730)
);

INVxp67_ASAP7_75t_SL g731 ( 
.A(n_537),
.Y(n_731)
);

CKINVDCx16_ASAP7_75t_R g732 ( 
.A(n_431),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_695),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_695),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_420),
.Y(n_735)
);

CKINVDCx20_ASAP7_75t_R g736 ( 
.A(n_486),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_492),
.B(n_0),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_695),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_695),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_695),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_695),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_560),
.B(n_0),
.Y(n_742)
);

INVxp33_ASAP7_75t_L g743 ( 
.A(n_702),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_437),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_537),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_437),
.Y(n_746)
);

BUFx3_ASAP7_75t_L g747 ( 
.A(n_568),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_437),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_437),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_437),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_422),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_425),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_518),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_518),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_568),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_518),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_518),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_518),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_427),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_445),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_525),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_429),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_525),
.Y(n_763)
);

INVxp33_ASAP7_75t_SL g764 ( 
.A(n_445),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_525),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_673),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_525),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_525),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_673),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_434),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_434),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_460),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_527),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_460),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_482),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_421),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_482),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_553),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_558),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_436),
.Y(n_780)
);

INVxp33_ASAP7_75t_SL g781 ( 
.A(n_558),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_436),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_455),
.Y(n_783)
);

INVxp67_ASAP7_75t_SL g784 ( 
.A(n_560),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_455),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_492),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_458),
.Y(n_787)
);

INVxp33_ASAP7_75t_SL g788 ( 
.A(n_430),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_458),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_495),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_476),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_470),
.B(n_1),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_476),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_481),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_481),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_483),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_483),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_487),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_487),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_506),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_506),
.Y(n_801)
);

BUFx5_ASAP7_75t_L g802 ( 
.A(n_516),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_516),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_438),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_524),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_524),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_495),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_442),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_443),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_555),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_555),
.Y(n_811)
);

INVxp33_ASAP7_75t_SL g812 ( 
.A(n_444),
.Y(n_812)
);

INVxp33_ASAP7_75t_SL g813 ( 
.A(n_461),
.Y(n_813)
);

INVxp33_ASAP7_75t_SL g814 ( 
.A(n_462),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_562),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_562),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_449),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_449),
.Y(n_818)
);

INVxp67_ASAP7_75t_SL g819 ( 
.A(n_560),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_570),
.Y(n_820)
);

INVxp33_ASAP7_75t_SL g821 ( 
.A(n_463),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_467),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_439),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_570),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_575),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_468),
.Y(n_826)
);

HB1xp67_ASAP7_75t_L g827 ( 
.A(n_475),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_603),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_575),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_581),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_581),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_584),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_584),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_592),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_449),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_495),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_480),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_592),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_L g839 ( 
.A(n_534),
.B(n_1),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_598),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_598),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_614),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_424),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_614),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_625),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_424),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_625),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_502),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_553),
.Y(n_849)
);

INVxp33_ASAP7_75t_SL g850 ( 
.A(n_488),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_588),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_588),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_495),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_659),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_489),
.Y(n_855)
);

INVxp67_ASAP7_75t_SL g856 ( 
.A(n_607),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_659),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_497),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_660),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_660),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_497),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_698),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_698),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_498),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_509),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_744),
.Y(n_866)
);

BUFx6f_ASAP7_75t_L g867 ( 
.A(n_758),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_744),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_758),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_746),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_861),
.B(n_731),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_L g872 ( 
.A1(n_764),
.A2(n_508),
.B1(n_539),
.B2(n_528),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_735),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_768),
.Y(n_874)
);

INVx5_ASAP7_75t_L g875 ( 
.A(n_776),
.Y(n_875)
);

BUFx6f_ASAP7_75t_L g876 ( 
.A(n_768),
.Y(n_876)
);

INVxp67_ASAP7_75t_L g877 ( 
.A(n_827),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_760),
.Y(n_878)
);

OAI22x1_ASAP7_75t_SL g879 ( 
.A1(n_764),
.A2(n_595),
.B1(n_597),
.B2(n_543),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_735),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_748),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_788),
.B(n_808),
.Y(n_883)
);

BUFx2_ASAP7_75t_L g884 ( 
.A(n_751),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_748),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_784),
.B(n_470),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_781),
.A2(n_690),
.B1(n_599),
.B2(n_520),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_745),
.B(n_624),
.Y(n_888)
);

AND2x6_ASAP7_75t_L g889 ( 
.A(n_728),
.B(n_421),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_819),
.B(n_499),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_749),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_776),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_856),
.B(n_499),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_749),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_750),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_750),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_753),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_747),
.B(n_501),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_742),
.B(n_583),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_728),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_753),
.Y(n_901)
);

HB1xp67_ASAP7_75t_L g902 ( 
.A(n_751),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_754),
.B(n_583),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_754),
.B(n_756),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_730),
.A2(n_706),
.B(n_686),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_747),
.B(n_686),
.Y(n_906)
);

AND2x4_ASAP7_75t_L g907 ( 
.A(n_756),
.B(n_706),
.Y(n_907)
);

INVx5_ASAP7_75t_L g908 ( 
.A(n_776),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_757),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_757),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_755),
.B(n_426),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_761),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_761),
.Y(n_913)
);

BUFx3_ASAP7_75t_L g914 ( 
.A(n_755),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_766),
.B(n_501),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_752),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_766),
.B(n_432),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_823),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_769),
.B(n_435),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_752),
.Y(n_920)
);

AND2x2_ASAP7_75t_SL g921 ( 
.A(n_792),
.B(n_621),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_733),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_763),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_763),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_759),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_765),
.Y(n_927)
);

BUFx2_ASAP7_75t_L g928 ( 
.A(n_759),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_765),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_767),
.Y(n_930)
);

INVx4_ASAP7_75t_L g931 ( 
.A(n_802),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_790),
.Y(n_932)
);

XOR2xp5_ASAP7_75t_L g933 ( 
.A(n_729),
.B(n_589),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_767),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_769),
.B(n_858),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_858),
.B(n_507),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_781),
.A2(n_565),
.B1(n_621),
.B2(n_683),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_738),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_737),
.A2(n_715),
.B1(n_523),
.B2(n_529),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_739),
.A2(n_629),
.B(n_627),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_740),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_780),
.B(n_627),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_782),
.B(n_629),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_741),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_783),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_802),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_790),
.Y(n_947)
);

INVx3_ASAP7_75t_L g948 ( 
.A(n_807),
.Y(n_948)
);

OAI22x1_ASAP7_75t_SL g949 ( 
.A1(n_848),
.A2(n_428),
.B1(n_433),
.B2(n_423),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_785),
.Y(n_950)
);

AND2x4_ASAP7_75t_L g951 ( 
.A(n_787),
.B(n_639),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_789),
.Y(n_952)
);

BUFx12f_ASAP7_75t_L g953 ( 
.A(n_762),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_791),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_793),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_794),
.B(n_795),
.Y(n_956)
);

INVxp33_ASAP7_75t_SL g957 ( 
.A(n_762),
.Y(n_957)
);

AND2x2_ASAP7_75t_SL g958 ( 
.A(n_727),
.B(n_639),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_770),
.Y(n_959)
);

BUFx12f_ASAP7_75t_L g960 ( 
.A(n_804),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_804),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_796),
.Y(n_962)
);

BUFx8_ASAP7_75t_SL g963 ( 
.A(n_760),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_802),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_797),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_798),
.B(n_507),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_817),
.B(n_440),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_799),
.Y(n_968)
);

INVx3_ASAP7_75t_L g969 ( 
.A(n_836),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_817),
.Y(n_970)
);

AND2x4_ASAP7_75t_L g971 ( 
.A(n_800),
.B(n_666),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_770),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_809),
.Y(n_973)
);

AOI22x1_ASAP7_75t_SL g974 ( 
.A1(n_736),
.A2(n_828),
.B1(n_773),
.B2(n_531),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_771),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_788),
.B(n_484),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_732),
.B(n_786),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_801),
.B(n_611),
.Y(n_978)
);

OAI21x1_ASAP7_75t_L g979 ( 
.A1(n_853),
.A2(n_671),
.B(n_666),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_853),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_802),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_803),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_878),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_916),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_938),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_885),
.Y(n_987)
);

BUFx8_ASAP7_75t_L g988 ( 
.A(n_916),
.Y(n_988)
);

BUFx6f_ASAP7_75t_SL g989 ( 
.A(n_958),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_914),
.B(n_805),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_R g991 ( 
.A(n_953),
.B(n_809),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_914),
.B(n_806),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_938),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_885),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_976),
.B(n_808),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_871),
.B(n_936),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_953),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_941),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_R g999 ( 
.A(n_960),
.B(n_822),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_SL g1000 ( 
.A1(n_937),
.A2(n_813),
.B1(n_814),
.B2(n_812),
.Y(n_1000)
);

BUFx8_ASAP7_75t_L g1001 ( 
.A(n_960),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_941),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_957),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_944),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_911),
.B(n_812),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_944),
.Y(n_1007)
);

BUFx2_ASAP7_75t_L g1008 ( 
.A(n_963),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_954),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_954),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_973),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_891),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_954),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_973),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_914),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_940),
.A2(n_811),
.B(n_810),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_878),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_955),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_955),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_974),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_878),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_955),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_974),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_878),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_898),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_881),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_881),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_871),
.B(n_822),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_940),
.A2(n_816),
.B(n_815),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_936),
.B(n_826),
.Y(n_1030)
);

CKINVDCx11_ASAP7_75t_R g1031 ( 
.A(n_884),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_SL g1032 ( 
.A(n_921),
.B(n_813),
.Y(n_1032)
);

CKINVDCx20_ASAP7_75t_R g1033 ( 
.A(n_933),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_982),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_982),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_898),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_982),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_886),
.B(n_802),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_884),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_956),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_891),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_942),
.B(n_820),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_915),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_956),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_932),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_933),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_894),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_956),
.Y(n_1048)
);

BUFx3_ASAP7_75t_L g1049 ( 
.A(n_915),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_945),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_894),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_886),
.B(n_824),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_956),
.Y(n_1053)
);

INVx3_ASAP7_75t_L g1054 ( 
.A(n_932),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_928),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_896),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_886),
.B(n_825),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_945),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_932),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_886),
.B(n_829),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_945),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_945),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_945),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_928),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_950),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_950),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_947),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_896),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_879),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_879),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_873),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_970),
.B(n_826),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_901),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_950),
.Y(n_1074)
);

CKINVDCx20_ASAP7_75t_R g1075 ( 
.A(n_872),
.Y(n_1075)
);

INVxp67_ASAP7_75t_L g1076 ( 
.A(n_883),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_950),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_902),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_920),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_926),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_888),
.B(n_830),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_947),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_947),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_889),
.B(n_495),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_921),
.B(n_814),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_952),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_961),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_952),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_952),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_R g1090 ( 
.A(n_970),
.B(n_837),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_952),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_952),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_947),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_962),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_877),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_942),
.B(n_831),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_966),
.B(n_837),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_967),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_901),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_979),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_917),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_962),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_948),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_962),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_919),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_872),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_927),
.Y(n_1107)
);

BUFx8_ASAP7_75t_L g1108 ( 
.A(n_966),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_962),
.Y(n_1109)
);

CKINVDCx14_ASAP7_75t_R g1110 ( 
.A(n_937),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_905),
.A2(n_833),
.B(n_832),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_978),
.B(n_855),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_962),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_958),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_958),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_939),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_978),
.B(n_855),
.Y(n_1117)
);

INVxp67_ASAP7_75t_L g1118 ( 
.A(n_935),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_965),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

CKINVDCx16_ASAP7_75t_R g1121 ( 
.A(n_939),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_965),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_965),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_942),
.B(n_943),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_949),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_965),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_927),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_968),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_949),
.Y(n_1129)
);

INVx3_ASAP7_75t_L g1130 ( 
.A(n_948),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_968),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_968),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_929),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_905),
.A2(n_838),
.B(n_834),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_942),
.B(n_943),
.Y(n_1135)
);

INVxp67_ASAP7_75t_L g1136 ( 
.A(n_893),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_SL g1137 ( 
.A(n_921),
.B(n_821),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_887),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_929),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_887),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_968),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_968),
.Y(n_1142)
);

CKINVDCx20_ASAP7_75t_R g1143 ( 
.A(n_977),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_922),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_934),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_922),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_934),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_922),
.Y(n_1148)
);

BUFx6f_ASAP7_75t_L g1149 ( 
.A(n_867),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_899),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_996),
.B(n_943),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1136),
.B(n_943),
.Y(n_1152)
);

AND2x2_ASAP7_75t_SL g1153 ( 
.A(n_1121),
.B(n_899),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1040),
.Y(n_1154)
);

INVx3_ASAP7_75t_L g1155 ( 
.A(n_1100),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_L g1156 ( 
.A(n_1076),
.B(n_821),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1100),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1038),
.B(n_890),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_987),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1036),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1124),
.A2(n_899),
.B1(n_971),
.B2(n_951),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1124),
.B(n_900),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1118),
.B(n_850),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_1124),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_SL g1165 ( 
.A(n_1135),
.B(n_900),
.Y(n_1165)
);

XOR2xp5_ASAP7_75t_L g1166 ( 
.A(n_985),
.B(n_864),
.Y(n_1166)
);

NAND2xp33_ASAP7_75t_SL g1167 ( 
.A(n_1116),
.B(n_1150),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_987),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_994),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1101),
.B(n_899),
.Y(n_1170)
);

INVx4_ASAP7_75t_L g1171 ( 
.A(n_1050),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_991),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1135),
.B(n_1150),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1003),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_994),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1025),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1044),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1048),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1053),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1012),
.Y(n_1180)
);

BUFx10_ASAP7_75t_L g1181 ( 
.A(n_1004),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1012),
.Y(n_1182)
);

BUFx4f_ASAP7_75t_L g1183 ( 
.A(n_1135),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1041),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1039),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1041),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1105),
.B(n_900),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1036),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1047),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1098),
.B(n_900),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1047),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1081),
.B(n_986),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1028),
.B(n_892),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_999),
.Y(n_1194)
);

INVx4_ASAP7_75t_L g1195 ( 
.A(n_1050),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_995),
.B(n_850),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1049),
.Y(n_1197)
);

AND3x2_ASAP7_75t_L g1198 ( 
.A(n_1008),
.B(n_689),
.C(n_779),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1049),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1042),
.A2(n_951),
.B1(n_971),
.B2(n_889),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_993),
.B(n_892),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_985),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1043),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1009),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_990),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1051),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1010),
.Y(n_1207)
);

INVx2_ASAP7_75t_SL g1208 ( 
.A(n_990),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1013),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1018),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1019),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1022),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1034),
.Y(n_1213)
);

INVx1_ASAP7_75t_SL g1214 ( 
.A(n_1095),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1035),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_990),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1032),
.A2(n_835),
.B1(n_818),
.B2(n_864),
.Y(n_1217)
);

NAND3xp33_ASAP7_75t_L g1218 ( 
.A(n_1116),
.B(n_865),
.C(n_906),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1026),
.Y(n_1219)
);

NOR2xp33_ASAP7_75t_L g1220 ( 
.A(n_1006),
.B(n_865),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1042),
.A2(n_951),
.B1(n_971),
.B2(n_889),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_998),
.B(n_892),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1037),
.Y(n_1223)
);

INVx4_ASAP7_75t_L g1224 ( 
.A(n_1050),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1050),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1097),
.B(n_843),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_992),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_1134),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1042),
.A2(n_951),
.B1(n_971),
.B2(n_889),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1002),
.B(n_892),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_SL g1231 ( 
.A(n_1137),
.B(n_924),
.Y(n_1231)
);

INVxp33_ASAP7_75t_L g1232 ( 
.A(n_1090),
.Y(n_1232)
);

INVxp33_ASAP7_75t_L g1233 ( 
.A(n_1030),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1005),
.B(n_924),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_992),
.Y(n_1235)
);

AND2x6_ASAP7_75t_L g1236 ( 
.A(n_1072),
.B(n_671),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1051),
.Y(n_1237)
);

AO21x2_ASAP7_75t_L g1238 ( 
.A1(n_1085),
.A2(n_1062),
.B(n_1058),
.Y(n_1238)
);

OR2x2_ASAP7_75t_L g1239 ( 
.A(n_1112),
.B(n_846),
.Y(n_1239)
);

NOR3xp33_ASAP7_75t_L g1240 ( 
.A(n_1000),
.B(n_839),
.C(n_835),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_992),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1117),
.B(n_818),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_L g1243 ( 
.A(n_1052),
.B(n_495),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1056),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1111),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1007),
.B(n_924),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1015),
.B(n_743),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1111),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1057),
.B(n_1060),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1056),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1096),
.B(n_946),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1134),
.Y(n_1252)
);

INVx4_ASAP7_75t_L g1253 ( 
.A(n_1061),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1068),
.Y(n_1254)
);

AND3x2_ASAP7_75t_L g1255 ( 
.A(n_1078),
.B(n_428),
.C(n_423),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1068),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1096),
.B(n_946),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1096),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1016),
.B(n_681),
.Y(n_1259)
);

AND2x4_ASAP7_75t_SL g1260 ( 
.A(n_984),
.B(n_503),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1073),
.Y(n_1261)
);

NAND3xp33_ASAP7_75t_L g1262 ( 
.A(n_1114),
.B(n_533),
.C(n_526),
.Y(n_1262)
);

BUFx8_ASAP7_75t_SL g1263 ( 
.A(n_1033),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1061),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1073),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1079),
.B(n_959),
.Y(n_1266)
);

INVx4_ASAP7_75t_L g1267 ( 
.A(n_1061),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1108),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1045),
.B(n_931),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_L g1270 ( 
.A(n_1115),
.B(n_541),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1115),
.B(n_547),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_1055),
.B(n_549),
.Y(n_1272)
);

AOI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_989),
.A2(n_448),
.B1(n_450),
.B2(n_441),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1144),
.B(n_681),
.Y(n_1274)
);

AND2x2_ASAP7_75t_SL g1275 ( 
.A(n_1084),
.B(n_692),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1099),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1016),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1029),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1099),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1029),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_1108),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1045),
.Y(n_1282)
);

AND2x4_ASAP7_75t_L g1283 ( 
.A(n_1054),
.B(n_692),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1061),
.Y(n_1284)
);

INVx4_ASAP7_75t_L g1285 ( 
.A(n_1074),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1107),
.Y(n_1286)
);

INVx3_ASAP7_75t_L g1287 ( 
.A(n_1054),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1059),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_989),
.A2(n_452),
.B1(n_453),
.B2(n_451),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_1108),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_SL g1291 ( 
.A(n_1059),
.B(n_931),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1149),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1067),
.B(n_964),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1138),
.B(n_504),
.Y(n_1294)
);

AND2x6_ASAP7_75t_L g1295 ( 
.A(n_1146),
.B(n_712),
.Y(n_1295)
);

INVxp33_ASAP7_75t_SL g1296 ( 
.A(n_1026),
.Y(n_1296)
);

INVx3_ASAP7_75t_L g1297 ( 
.A(n_1067),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1082),
.B(n_981),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1082),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1082),
.B(n_959),
.Y(n_1300)
);

AND2x4_ASAP7_75t_L g1301 ( 
.A(n_1083),
.B(n_712),
.Y(n_1301)
);

BUFx3_ASAP7_75t_L g1302 ( 
.A(n_988),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1027),
.B(n_424),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1107),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1083),
.B(n_495),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_988),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1127),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1083),
.Y(n_1308)
);

NOR2x1p5_ASAP7_75t_L g1309 ( 
.A(n_1024),
.B(n_611),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1093),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1148),
.A2(n_889),
.B1(n_907),
.B2(n_903),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1127),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1093),
.Y(n_1313)
);

NOR2xp33_ASAP7_75t_L g1314 ( 
.A(n_1138),
.B(n_551),
.Y(n_1314)
);

AND3x2_ASAP7_75t_L g1315 ( 
.A(n_1110),
.B(n_447),
.C(n_433),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1140),
.B(n_504),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1133),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_988),
.Y(n_1318)
);

HB1xp67_ASAP7_75t_L g1319 ( 
.A(n_1027),
.Y(n_1319)
);

AND2x4_ASAP7_75t_L g1320 ( 
.A(n_1093),
.B(n_979),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1103),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1103),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1103),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1130),
.A2(n_889),
.B1(n_907),
.B2(n_903),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1133),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1149),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1130),
.Y(n_1327)
);

NAND3xp33_ASAP7_75t_L g1328 ( 
.A(n_1140),
.B(n_569),
.C(n_566),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1074),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1130),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1139),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1139),
.Y(n_1332)
);

OR2x6_ASAP7_75t_L g1333 ( 
.A(n_989),
.B(n_590),
.Y(n_1333)
);

BUFx10_ASAP7_75t_L g1334 ( 
.A(n_997),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1145),
.Y(n_1335)
);

BUFx3_ASAP7_75t_L g1336 ( 
.A(n_1174),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1300),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1300),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1159),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1154),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1266),
.B(n_1064),
.Y(n_1341)
);

AND2x4_ASAP7_75t_SL g1342 ( 
.A(n_1181),
.B(n_984),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1177),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1151),
.B(n_1145),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1178),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1263),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1159),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1179),
.Y(n_1348)
);

INVxp33_ASAP7_75t_L g1349 ( 
.A(n_1247),
.Y(n_1349)
);

OAI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1275),
.A2(n_1110),
.B1(n_1106),
.B2(n_1075),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1164),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1168),
.Y(n_1352)
);

OA22x2_ASAP7_75t_L g1353 ( 
.A1(n_1315),
.A2(n_1129),
.B1(n_1125),
.B2(n_1064),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1160),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1164),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1164),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1288),
.Y(n_1357)
);

INVx8_ASAP7_75t_L g1358 ( 
.A(n_1236),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_1263),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1308),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1157),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1310),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1266),
.B(n_1071),
.Y(n_1363)
);

NAND2x1p5_ASAP7_75t_L g1364 ( 
.A(n_1183),
.B(n_1074),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1151),
.B(n_1147),
.Y(n_1365)
);

INVx4_ASAP7_75t_L g1366 ( 
.A(n_1199),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1321),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1322),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1160),
.Y(n_1369)
);

AO22x2_ASAP7_75t_L g1370 ( 
.A1(n_1231),
.A2(n_590),
.B1(n_459),
.B2(n_465),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1220),
.B(n_1071),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1323),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1330),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1199),
.Y(n_1374)
);

OAI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1196),
.A2(n_1087),
.B(n_1080),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1332),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1335),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1168),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1169),
.Y(n_1379)
);

INVx4_ASAP7_75t_L g1380 ( 
.A(n_1199),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1249),
.B(n_1147),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1166),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1169),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1175),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1175),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1233),
.B(n_1080),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1183),
.B(n_1074),
.Y(n_1387)
);

AND2x6_ASAP7_75t_L g1388 ( 
.A(n_1155),
.B(n_1063),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1180),
.Y(n_1389)
);

AND2x4_ASAP7_75t_L g1390 ( 
.A(n_1216),
.B(n_1143),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1163),
.B(n_1087),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1172),
.Y(n_1392)
);

BUFx2_ASAP7_75t_L g1393 ( 
.A(n_1185),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1157),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1214),
.Y(n_1395)
);

INVxp67_ASAP7_75t_L g1396 ( 
.A(n_1152),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1216),
.B(n_1143),
.Y(n_1397)
);

AOI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1193),
.A2(n_1106),
.B1(n_1075),
.B2(n_1066),
.Y(n_1398)
);

AND2x2_ASAP7_75t_SL g1399 ( 
.A(n_1275),
.B(n_1084),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1180),
.Y(n_1400)
);

AND2x4_ASAP7_75t_L g1401 ( 
.A(n_1235),
.B(n_972),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1242),
.B(n_1014),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1182),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1172),
.Y(n_1404)
);

NAND3xp33_ASAP7_75t_L g1405 ( 
.A(n_1314),
.B(n_1129),
.C(n_1125),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1235),
.B(n_972),
.Y(n_1406)
);

NOR2xp33_ASAP7_75t_L g1407 ( 
.A(n_1233),
.B(n_1156),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1157),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1232),
.B(n_1024),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1258),
.B(n_1188),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1236),
.A2(n_459),
.B1(n_465),
.B2(n_447),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1249),
.B(n_1158),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1158),
.B(n_1192),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1187),
.B(n_1065),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1182),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1184),
.Y(n_1416)
);

BUFx6f_ASAP7_75t_L g1417 ( 
.A(n_1157),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1184),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1186),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1152),
.B(n_1031),
.Y(n_1420)
);

OR2x6_ASAP7_75t_L g1421 ( 
.A(n_1306),
.B(n_1001),
.Y(n_1421)
);

BUFx6f_ASAP7_75t_L g1422 ( 
.A(n_1199),
.Y(n_1422)
);

AND2x6_ASAP7_75t_L g1423 ( 
.A(n_1155),
.B(n_1077),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1186),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1181),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1189),
.Y(n_1426)
);

INVx5_ASAP7_75t_L g1427 ( 
.A(n_1155),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1189),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_1176),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1191),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1191),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1206),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_L g1433 ( 
.A(n_1270),
.B(n_1031),
.C(n_1011),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1206),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1181),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1237),
.Y(n_1436)
);

NAND3xp33_ASAP7_75t_L g1437 ( 
.A(n_1271),
.B(n_1011),
.C(n_997),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1237),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1203),
.Y(n_1439)
);

XNOR2xp5_ASAP7_75t_L g1440 ( 
.A(n_1153),
.B(n_1017),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1244),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1193),
.A2(n_1086),
.B1(n_1089),
.B2(n_1088),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1232),
.B(n_1226),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1287),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1231),
.A2(n_1102),
.B1(n_1104),
.B2(n_1094),
.Y(n_1445)
);

NAND3xp33_ASAP7_75t_L g1446 ( 
.A(n_1272),
.B(n_1070),
.C(n_1069),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1287),
.Y(n_1447)
);

INVx5_ASAP7_75t_L g1448 ( 
.A(n_1292),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_L g1449 ( 
.A(n_1183),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1194),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1190),
.B(n_1091),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1292),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1170),
.B(n_1091),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1171),
.B(n_1091),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1292),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1197),
.B(n_975),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1244),
.Y(n_1457)
);

OR2x2_ASAP7_75t_SL g1458 ( 
.A(n_1328),
.B(n_1069),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1292),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1228),
.B(n_1109),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1205),
.B(n_975),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1250),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1250),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1161),
.A2(n_472),
.B1(n_490),
.B2(n_469),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1254),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1219),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1326),
.Y(n_1467)
);

BUFx3_ASAP7_75t_L g1468 ( 
.A(n_1306),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1254),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1239),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1319),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1256),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1228),
.B(n_1119),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1256),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1261),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1261),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1205),
.B(n_983),
.Y(n_1477)
);

AO22x2_ASAP7_75t_L g1478 ( 
.A1(n_1294),
.A2(n_472),
.B1(n_490),
.B2(n_469),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1252),
.B(n_1120),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1306),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1265),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1296),
.A2(n_1046),
.B1(n_1033),
.B2(n_1070),
.Y(n_1482)
);

AND2x6_ASAP7_75t_L g1483 ( 
.A(n_1252),
.B(n_1122),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1303),
.B(n_1017),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1153),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1316),
.B(n_1021),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1371),
.A2(n_1407),
.B1(n_1167),
.B2(n_1391),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_SL g1488 ( 
.A(n_1399),
.B(n_1167),
.Y(n_1488)
);

AOI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1371),
.A2(n_1173),
.B1(n_1218),
.B2(n_1262),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1340),
.Y(n_1490)
);

AND2x6_ASAP7_75t_SL g1491 ( 
.A(n_1421),
.B(n_1333),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1399),
.B(n_1208),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1363),
.B(n_1217),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_L g1494 ( 
.A(n_1358),
.B(n_1236),
.Y(n_1494)
);

NAND2x1p5_ASAP7_75t_L g1495 ( 
.A(n_1449),
.B(n_1208),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1413),
.B(n_1236),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1343),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1413),
.B(n_1236),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1339),
.Y(n_1499)
);

INVx2_ASAP7_75t_SL g1500 ( 
.A(n_1336),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1449),
.B(n_1251),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1427),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1347),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1349),
.B(n_1296),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1345),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1449),
.B(n_1257),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1407),
.A2(n_1386),
.B1(n_1396),
.B2(n_1173),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1396),
.B(n_1236),
.Y(n_1508)
);

AND2x6_ASAP7_75t_SL g1509 ( 
.A(n_1421),
.B(n_1333),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1337),
.A2(n_1241),
.B(n_1227),
.C(n_1204),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1410),
.A2(n_1209),
.B1(n_1210),
.B2(n_1207),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1395),
.B(n_1333),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1348),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1338),
.B(n_1211),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1352),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1361),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1341),
.B(n_1333),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1461),
.B(n_1212),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1461),
.B(n_1213),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1477),
.B(n_1215),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1470),
.B(n_1393),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1427),
.B(n_1287),
.Y(n_1522)
);

AOI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1386),
.A2(n_1273),
.B1(n_1289),
.B2(n_1223),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1477),
.B(n_1283),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1378),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1412),
.B(n_1283),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1412),
.B(n_1283),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1383),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1379),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1414),
.B(n_1301),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1414),
.B(n_1301),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1344),
.B(n_1301),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1384),
.Y(n_1533)
);

NOR2x1p5_ASAP7_75t_L g1534 ( 
.A(n_1468),
.B(n_1302),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1361),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_L g1536 ( 
.A1(n_1453),
.A2(n_1259),
.B(n_1245),
.C(n_1248),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1350),
.B(n_1202),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1349),
.B(n_1194),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_SL g1539 ( 
.A(n_1427),
.B(n_1297),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1366),
.B(n_1171),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1344),
.B(n_1297),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1365),
.B(n_1297),
.Y(n_1542)
);

NAND2xp33_ASAP7_75t_L g1543 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1400),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1385),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_1427),
.B(n_1299),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1365),
.B(n_1313),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1356),
.B(n_1299),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1410),
.A2(n_1165),
.B1(n_1162),
.B2(n_1238),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1411),
.A2(n_1165),
.B1(n_1162),
.B2(n_1238),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1366),
.B(n_1171),
.Y(n_1551)
);

AND2x2_ASAP7_75t_SL g1552 ( 
.A(n_1411),
.B(n_1240),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1443),
.B(n_1485),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1389),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1401),
.A2(n_1238),
.B1(n_1221),
.B2(n_1229),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1401),
.B(n_1327),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1398),
.A2(n_1243),
.B1(n_1309),
.B2(n_1200),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1406),
.A2(n_1243),
.B1(n_1295),
.B2(n_1274),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1406),
.B(n_1327),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1350),
.B(n_1202),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1361),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1370),
.B(n_1327),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1336),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_1450),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1370),
.A2(n_1295),
.B1(n_1274),
.B2(n_1246),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_SL g1566 ( 
.A(n_1359),
.B(n_1021),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1356),
.B(n_1299),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1403),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_1359),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1415),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1466),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1351),
.A2(n_1355),
.B1(n_1447),
.B2(n_1444),
.Y(n_1572)
);

BUFx4f_ASAP7_75t_L g1573 ( 
.A(n_1425),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_SL g1574 ( 
.A1(n_1382),
.A2(n_1046),
.B1(n_1482),
.B2(n_1023),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1381),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1499),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_R g1577 ( 
.A(n_1564),
.B(n_1392),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1487),
.B(n_1375),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1569),
.Y(n_1579)
);

INVx3_ASAP7_75t_L g1580 ( 
.A(n_1502),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_1569),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_R g1582 ( 
.A(n_1538),
.B(n_1392),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1552),
.A2(n_1464),
.B1(n_1488),
.B2(n_1370),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1521),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1504),
.B(n_1429),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_SL g1586 ( 
.A(n_1534),
.B(n_1404),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1499),
.Y(n_1587)
);

OR2x6_ASAP7_75t_L g1588 ( 
.A(n_1492),
.B(n_1358),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1503),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1503),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1515),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1354),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1488),
.B(n_1381),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1573),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1531),
.B(n_1376),
.Y(n_1595)
);

NOR2x1_ASAP7_75t_R g1596 ( 
.A(n_1571),
.B(n_1404),
.Y(n_1596)
);

INVx3_ASAP7_75t_L g1597 ( 
.A(n_1502),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_R g1598 ( 
.A(n_1573),
.B(n_1346),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1552),
.B(n_1444),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1507),
.B(n_1390),
.Y(n_1600)
);

CKINVDCx6p67_ASAP7_75t_R g1601 ( 
.A(n_1563),
.Y(n_1601)
);

OR2x4_ASAP7_75t_L g1602 ( 
.A(n_1537),
.B(n_1409),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1563),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1571),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1492),
.B(n_1451),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1515),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1493),
.B(n_1553),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1528),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1526),
.B(n_1527),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1532),
.B(n_1377),
.Y(n_1610)
);

BUFx3_ASAP7_75t_L g1611 ( 
.A(n_1516),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1528),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1489),
.A2(n_1409),
.B(n_1464),
.C(n_1453),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1538),
.Y(n_1614)
);

BUFx6f_ASAP7_75t_L g1615 ( 
.A(n_1516),
.Y(n_1615)
);

BUFx10_ASAP7_75t_L g1616 ( 
.A(n_1504),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1560),
.B(n_1429),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1544),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1523),
.B(n_1390),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1544),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1568),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1559),
.B(n_1524),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1502),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1568),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1517),
.B(n_1471),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1516),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1535),
.B(n_1354),
.Y(n_1627)
);

HAxp5_ASAP7_75t_L g1628 ( 
.A(n_1582),
.B(n_1478),
.CON(n_1628),
.SN(n_1628)
);

AOI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1578),
.A2(n_1600),
.B(n_1619),
.Y(n_1629)
);

AO21x1_ASAP7_75t_L g1630 ( 
.A1(n_1605),
.A2(n_1562),
.B(n_1506),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1605),
.A2(n_1536),
.B(n_1506),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1613),
.A2(n_1498),
.B(n_1496),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1614),
.A2(n_1471),
.B1(n_1437),
.B2(n_1440),
.Y(n_1633)
);

A2O1A1Ixp33_ASAP7_75t_L g1634 ( 
.A1(n_1583),
.A2(n_1557),
.B(n_1555),
.C(n_1494),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1501),
.B(n_1451),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1575),
.A2(n_1494),
.B(n_1543),
.Y(n_1636)
);

AO31x2_ASAP7_75t_L g1637 ( 
.A1(n_1575),
.A2(n_1510),
.A3(n_1572),
.B(n_1508),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1595),
.A2(n_1543),
.B(n_1542),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1583),
.A2(n_1550),
.B(n_1510),
.C(n_1490),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1609),
.B(n_1607),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1592),
.B(n_1622),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1587),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1609),
.B(n_1397),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1588),
.B(n_1421),
.Y(n_1644)
);

AOI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1595),
.A2(n_1547),
.B(n_1541),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1605),
.A2(n_1501),
.B(n_1522),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1607),
.B(n_1397),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1588),
.A2(n_1539),
.B(n_1522),
.Y(n_1648)
);

INVx3_ASAP7_75t_L g1649 ( 
.A(n_1580),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1580),
.A2(n_1546),
.B(n_1539),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1580),
.A2(n_1546),
.B(n_1548),
.Y(n_1651)
);

OAI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1610),
.A2(n_1519),
.B(n_1518),
.Y(n_1652)
);

A2O1A1Ixp33_ASAP7_75t_L g1653 ( 
.A1(n_1610),
.A2(n_1497),
.B(n_1513),
.C(n_1505),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_SL g1654 ( 
.A(n_1588),
.B(n_1394),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1617),
.A2(n_1405),
.B1(n_1511),
.B2(n_1425),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1587),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1584),
.B(n_1512),
.Y(n_1657)
);

OAI21x1_ASAP7_75t_L g1658 ( 
.A1(n_1580),
.A2(n_1567),
.B(n_1548),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1616),
.B(n_1622),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1585),
.A2(n_1520),
.B(n_1622),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1597),
.A2(n_1567),
.B(n_1473),
.Y(n_1661)
);

OAI21x1_ASAP7_75t_L g1662 ( 
.A1(n_1597),
.A2(n_1473),
.B(n_1460),
.Y(n_1662)
);

BUFx3_ASAP7_75t_L g1663 ( 
.A(n_1594),
.Y(n_1663)
);

BUFx2_ASAP7_75t_L g1664 ( 
.A(n_1604),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1622),
.A2(n_1565),
.B(n_1234),
.Y(n_1665)
);

INVxp67_ASAP7_75t_L g1666 ( 
.A(n_1584),
.Y(n_1666)
);

BUFx3_ASAP7_75t_L g1667 ( 
.A(n_1594),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1625),
.B(n_1439),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1576),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1597),
.A2(n_1479),
.B(n_1460),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1593),
.A2(n_1549),
.B(n_1514),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1588),
.A2(n_1448),
.B(n_1225),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1597),
.A2(n_1479),
.B(n_1278),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1577),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1593),
.B(n_1599),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1623),
.A2(n_1280),
.B(n_1277),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1593),
.B(n_1439),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1642),
.Y(n_1678)
);

AO31x2_ASAP7_75t_L g1679 ( 
.A1(n_1630),
.A2(n_1589),
.A3(n_1612),
.B(n_1576),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1599),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1643),
.B(n_1602),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_L g1682 ( 
.A1(n_1647),
.A2(n_1599),
.B1(n_1616),
.B2(n_1486),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1663),
.Y(n_1683)
);

AND2x4_ASAP7_75t_L g1684 ( 
.A(n_1641),
.B(n_1588),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1660),
.B(n_1616),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1652),
.B(n_1616),
.Y(n_1687)
);

CKINVDCx20_ASAP7_75t_R g1688 ( 
.A(n_1674),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1663),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1641),
.B(n_1588),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1673),
.A2(n_1623),
.B(n_1589),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1656),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1667),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1669),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1677),
.B(n_1592),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1647),
.B(n_1602),
.Y(n_1696)
);

AO21x2_ASAP7_75t_L g1697 ( 
.A1(n_1632),
.A2(n_1442),
.B(n_1445),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1664),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1673),
.Y(n_1700)
);

O2A1O1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1655),
.A2(n_1446),
.B(n_510),
.C(n_530),
.Y(n_1701)
);

INVxp67_ASAP7_75t_L g1702 ( 
.A(n_1668),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1662),
.Y(n_1703)
);

BUFx3_ASAP7_75t_L g1704 ( 
.A(n_1667),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1675),
.B(n_1576),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1662),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1670),
.Y(n_1707)
);

CKINVDCx5p33_ASAP7_75t_R g1708 ( 
.A(n_1633),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1644),
.A2(n_1484),
.B1(n_1420),
.B2(n_1433),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1641),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1666),
.B(n_1592),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1671),
.B(n_1589),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1653),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1644),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1653),
.Y(n_1715)
);

INVx4_ASAP7_75t_L g1716 ( 
.A(n_1644),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1645),
.B(n_1592),
.Y(n_1717)
);

O2A1O1Ixp33_ASAP7_75t_L g1718 ( 
.A1(n_1628),
.A2(n_510),
.B(n_530),
.C(n_514),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1670),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1649),
.Y(n_1720)
);

BUFx12f_ASAP7_75t_L g1721 ( 
.A(n_1628),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1634),
.A2(n_1402),
.B1(n_1602),
.B2(n_1020),
.Y(n_1722)
);

BUFx3_ASAP7_75t_L g1723 ( 
.A(n_1649),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1724)
);

NOR2xp67_ASAP7_75t_L g1725 ( 
.A(n_1649),
.B(n_1435),
.Y(n_1725)
);

INVx2_ASAP7_75t_SL g1726 ( 
.A(n_1659),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1646),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1676),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1659),
.Y(n_1729)
);

INVx6_ASAP7_75t_L g1730 ( 
.A(n_1654),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1637),
.B(n_1612),
.Y(n_1731)
);

INVx3_ASAP7_75t_SL g1732 ( 
.A(n_1639),
.Y(n_1732)
);

INVxp67_ASAP7_75t_L g1733 ( 
.A(n_1665),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1638),
.B(n_1590),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1648),
.B(n_1623),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1646),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1635),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1650),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1639),
.B(n_1590),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1636),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1676),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1635),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1634),
.B(n_1591),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1658),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1661),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1658),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1672),
.A2(n_1448),
.B(n_1540),
.Y(n_1747)
);

INVx4_ASAP7_75t_L g1748 ( 
.A(n_1650),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1637),
.B(n_1591),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1631),
.A2(n_1623),
.B(n_1618),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1651),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1651),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1637),
.B(n_1612),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1631),
.A2(n_1448),
.B(n_1540),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1661),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1637),
.A2(n_1448),
.B(n_1551),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1660),
.B(n_1422),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1664),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1642),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1642),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1675),
.B(n_1618),
.Y(n_1762)
);

AND2x4_ASAP7_75t_L g1763 ( 
.A(n_1641),
.B(n_1606),
.Y(n_1763)
);

INVx4_ASAP7_75t_L g1764 ( 
.A(n_1689),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1678),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1704),
.Y(n_1766)
);

INVx3_ASAP7_75t_L g1767 ( 
.A(n_1704),
.Y(n_1767)
);

BUFx2_ASAP7_75t_L g1768 ( 
.A(n_1683),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1685),
.B(n_1604),
.Y(n_1769)
);

OAI21x1_ASAP7_75t_L g1770 ( 
.A1(n_1754),
.A2(n_1387),
.B(n_1364),
.Y(n_1770)
);

OAI21x1_ASAP7_75t_L g1771 ( 
.A1(n_1756),
.A2(n_1387),
.B(n_1364),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1710),
.B(n_1601),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1691),
.A2(n_1620),
.B(n_1618),
.Y(n_1773)
);

CKINVDCx6p67_ASAP7_75t_R g1774 ( 
.A(n_1688),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1691),
.A2(n_1620),
.B(n_1495),
.Y(n_1775)
);

OAI21x1_ASAP7_75t_L g1776 ( 
.A1(n_1736),
.A2(n_1620),
.B(n_1495),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_SL g1777 ( 
.A(n_1688),
.B(n_1579),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1708),
.A2(n_1478),
.B1(n_682),
.B2(n_717),
.Y(n_1778)
);

OAI21x1_ASAP7_75t_L g1779 ( 
.A1(n_1736),
.A2(n_1621),
.B(n_1608),
.Y(n_1779)
);

INVxp67_ASAP7_75t_SL g1780 ( 
.A(n_1744),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1700),
.A2(n_841),
.B(n_840),
.Y(n_1781)
);

OR2x2_ASAP7_75t_SL g1782 ( 
.A(n_1724),
.B(n_1425),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1692),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1689),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1689),
.Y(n_1785)
);

OAI21x1_ASAP7_75t_L g1786 ( 
.A1(n_1747),
.A2(n_1551),
.B(n_1608),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1708),
.A2(n_1478),
.B1(n_682),
.B2(n_717),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1760),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1761),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1750),
.A2(n_1624),
.B(n_1621),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1750),
.A2(n_1624),
.B(n_1529),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1702),
.B(n_1601),
.Y(n_1792)
);

OAI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1736),
.A2(n_1706),
.B(n_1703),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1729),
.Y(n_1794)
);

NAND2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1716),
.B(n_1713),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1689),
.Y(n_1796)
);

OAI21x1_ASAP7_75t_L g1797 ( 
.A1(n_1700),
.A2(n_1454),
.B(n_1525),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1698),
.Y(n_1798)
);

INVx1_ASAP7_75t_SL g1799 ( 
.A(n_1693),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1680),
.B(n_1601),
.Y(n_1800)
);

OA21x2_ASAP7_75t_L g1801 ( 
.A1(n_1703),
.A2(n_844),
.B(n_842),
.Y(n_1801)
);

OAI21x1_ASAP7_75t_L g1802 ( 
.A1(n_1706),
.A2(n_1454),
.B(n_1533),
.Y(n_1802)
);

AND3x2_ASAP7_75t_L g1803 ( 
.A(n_1733),
.B(n_1566),
.C(n_643),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_SL g1804 ( 
.A1(n_1740),
.A2(n_1260),
.B1(n_1020),
.B2(n_1023),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1732),
.A2(n_655),
.B1(n_540),
.B2(n_559),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1695),
.B(n_1603),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1694),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1726),
.Y(n_1808)
);

OA21x2_ASAP7_75t_L g1809 ( 
.A1(n_1707),
.A2(n_847),
.B(n_845),
.Y(n_1809)
);

INVx2_ASAP7_75t_SL g1810 ( 
.A(n_1693),
.Y(n_1810)
);

AOI21x1_ASAP7_75t_L g1811 ( 
.A1(n_1734),
.A2(n_1259),
.B(n_1305),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1717),
.B(n_1458),
.Y(n_1812)
);

BUFx6f_ASAP7_75t_L g1813 ( 
.A(n_1693),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1705),
.B(n_1500),
.Y(n_1814)
);

BUFx2_ASAP7_75t_L g1815 ( 
.A(n_1693),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1705),
.B(n_1596),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1762),
.B(n_1627),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1726),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1707),
.A2(n_1554),
.B(n_1545),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1749),
.Y(n_1820)
);

AOI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1701),
.A2(n_586),
.B1(n_587),
.B2(n_585),
.C(n_574),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1762),
.B(n_1627),
.Y(n_1822)
);

AO32x2_ASAP7_75t_L g1823 ( 
.A1(n_1698),
.A2(n_1574),
.A3(n_1626),
.B1(n_1561),
.B2(n_1535),
.Y(n_1823)
);

CKINVDCx5p33_ASAP7_75t_R g1824 ( 
.A(n_1758),
.Y(n_1824)
);

OAI21x1_ASAP7_75t_L g1825 ( 
.A1(n_1719),
.A2(n_1570),
.B(n_1408),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1758),
.Y(n_1826)
);

AOI21xp5_ASAP7_75t_L g1827 ( 
.A1(n_1697),
.A2(n_1558),
.B(n_1380),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1716),
.B(n_1611),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1699),
.Y(n_1829)
);

OAI21xp5_ASAP7_75t_L g1830 ( 
.A1(n_1722),
.A2(n_1586),
.B(n_1353),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1711),
.B(n_1596),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1719),
.A2(n_1408),
.B(n_1419),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1732),
.A2(n_655),
.B1(n_540),
.B2(n_559),
.Y(n_1833)
);

AO32x2_ASAP7_75t_L g1834 ( 
.A1(n_1716),
.A2(n_1626),
.A3(n_1561),
.B1(n_1535),
.B2(n_1374),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1699),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_SL g1836 ( 
.A1(n_1740),
.A2(n_571),
.B1(n_576),
.B2(n_514),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1728),
.A2(n_1428),
.B(n_1424),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1679),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1749),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1696),
.B(n_1627),
.Y(n_1840)
);

OA21x2_ASAP7_75t_L g1841 ( 
.A1(n_1751),
.A2(n_774),
.B(n_772),
.Y(n_1841)
);

INVx4_ASAP7_75t_L g1842 ( 
.A(n_1730),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1679),
.Y(n_1843)
);

OAI21x1_ASAP7_75t_L g1844 ( 
.A1(n_1727),
.A2(n_1742),
.B(n_1737),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1731),
.Y(n_1845)
);

OAI21x1_ASAP7_75t_L g1846 ( 
.A1(n_1745),
.A2(n_1360),
.B(n_1357),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_SL g1847 ( 
.A1(n_1721),
.A2(n_1260),
.B1(n_1382),
.B2(n_1001),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1679),
.Y(n_1848)
);

OAI21x1_ASAP7_75t_L g1849 ( 
.A1(n_1745),
.A2(n_1367),
.B(n_1362),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1731),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_L g1851 ( 
.A1(n_1752),
.A2(n_1372),
.B(n_1368),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1714),
.B(n_1611),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1753),
.Y(n_1853)
);

AOI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1696),
.A2(n_1353),
.B1(n_1281),
.B2(n_1290),
.Y(n_1854)
);

OAI21x1_ASAP7_75t_L g1855 ( 
.A1(n_1728),
.A2(n_1373),
.B(n_1430),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1697),
.A2(n_1380),
.B(n_1374),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1753),
.Y(n_1857)
);

AO21x2_ASAP7_75t_L g1858 ( 
.A1(n_1746),
.A2(n_1259),
.B(n_1305),
.Y(n_1858)
);

AO31x2_ASAP7_75t_L g1859 ( 
.A1(n_1748),
.A2(n_1738),
.A3(n_1741),
.B(n_1755),
.Y(n_1859)
);

AOI31xp67_ASAP7_75t_L g1860 ( 
.A1(n_1741),
.A2(n_1418),
.A3(n_1426),
.B(n_1416),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1712),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1712),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1720),
.Y(n_1863)
);

OAI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1709),
.A2(n_576),
.B1(n_579),
.B2(n_571),
.Y(n_1864)
);

OAI21xp5_ASAP7_75t_L g1865 ( 
.A1(n_1681),
.A2(n_1627),
.B(n_593),
.Y(n_1865)
);

INVx4_ASAP7_75t_L g1866 ( 
.A(n_1730),
.Y(n_1866)
);

CKINVDCx14_ASAP7_75t_R g1867 ( 
.A(n_1681),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1682),
.A2(n_1594),
.B1(n_1581),
.B2(n_1435),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_SL g1869 ( 
.A(n_1687),
.B(n_1422),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1718),
.A2(n_1686),
.B(n_1757),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1679),
.Y(n_1871)
);

INVx5_ASAP7_75t_L g1872 ( 
.A(n_1748),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1763),
.Y(n_1873)
);

OAI21x1_ASAP7_75t_L g1874 ( 
.A1(n_1739),
.A2(n_1434),
.B(n_1431),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1735),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1721),
.A2(n_1281),
.B1(n_1290),
.B2(n_1268),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1697),
.A2(n_593),
.B1(n_602),
.B2(n_579),
.Y(n_1877)
);

OA21x2_ASAP7_75t_L g1878 ( 
.A1(n_1715),
.A2(n_774),
.B(n_772),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1735),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1714),
.Y(n_1880)
);

INVx3_ASAP7_75t_L g1881 ( 
.A(n_1723),
.Y(n_1881)
);

AOI21x1_ASAP7_75t_L g1882 ( 
.A1(n_1725),
.A2(n_777),
.B(n_775),
.Y(n_1882)
);

AO21x2_ASAP7_75t_L g1883 ( 
.A1(n_1757),
.A2(n_606),
.B(n_602),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1759),
.B(n_591),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1735),
.Y(n_1885)
);

AO21x2_ASAP7_75t_L g1886 ( 
.A1(n_1743),
.A2(n_612),
.B(n_606),
.Y(n_1886)
);

OAI21x1_ASAP7_75t_L g1887 ( 
.A1(n_1748),
.A2(n_1441),
.B(n_1438),
.Y(n_1887)
);

BUFx8_ASAP7_75t_SL g1888 ( 
.A(n_1763),
.Y(n_1888)
);

OAI21x1_ASAP7_75t_L g1889 ( 
.A1(n_1730),
.A2(n_1465),
.B(n_1463),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1684),
.B(n_1611),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1763),
.B(n_1723),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1684),
.B(n_596),
.Y(n_1892)
);

NAND2x1p5_ASAP7_75t_L g1893 ( 
.A(n_1684),
.B(n_1615),
.Y(n_1893)
);

AOI221xp5_ASAP7_75t_L g1894 ( 
.A1(n_1690),
.A2(n_609),
.B1(n_610),
.B2(n_605),
.C(n_600),
.Y(n_1894)
);

BUFx2_ASAP7_75t_L g1895 ( 
.A(n_1690),
.Y(n_1895)
);

AND2x4_ASAP7_75t_L g1896 ( 
.A(n_1690),
.B(n_1626),
.Y(n_1896)
);

A2O1A1Ixp33_ASAP7_75t_L g1897 ( 
.A1(n_1730),
.A2(n_643),
.B(n_648),
.C(n_612),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1678),
.Y(n_1898)
);

BUFx2_ASAP7_75t_SL g1899 ( 
.A(n_1688),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1704),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1678),
.Y(n_1901)
);

OAI21x1_ASAP7_75t_L g1902 ( 
.A1(n_1754),
.A2(n_1475),
.B(n_1469),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1708),
.A2(n_649),
.B1(n_650),
.B2(n_648),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1678),
.Y(n_1904)
);

INVxp67_ASAP7_75t_SL g1905 ( 
.A(n_1744),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1710),
.B(n_1466),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1708),
.A2(n_1268),
.B1(n_1342),
.B2(n_1318),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1710),
.B(n_1615),
.Y(n_1908)
);

CKINVDCx12_ASAP7_75t_R g1909 ( 
.A(n_1688),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1744),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1678),
.Y(n_1911)
);

OAI22xp5_ASAP7_75t_L g1912 ( 
.A1(n_1708),
.A2(n_1318),
.B1(n_1302),
.B2(n_1468),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1678),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1678),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1704),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1861),
.B(n_775),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1904),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1904),
.Y(n_1918)
);

AOI22xp33_ASAP7_75t_L g1919 ( 
.A1(n_1867),
.A2(n_495),
.B1(n_517),
.B2(n_503),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1765),
.Y(n_1920)
);

INVxp67_ASAP7_75t_L g1921 ( 
.A(n_1826),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1824),
.Y(n_1922)
);

OAI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1793),
.A2(n_1481),
.B(n_1476),
.Y(n_1923)
);

NAND4xp25_ASAP7_75t_L g1924 ( 
.A(n_1903),
.B(n_649),
.C(n_651),
.D(n_650),
.Y(n_1924)
);

AND2x4_ASAP7_75t_L g1925 ( 
.A(n_1875),
.B(n_1615),
.Y(n_1925)
);

INVx6_ASAP7_75t_L g1926 ( 
.A(n_1813),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1867),
.A2(n_495),
.B1(n_517),
.B2(n_503),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1783),
.Y(n_1928)
);

OAI22xp5_ASAP7_75t_L g1929 ( 
.A1(n_1778),
.A2(n_652),
.B1(n_663),
.B2(n_651),
.Y(n_1929)
);

OAI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1854),
.A2(n_663),
.B1(n_667),
.B2(n_652),
.Y(n_1930)
);

INVxp67_ASAP7_75t_SL g1931 ( 
.A(n_1910),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_1774),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1788),
.Y(n_1933)
);

AOI22xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1865),
.A2(n_1001),
.B1(n_517),
.B2(n_626),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1789),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1898),
.Y(n_1936)
);

AND2x4_ASAP7_75t_L g1937 ( 
.A(n_1875),
.B(n_1615),
.Y(n_1937)
);

BUFx4f_ASAP7_75t_SL g1938 ( 
.A(n_1880),
.Y(n_1938)
);

AOI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1864),
.A2(n_580),
.B1(n_626),
.B2(n_667),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1864),
.A2(n_669),
.B1(n_685),
.B2(n_677),
.Y(n_1940)
);

NAND2xp33_ASAP7_75t_SL g1941 ( 
.A(n_1880),
.B(n_1598),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1901),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1911),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1895),
.B(n_669),
.Y(n_1944)
);

CKINVDCx12_ASAP7_75t_R g1945 ( 
.A(n_1906),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1862),
.B(n_677),
.Y(n_1946)
);

HB1xp67_ASAP7_75t_L g1947 ( 
.A(n_1798),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1913),
.Y(n_1948)
);

BUFx4f_ASAP7_75t_L g1949 ( 
.A(n_1813),
.Y(n_1949)
);

AOI22xp5_ASAP7_75t_L g1950 ( 
.A1(n_1778),
.A2(n_685),
.B1(n_693),
.B2(n_687),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1804),
.A2(n_693),
.B1(n_697),
.B2(n_687),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1787),
.A2(n_699),
.B1(n_701),
.B2(n_697),
.Y(n_1952)
);

BUFx3_ASAP7_75t_L g1953 ( 
.A(n_1824),
.Y(n_1953)
);

HB1xp67_ASAP7_75t_L g1954 ( 
.A(n_1798),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_SL g1955 ( 
.A(n_1836),
.B(n_1334),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1794),
.B(n_699),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1812),
.A2(n_580),
.B1(n_626),
.B2(n_701),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1768),
.B(n_722),
.Y(n_1958)
);

BUFx4f_ASAP7_75t_SL g1959 ( 
.A(n_1796),
.Y(n_1959)
);

AOI22xp33_ASAP7_75t_L g1960 ( 
.A1(n_1870),
.A2(n_580),
.B1(n_722),
.B2(n_705),
.Y(n_1960)
);

BUFx12f_ASAP7_75t_L g1961 ( 
.A(n_1782),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1914),
.Y(n_1962)
);

OAI22xp5_ASAP7_75t_L g1963 ( 
.A1(n_1787),
.A2(n_1480),
.B1(n_615),
.B2(n_616),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1769),
.B(n_777),
.Y(n_1964)
);

INVx3_ASAP7_75t_L g1965 ( 
.A(n_1813),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1879),
.B(n_1615),
.Y(n_1966)
);

BUFx2_ASAP7_75t_L g1967 ( 
.A(n_1888),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1873),
.B(n_778),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1808),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_SL g1970 ( 
.A1(n_1804),
.A2(n_617),
.B1(n_618),
.B2(n_613),
.Y(n_1970)
);

AOI222xp33_ASAP7_75t_L g1971 ( 
.A1(n_1903),
.A2(n_705),
.B1(n_714),
.B2(n_496),
.C1(n_622),
.C2(n_623),
.Y(n_1971)
);

AOI22xp33_ASAP7_75t_SL g1972 ( 
.A1(n_1830),
.A2(n_705),
.B1(n_714),
.B2(n_496),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_L g1973 ( 
.A1(n_1805),
.A2(n_620),
.B(n_631),
.C(n_619),
.Y(n_1973)
);

INVx1_ASAP7_75t_L g1974 ( 
.A(n_1807),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1805),
.A2(n_1480),
.B1(n_635),
.B2(n_636),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1887),
.A2(n_1436),
.B(n_1432),
.Y(n_1976)
);

OAI21x1_ASAP7_75t_L g1977 ( 
.A1(n_1887),
.A2(n_1462),
.B(n_1457),
.Y(n_1977)
);

OR2x6_ASAP7_75t_L g1978 ( 
.A(n_1795),
.B(n_1615),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_SL g1979 ( 
.A1(n_1886),
.A2(n_714),
.B1(n_496),
.B2(n_1334),
.Y(n_1979)
);

BUFx5_ASAP7_75t_L g1980 ( 
.A(n_1885),
.Y(n_1980)
);

AOI22xp33_ASAP7_75t_SL g1981 ( 
.A1(n_1886),
.A2(n_1334),
.B1(n_638),
.B2(n_641),
.Y(n_1981)
);

AOI22xp33_ASAP7_75t_L g1982 ( 
.A1(n_1877),
.A2(n_1295),
.B1(n_1274),
.B2(n_849),
.Y(n_1982)
);

INVx2_ASAP7_75t_SL g1983 ( 
.A(n_1813),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1877),
.A2(n_1295),
.B1(n_1274),
.B2(n_849),
.Y(n_1984)
);

AOI21x1_ASAP7_75t_L g1985 ( 
.A1(n_1892),
.A2(n_1869),
.B(n_1882),
.Y(n_1985)
);

AND2x2_ASAP7_75t_L g1986 ( 
.A(n_1900),
.B(n_778),
.Y(n_1986)
);

NAND2xp33_ASAP7_75t_R g1987 ( 
.A(n_1803),
.B(n_1198),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1796),
.Y(n_1988)
);

NAND2xp33_ASAP7_75t_SL g1989 ( 
.A(n_1833),
.B(n_632),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_SL g1990 ( 
.A(n_1777),
.B(n_1899),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1845),
.B(n_851),
.Y(n_1991)
);

BUFx8_ASAP7_75t_L g1992 ( 
.A(n_1915),
.Y(n_1992)
);

AOI221xp5_ASAP7_75t_L g1993 ( 
.A1(n_1833),
.A2(n_656),
.B1(n_657),
.B2(n_647),
.C(n_645),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1785),
.B(n_851),
.Y(n_1994)
);

BUFx3_ASAP7_75t_L g1995 ( 
.A(n_1815),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1827),
.A2(n_1417),
.B(n_1394),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1818),
.Y(n_1997)
);

BUFx6f_ASAP7_75t_L g1998 ( 
.A(n_1764),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1897),
.A2(n_854),
.B(n_852),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1814),
.B(n_1800),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1829),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1890),
.B(n_1817),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1829),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1835),
.Y(n_2004)
);

OAI22xp5_ASAP7_75t_L g2005 ( 
.A1(n_1847),
.A2(n_662),
.B1(n_664),
.B2(n_661),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1856),
.A2(n_1417),
.B(n_1394),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1784),
.Y(n_2007)
);

OAI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1831),
.A2(n_668),
.B1(n_670),
.B2(n_665),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1835),
.Y(n_2009)
);

O2A1O1Ixp33_ASAP7_75t_SL g2010 ( 
.A1(n_1897),
.A2(n_1509),
.B(n_1491),
.C(n_854),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1822),
.B(n_852),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1863),
.B(n_857),
.Y(n_2012)
);

OAI221xp5_ASAP7_75t_L g2013 ( 
.A1(n_1894),
.A2(n_684),
.B1(n_688),
.B2(n_675),
.C(n_672),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1847),
.A2(n_1912),
.B1(n_1868),
.B2(n_1907),
.Y(n_2014)
);

AOI22xp5_ASAP7_75t_L g2015 ( 
.A1(n_1803),
.A2(n_1876),
.B1(n_1806),
.B2(n_1816),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1910),
.Y(n_2016)
);

AO21x2_ASAP7_75t_L g2017 ( 
.A1(n_1838),
.A2(n_859),
.B(n_857),
.Y(n_2017)
);

INVx6_ASAP7_75t_L g2018 ( 
.A(n_1764),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1891),
.B(n_859),
.Y(n_2019)
);

OR2x6_ASAP7_75t_L g2020 ( 
.A(n_1795),
.B(n_1516),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1850),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1869),
.B(n_860),
.Y(n_2022)
);

AOI21xp33_ASAP7_75t_L g2023 ( 
.A1(n_1884),
.A2(n_862),
.B(n_860),
.Y(n_2023)
);

AOI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_1821),
.A2(n_694),
.B(n_696),
.C(n_691),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1890),
.B(n_862),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1792),
.A2(n_703),
.B1(n_704),
.B2(n_700),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1853),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1857),
.Y(n_2028)
);

AND2x4_ASAP7_75t_L g2029 ( 
.A(n_1863),
.B(n_863),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1840),
.A2(n_1883),
.B1(n_1909),
.B2(n_1772),
.Y(n_2030)
);

INVx2_ASAP7_75t_L g2031 ( 
.A(n_1766),
.Y(n_2031)
);

NAND2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1842),
.B(n_1866),
.Y(n_2032)
);

OAI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1842),
.A2(n_718),
.B1(n_720),
.B2(n_709),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1766),
.B(n_863),
.Y(n_2034)
);

OAI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1889),
.A2(n_983),
.B(n_724),
.Y(n_2035)
);

AOI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1883),
.A2(n_725),
.B1(n_726),
.B2(n_723),
.Y(n_2036)
);

BUFx6f_ASAP7_75t_L g2037 ( 
.A(n_1784),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1820),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1839),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1780),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1890),
.B(n_3),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1896),
.B(n_3),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1780),
.Y(n_2043)
);

NAND2xp33_ASAP7_75t_L g2044 ( 
.A(n_1810),
.B(n_1422),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1889),
.A2(n_1417),
.B(n_1269),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1905),
.Y(n_2046)
);

AOI22xp33_ASAP7_75t_L g2047 ( 
.A1(n_1896),
.A2(n_1295),
.B1(n_1274),
.B2(n_1456),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1896),
.A2(n_1295),
.B1(n_1274),
.B2(n_1456),
.Y(n_2048)
);

OAI22xp5_ASAP7_75t_L g2049 ( 
.A1(n_1866),
.A2(n_1369),
.B1(n_1561),
.B2(n_456),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_1905),
.A2(n_464),
.B1(n_466),
.B2(n_457),
.C(n_454),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_1893),
.A2(n_1369),
.B1(n_473),
.B2(n_474),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1852),
.A2(n_907),
.B1(n_903),
.B2(n_477),
.Y(n_2052)
);

AND2x2_ASAP7_75t_L g2053 ( 
.A(n_1767),
.B(n_4),
.Y(n_2053)
);

OAI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_1893),
.A2(n_479),
.B1(n_485),
.B2(n_478),
.C(n_471),
.Y(n_2054)
);

OAI21x1_ASAP7_75t_L g2055 ( 
.A1(n_1844),
.A2(n_1474),
.B(n_1472),
.Y(n_2055)
);

NOR3xp33_ASAP7_75t_SL g2056 ( 
.A(n_1823),
.B(n_493),
.C(n_491),
.Y(n_2056)
);

INVx2_ASAP7_75t_SL g2057 ( 
.A(n_1767),
.Y(n_2057)
);

AOI22xp33_ASAP7_75t_L g2058 ( 
.A1(n_1852),
.A2(n_1828),
.B1(n_1888),
.B2(n_1881),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1799),
.B(n_1255),
.Y(n_2059)
);

BUFx3_ASAP7_75t_L g2060 ( 
.A(n_1852),
.Y(n_2060)
);

OAI211xp5_ASAP7_75t_SL g2061 ( 
.A1(n_1881),
.A2(n_868),
.B(n_870),
.C(n_866),
.Y(n_2061)
);

AND2x2_ASAP7_75t_SL g2062 ( 
.A(n_1828),
.B(n_903),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1828),
.A2(n_500),
.B1(n_505),
.B2(n_494),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1908),
.B(n_5),
.Y(n_2064)
);

BUFx2_ASAP7_75t_SL g2065 ( 
.A(n_1872),
.Y(n_2065)
);

INVx3_ASAP7_75t_L g2066 ( 
.A(n_1872),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_1779),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1859),
.Y(n_2068)
);

OAI22xp5_ASAP7_75t_L g2069 ( 
.A1(n_1872),
.A2(n_512),
.B1(n_513),
.B2(n_511),
.Y(n_2069)
);

INVxp33_ASAP7_75t_L g2070 ( 
.A(n_1819),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1779),
.Y(n_2071)
);

AOI21xp5_ASAP7_75t_L g2072 ( 
.A1(n_1874),
.A2(n_1786),
.B(n_1878),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1859),
.Y(n_2073)
);

AOI221xp5_ASAP7_75t_L g2074 ( 
.A1(n_1838),
.A2(n_521),
.B1(n_522),
.B2(n_519),
.C(n_515),
.Y(n_2074)
);

AOI22xp33_ASAP7_75t_L g2075 ( 
.A1(n_1858),
.A2(n_907),
.B1(n_535),
.B2(n_536),
.Y(n_2075)
);

NAND3xp33_ASAP7_75t_SL g2076 ( 
.A(n_1843),
.B(n_538),
.C(n_532),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2040),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2043),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2046),
.Y(n_2079)
);

OAI33xp33_ASAP7_75t_L g2080 ( 
.A1(n_1970),
.A2(n_1848),
.A3(n_1871),
.B1(n_1843),
.B2(n_546),
.B3(n_544),
.Y(n_2080)
);

HB1xp67_ASAP7_75t_L g2081 ( 
.A(n_1947),
.Y(n_2081)
);

OAI21x1_ASAP7_75t_L g2082 ( 
.A1(n_2072),
.A2(n_1871),
.B(n_1848),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_1954),
.B(n_1859),
.Y(n_2083)
);

INVx2_ASAP7_75t_L g2084 ( 
.A(n_2073),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2038),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2068),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_2067),
.A2(n_2071),
.B(n_1996),
.Y(n_2087)
);

AOI22xp33_ASAP7_75t_L g2088 ( 
.A1(n_1934),
.A2(n_1858),
.B1(n_1874),
.B2(n_1770),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1917),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_2016),
.B(n_1859),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2002),
.B(n_1872),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1918),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1931),
.Y(n_2093)
);

BUFx2_ASAP7_75t_L g2094 ( 
.A(n_1992),
.Y(n_2094)
);

INVx3_ASAP7_75t_L g2095 ( 
.A(n_2066),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_1992),
.Y(n_2096)
);

BUFx6f_ASAP7_75t_L g2097 ( 
.A(n_1998),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_2066),
.A2(n_1802),
.B(n_1797),
.Y(n_2098)
);

AOI21x1_ASAP7_75t_L g2099 ( 
.A1(n_2034),
.A2(n_1841),
.B(n_1809),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2001),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2039),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2004),
.Y(n_2102)
);

OA21x2_ASAP7_75t_L g2103 ( 
.A1(n_2056),
.A2(n_1802),
.B(n_1797),
.Y(n_2103)
);

INVxp67_ASAP7_75t_L g2104 ( 
.A(n_1986),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1980),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_2009),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_2021),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_2003),
.Y(n_2108)
);

INVxp67_ASAP7_75t_SL g2109 ( 
.A(n_2019),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2027),
.B(n_1841),
.Y(n_2110)
);

INVx2_ASAP7_75t_SL g2111 ( 
.A(n_2018),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_2006),
.A2(n_1825),
.B(n_1832),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1969),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1997),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1920),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_2018),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1928),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1935),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1936),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1942),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_2028),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1943),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1948),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1933),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1962),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_1995),
.B(n_1823),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1980),
.Y(n_2127)
);

OAI21x1_ASAP7_75t_L g2128 ( 
.A1(n_1976),
.A2(n_1832),
.B(n_1809),
.Y(n_2128)
);

AOI21x1_ASAP7_75t_L g2129 ( 
.A1(n_1985),
.A2(n_1841),
.B(n_1809),
.Y(n_2129)
);

AO21x2_ASAP7_75t_L g2130 ( 
.A1(n_2017),
.A2(n_1776),
.B(n_1775),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1980),
.Y(n_2131)
);

NOR2x1_ASAP7_75t_L g2132 ( 
.A(n_2065),
.B(n_1781),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_1938),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1980),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1974),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_1980),
.Y(n_2136)
);

NAND2x1p5_ASAP7_75t_L g2137 ( 
.A(n_1949),
.B(n_1781),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_2060),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1916),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1991),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1967),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_2031),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1994),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_1965),
.Y(n_2144)
);

HB1xp67_ASAP7_75t_L g2145 ( 
.A(n_2057),
.Y(n_2145)
);

INVx6_ASAP7_75t_L g2146 ( 
.A(n_1961),
.Y(n_2146)
);

INVx2_ASAP7_75t_L g2147 ( 
.A(n_1965),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1968),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_2025),
.Y(n_2149)
);

AO21x2_ASAP7_75t_L g2150 ( 
.A1(n_2017),
.A2(n_1776),
.B(n_1775),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2037),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2037),
.Y(n_2152)
);

INVx3_ASAP7_75t_L g2153 ( 
.A(n_2037),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_2007),
.Y(n_2154)
);

INVx3_ASAP7_75t_L g2155 ( 
.A(n_1998),
.Y(n_2155)
);

INVx2_ASAP7_75t_L g2156 ( 
.A(n_2012),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_1978),
.B(n_1790),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1921),
.B(n_1823),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1946),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2070),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_2000),
.Y(n_2161)
);

OAI21x1_ASAP7_75t_L g2162 ( 
.A1(n_1977),
.A2(n_1801),
.B(n_1781),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2012),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_1988),
.B(n_1823),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1956),
.Y(n_2165)
);

BUFx6f_ASAP7_75t_L g2166 ( 
.A(n_1998),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1925),
.Y(n_2167)
);

AO21x2_ASAP7_75t_L g2168 ( 
.A1(n_2022),
.A2(n_1837),
.B(n_1773),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1983),
.B(n_1801),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2029),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_1926),
.Y(n_2171)
);

AOI22xp33_ASAP7_75t_L g2172 ( 
.A1(n_1972),
.A2(n_1770),
.B1(n_1771),
.B2(n_1878),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1926),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2029),
.Y(n_2174)
);

BUFx3_ASAP7_75t_L g2175 ( 
.A(n_2032),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_1953),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1925),
.Y(n_2177)
);

BUFx3_ASAP7_75t_L g2178 ( 
.A(n_1932),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1937),
.Y(n_2179)
);

BUFx3_ASAP7_75t_L g2180 ( 
.A(n_1944),
.Y(n_2180)
);

OR2x6_ASAP7_75t_L g2181 ( 
.A(n_1978),
.B(n_1771),
.Y(n_2181)
);

INVx2_ASAP7_75t_SL g2182 ( 
.A(n_1922),
.Y(n_2182)
);

AND2x2_ASAP7_75t_L g2183 ( 
.A(n_1937),
.B(n_1801),
.Y(n_2183)
);

BUFx2_ASAP7_75t_SL g2184 ( 
.A(n_1958),
.Y(n_2184)
);

AOI21x1_ASAP7_75t_L g2185 ( 
.A1(n_1964),
.A2(n_1878),
.B(n_1811),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2058),
.B(n_1773),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2030),
.B(n_1834),
.Y(n_2187)
);

BUFx6f_ASAP7_75t_L g2188 ( 
.A(n_2020),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1966),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2030),
.B(n_1834),
.Y(n_2190)
);

BUFx4f_ASAP7_75t_L g2191 ( 
.A(n_2062),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_1966),
.B(n_1834),
.Y(n_2192)
);

NOR2xp33_ASAP7_75t_L g2193 ( 
.A(n_1990),
.B(n_6),
.Y(n_2193)
);

INVx2_ASAP7_75t_L g2194 ( 
.A(n_1978),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2011),
.Y(n_2195)
);

OAI21x1_ASAP7_75t_L g2196 ( 
.A1(n_1923),
.A2(n_1837),
.B(n_1791),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_2020),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2020),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2041),
.B(n_1834),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2055),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2064),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2042),
.B(n_1902),
.Y(n_2202)
);

OAI21x1_ASAP7_75t_SL g2203 ( 
.A1(n_2014),
.A2(n_1851),
.B(n_1849),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2053),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1945),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1949),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1959),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2044),
.Y(n_2208)
);

AND2x4_ASAP7_75t_L g2209 ( 
.A(n_2015),
.B(n_1902),
.Y(n_2209)
);

OR2x6_ASAP7_75t_L g2210 ( 
.A(n_2045),
.B(n_1855),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2061),
.Y(n_2211)
);

OR2x6_ASAP7_75t_L g2212 ( 
.A(n_2035),
.B(n_1846),
.Y(n_2212)
);

OR2x2_ASAP7_75t_L g2213 ( 
.A(n_2015),
.B(n_6),
.Y(n_2213)
);

BUFx3_ASAP7_75t_L g2214 ( 
.A(n_2059),
.Y(n_2214)
);

OR2x6_ASAP7_75t_L g2215 ( 
.A(n_1955),
.B(n_1860),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1930),
.B(n_7),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_2063),
.B(n_7),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_1919),
.B(n_8),
.Y(n_2218)
);

BUFx3_ASAP7_75t_L g2219 ( 
.A(n_2063),
.Y(n_2219)
);

OA21x2_ASAP7_75t_L g2220 ( 
.A1(n_2075),
.A2(n_868),
.B(n_866),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1999),
.Y(n_2221)
);

BUFx3_ASAP7_75t_L g2222 ( 
.A(n_1951),
.Y(n_2222)
);

INVx8_ASAP7_75t_L g2223 ( 
.A(n_1941),
.Y(n_2223)
);

AND2x2_ASAP7_75t_SL g2224 ( 
.A(n_1960),
.B(n_8),
.Y(n_2224)
);

AO21x2_ASAP7_75t_L g2225 ( 
.A1(n_2076),
.A2(n_880),
.B(n_870),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_1927),
.B(n_9),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_1924),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2036),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2036),
.Y(n_2229)
);

AND2x2_ASAP7_75t_L g2230 ( 
.A(n_1979),
.B(n_9),
.Y(n_2230)
);

AND2x2_ASAP7_75t_L g2231 ( 
.A(n_2026),
.B(n_10),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1940),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1940),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2051),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_2069),
.Y(n_2235)
);

OAI21x1_ASAP7_75t_L g2236 ( 
.A1(n_2049),
.A2(n_1447),
.B(n_882),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1951),
.Y(n_2237)
);

INVxp67_ASAP7_75t_L g2238 ( 
.A(n_1987),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2054),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2010),
.Y(n_2240)
);

INVx1_ASAP7_75t_SL g2241 ( 
.A(n_2184),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_2132),
.A2(n_2033),
.B(n_1957),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2125),
.Y(n_2243)
);

AND2x4_ASAP7_75t_SL g2244 ( 
.A(n_2207),
.B(n_1950),
.Y(n_2244)
);

AOI22xp5_ASAP7_75t_L g2245 ( 
.A1(n_2219),
.A2(n_1970),
.B1(n_1950),
.B2(n_1981),
.Y(n_2245)
);

INVxp67_ASAP7_75t_L g2246 ( 
.A(n_2184),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2125),
.Y(n_2247)
);

AND2x2_ASAP7_75t_L g2248 ( 
.A(n_2091),
.B(n_2047),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2222),
.A2(n_1939),
.B1(n_2024),
.B2(n_1952),
.Y(n_2249)
);

OAI221xp5_ASAP7_75t_L g2250 ( 
.A1(n_2219),
.A2(n_1971),
.B1(n_2024),
.B2(n_1989),
.C(n_2005),
.Y(n_2250)
);

OR2x2_ASAP7_75t_L g2251 ( 
.A(n_2161),
.B(n_2023),
.Y(n_2251)
);

AOI222xp33_ASAP7_75t_L g2252 ( 
.A1(n_2224),
.A2(n_1929),
.B1(n_1993),
.B2(n_2013),
.C1(n_1973),
.C2(n_2008),
.Y(n_2252)
);

AOI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2219),
.A2(n_2074),
.B1(n_2050),
.B2(n_2048),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_SL g2254 ( 
.A1(n_2229),
.A2(n_1963),
.B1(n_1975),
.B2(n_545),
.Y(n_2254)
);

OR2x2_ASAP7_75t_L g2255 ( 
.A(n_2081),
.B(n_2052),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2091),
.B(n_11),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2115),
.Y(n_2257)
);

NOR2x1p5_ASAP7_75t_L g2258 ( 
.A(n_2096),
.B(n_542),
.Y(n_2258)
);

AOI22xp33_ASAP7_75t_L g2259 ( 
.A1(n_2229),
.A2(n_2228),
.B1(n_2239),
.B2(n_2080),
.Y(n_2259)
);

INVxp67_ASAP7_75t_L g2260 ( 
.A(n_2143),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2144),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_L g2262 ( 
.A1(n_2222),
.A2(n_1984),
.B1(n_1982),
.B2(n_550),
.Y(n_2262)
);

OAI22xp5_ASAP7_75t_L g2263 ( 
.A1(n_2228),
.A2(n_552),
.B1(n_554),
.B2(n_548),
.Y(n_2263)
);

O2A1O1Ixp33_ASAP7_75t_L g2264 ( 
.A1(n_2213),
.A2(n_14),
.B(n_12),
.C(n_13),
.Y(n_2264)
);

AOI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2094),
.A2(n_882),
.B(n_880),
.Y(n_2265)
);

OA21x2_ASAP7_75t_L g2266 ( 
.A1(n_2160),
.A2(n_557),
.B(n_556),
.Y(n_2266)
);

AOI22xp33_ASAP7_75t_L g2267 ( 
.A1(n_2239),
.A2(n_2224),
.B1(n_2217),
.B2(n_2191),
.Y(n_2267)
);

AOI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2224),
.A2(n_1126),
.B1(n_1131),
.B2(n_1123),
.Y(n_2268)
);

AND2x4_ASAP7_75t_L g2269 ( 
.A(n_2175),
.B(n_12),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2132),
.A2(n_910),
.B(n_895),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_2115),
.Y(n_2271)
);

BUFx2_ASAP7_75t_L g2272 ( 
.A(n_2094),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2139),
.B(n_13),
.Y(n_2273)
);

OAI221xp5_ASAP7_75t_L g2274 ( 
.A1(n_2213),
.A2(n_564),
.B1(n_567),
.B2(n_563),
.C(n_561),
.Y(n_2274)
);

INVx3_ASAP7_75t_L g2275 ( 
.A(n_2097),
.Y(n_2275)
);

HB1xp67_ASAP7_75t_L g2276 ( 
.A(n_2093),
.Y(n_2276)
);

OAI221xp5_ASAP7_75t_SL g2277 ( 
.A1(n_2230),
.A2(n_2216),
.B1(n_2237),
.B2(n_2218),
.C(n_2226),
.Y(n_2277)
);

AOI22xp33_ASAP7_75t_L g2278 ( 
.A1(n_2217),
.A2(n_1141),
.B1(n_573),
.B2(n_577),
.Y(n_2278)
);

OAI33xp33_ASAP7_75t_L g2279 ( 
.A1(n_2159),
.A2(n_594),
.A3(n_578),
.B1(n_601),
.B2(n_582),
.B3(n_572),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2117),
.Y(n_2280)
);

AOI22xp33_ASAP7_75t_SL g2281 ( 
.A1(n_2217),
.A2(n_608),
.B1(n_628),
.B2(n_604),
.Y(n_2281)
);

OA21x2_ASAP7_75t_L g2282 ( 
.A1(n_2160),
.A2(n_633),
.B(n_630),
.Y(n_2282)
);

AOI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_2217),
.A2(n_637),
.B1(n_640),
.B2(n_634),
.Y(n_2283)
);

INVx2_ASAP7_75t_SL g2284 ( 
.A(n_2141),
.Y(n_2284)
);

OAI22xp33_ASAP7_75t_L g2285 ( 
.A1(n_2191),
.A2(n_2221),
.B1(n_2212),
.B2(n_2232),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2117),
.Y(n_2286)
);

AO31x2_ASAP7_75t_L g2287 ( 
.A1(n_2084),
.A2(n_910),
.A3(n_912),
.B(n_895),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_2083),
.Y(n_2288)
);

INVx2_ASAP7_75t_L g2289 ( 
.A(n_2144),
.Y(n_2289)
);

AND2x2_ASAP7_75t_L g2290 ( 
.A(n_2138),
.B(n_14),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2083),
.B(n_15),
.Y(n_2291)
);

AO21x2_ASAP7_75t_L g2292 ( 
.A1(n_2084),
.A2(n_923),
.B(n_912),
.Y(n_2292)
);

OAI211xp5_ASAP7_75t_L g2293 ( 
.A1(n_2230),
.A2(n_644),
.B(n_646),
.C(n_642),
.Y(n_2293)
);

OAI21xp5_ASAP7_75t_L g2294 ( 
.A1(n_2193),
.A2(n_654),
.B(n_653),
.Y(n_2294)
);

AOI22xp33_ASAP7_75t_L g2295 ( 
.A1(n_2191),
.A2(n_2221),
.B1(n_2234),
.B2(n_2223),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2139),
.B(n_2140),
.Y(n_2296)
);

BUFx3_ASAP7_75t_L g2297 ( 
.A(n_2178),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_L g2298 ( 
.A1(n_2234),
.A2(n_674),
.B1(n_676),
.B2(n_658),
.Y(n_2298)
);

OR2x6_ASAP7_75t_L g2299 ( 
.A(n_2223),
.B(n_1452),
.Y(n_2299)
);

NAND3xp33_ASAP7_75t_L g2300 ( 
.A(n_2088),
.B(n_679),
.C(n_678),
.Y(n_2300)
);

OAI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2237),
.A2(n_707),
.B1(n_708),
.B2(n_680),
.Y(n_2301)
);

AOI21x1_ASAP7_75t_L g2302 ( 
.A1(n_2165),
.A2(n_925),
.B(n_923),
.Y(n_2302)
);

OAI21x1_ASAP7_75t_SL g2303 ( 
.A1(n_2182),
.A2(n_15),
.B(n_16),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_2223),
.A2(n_711),
.B1(n_713),
.B2(n_710),
.Y(n_2304)
);

AOI221xp5_ASAP7_75t_L g2305 ( 
.A1(n_2232),
.A2(n_721),
.B1(n_719),
.B2(n_716),
.C(n_19),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_2107),
.B(n_16),
.Y(n_2306)
);

OAI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2233),
.A2(n_21),
.B1(n_18),
.B2(n_20),
.Y(n_2307)
);

NOR3xp33_ASAP7_75t_L g2308 ( 
.A(n_2109),
.B(n_925),
.C(n_18),
.Y(n_2308)
);

AND2x4_ASAP7_75t_L g2309 ( 
.A(n_2175),
.B(n_20),
.Y(n_2309)
);

AND2x2_ASAP7_75t_L g2310 ( 
.A(n_2138),
.B(n_21),
.Y(n_2310)
);

AOI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2223),
.A2(n_889),
.B1(n_909),
.B2(n_897),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2118),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2179),
.B(n_24),
.Y(n_2313)
);

OAI211xp5_ASAP7_75t_L g2314 ( 
.A1(n_2231),
.A2(n_29),
.B(n_26),
.C(n_27),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2118),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2119),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2223),
.A2(n_909),
.B1(n_913),
.B2(n_897),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2119),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2120),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2179),
.B(n_26),
.Y(n_2320)
);

OA21x2_ASAP7_75t_L g2321 ( 
.A1(n_2127),
.A2(n_1276),
.B(n_1265),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2147),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2235),
.A2(n_909),
.B1(n_913),
.B2(n_897),
.Y(n_2323)
);

CKINVDCx20_ASAP7_75t_R g2324 ( 
.A(n_2178),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2120),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2122),
.Y(n_2326)
);

AOI21xp33_ASAP7_75t_L g2327 ( 
.A1(n_2218),
.A2(n_30),
.B(n_32),
.Y(n_2327)
);

BUFx12f_ASAP7_75t_L g2328 ( 
.A(n_2146),
.Y(n_2328)
);

INVx1_ASAP7_75t_SL g2329 ( 
.A(n_2180),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2147),
.Y(n_2330)
);

AOI221xp5_ASAP7_75t_L g2331 ( 
.A1(n_2233),
.A2(n_34),
.B1(n_30),
.B2(n_32),
.C(n_36),
.Y(n_2331)
);

INVx2_ASAP7_75t_L g2332 ( 
.A(n_2095),
.Y(n_2332)
);

AOI22xp33_ASAP7_75t_L g2333 ( 
.A1(n_2235),
.A2(n_2212),
.B1(n_2209),
.B2(n_2227),
.Y(n_2333)
);

AOI221xp5_ASAP7_75t_L g2334 ( 
.A1(n_2231),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.C(n_41),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2212),
.A2(n_2209),
.B1(n_2227),
.B2(n_2195),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2095),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2122),
.Y(n_2337)
);

AOI21x1_ASAP7_75t_L g2338 ( 
.A1(n_2165),
.A2(n_1279),
.B(n_1276),
.Y(n_2338)
);

CKINVDCx11_ASAP7_75t_R g2339 ( 
.A(n_2133),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2189),
.B(n_2199),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2212),
.A2(n_43),
.B1(n_39),
.B2(n_42),
.Y(n_2341)
);

INVx1_ASAP7_75t_SL g2342 ( 
.A(n_2180),
.Y(n_2342)
);

AOI22xp33_ASAP7_75t_SL g2343 ( 
.A1(n_2187),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_2343)
);

AOI22xp33_ASAP7_75t_SL g2344 ( 
.A1(n_2187),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_2141),
.Y(n_2345)
);

AOI22xp33_ASAP7_75t_L g2346 ( 
.A1(n_2212),
.A2(n_909),
.B1(n_913),
.B2(n_897),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2189),
.B(n_46),
.Y(n_2347)
);

OR2x2_ASAP7_75t_SL g2348 ( 
.A(n_2205),
.B(n_2146),
.Y(n_2348)
);

AND2x4_ASAP7_75t_L g2349 ( 
.A(n_2175),
.B(n_47),
.Y(n_2349)
);

OAI211xp5_ASAP7_75t_L g2350 ( 
.A1(n_2190),
.A2(n_50),
.B(n_47),
.C(n_48),
.Y(n_2350)
);

OAI22xp33_ASAP7_75t_L g2351 ( 
.A1(n_2205),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2199),
.B(n_51),
.Y(n_2352)
);

AND2x2_ASAP7_75t_L g2353 ( 
.A(n_2167),
.B(n_53),
.Y(n_2353)
);

AOI221xp5_ASAP7_75t_L g2354 ( 
.A1(n_2226),
.A2(n_59),
.B1(n_54),
.B2(n_58),
.C(n_60),
.Y(n_2354)
);

OAI211xp5_ASAP7_75t_L g2355 ( 
.A1(n_2240),
.A2(n_2172),
.B(n_2238),
.C(n_2190),
.Y(n_2355)
);

OR2x2_ASAP7_75t_L g2356 ( 
.A(n_2140),
.B(n_54),
.Y(n_2356)
);

AOI22xp33_ASAP7_75t_L g2357 ( 
.A1(n_2209),
.A2(n_909),
.B1(n_913),
.B2(n_897),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2204),
.B(n_58),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2204),
.B(n_61),
.Y(n_2359)
);

AOI22xp33_ASAP7_75t_L g2360 ( 
.A1(n_2209),
.A2(n_913),
.B1(n_930),
.B2(n_1279),
.Y(n_2360)
);

INVx2_ASAP7_75t_SL g2361 ( 
.A(n_2096),
.Y(n_2361)
);

OAI221xp5_ASAP7_75t_L g2362 ( 
.A1(n_2240),
.A2(n_64),
.B1(n_62),
.B2(n_63),
.C(n_65),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2123),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2123),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2095),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2340),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2261),
.Y(n_2367)
);

OR2x2_ASAP7_75t_L g2368 ( 
.A(n_2296),
.B(n_2201),
.Y(n_2368)
);

AND2x2_ASAP7_75t_L g2369 ( 
.A(n_2272),
.B(n_2329),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_SL g2370 ( 
.A(n_2324),
.B(n_2176),
.Y(n_2370)
);

HB1xp67_ASAP7_75t_L g2371 ( 
.A(n_2276),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2289),
.Y(n_2372)
);

OR2x2_ASAP7_75t_L g2373 ( 
.A(n_2251),
.B(n_2201),
.Y(n_2373)
);

AND2x2_ASAP7_75t_L g2374 ( 
.A(n_2329),
.B(n_2342),
.Y(n_2374)
);

INVxp67_ASAP7_75t_SL g2375 ( 
.A(n_2291),
.Y(n_2375)
);

NAND2x1p5_ASAP7_75t_L g2376 ( 
.A(n_2241),
.B(n_2188),
.Y(n_2376)
);

AND2x4_ASAP7_75t_L g2377 ( 
.A(n_2299),
.B(n_2241),
.Y(n_2377)
);

INVxp67_ASAP7_75t_L g2378 ( 
.A(n_2242),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2257),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2260),
.B(n_2148),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_2322),
.Y(n_2381)
);

AOI22xp33_ASAP7_75t_SL g2382 ( 
.A1(n_2350),
.A2(n_2164),
.B1(n_2203),
.B2(n_2146),
.Y(n_2382)
);

BUFx3_ASAP7_75t_L g2383 ( 
.A(n_2328),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2271),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2280),
.Y(n_2385)
);

AND2x2_ASAP7_75t_L g2386 ( 
.A(n_2342),
.B(n_2116),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2286),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2312),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2259),
.B(n_2148),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2291),
.B(n_2306),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2315),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2316),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2318),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_2306),
.B(n_2104),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2352),
.B(n_2159),
.Y(n_2395)
);

AND2x2_ASAP7_75t_L g2396 ( 
.A(n_2248),
.B(n_2116),
.Y(n_2396)
);

AND2x4_ASAP7_75t_L g2397 ( 
.A(n_2299),
.B(n_2181),
.Y(n_2397)
);

BUFx2_ASAP7_75t_L g2398 ( 
.A(n_2348),
.Y(n_2398)
);

AOI21xp5_ASAP7_75t_SL g2399 ( 
.A1(n_2264),
.A2(n_2220),
.B(n_2176),
.Y(n_2399)
);

INVx1_ASAP7_75t_SL g2400 ( 
.A(n_2339),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2330),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2284),
.B(n_2116),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2319),
.Y(n_2403)
);

AND2x4_ASAP7_75t_L g2404 ( 
.A(n_2299),
.B(n_2181),
.Y(n_2404)
);

AND2x2_ASAP7_75t_L g2405 ( 
.A(n_2345),
.B(n_2111),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2246),
.B(n_2111),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2313),
.B(n_2195),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2333),
.B(n_2158),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_2320),
.B(n_2149),
.Y(n_2409)
);

AND2x4_ASAP7_75t_SL g2410 ( 
.A(n_2269),
.B(n_2309),
.Y(n_2410)
);

AND2x4_ASAP7_75t_L g2411 ( 
.A(n_2275),
.B(n_2181),
.Y(n_2411)
);

INVxp67_ASAP7_75t_SL g2412 ( 
.A(n_2288),
.Y(n_2412)
);

INVx2_ASAP7_75t_L g2413 ( 
.A(n_2325),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2341),
.A2(n_2186),
.B1(n_2202),
.B2(n_2164),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2326),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2275),
.B(n_2158),
.Y(n_2416)
);

INVx1_ASAP7_75t_L g2417 ( 
.A(n_2337),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2363),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2335),
.B(n_2167),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2295),
.B(n_2177),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2364),
.Y(n_2421)
);

OAI21xp5_ASAP7_75t_L g2422 ( 
.A1(n_2355),
.A2(n_2285),
.B(n_2245),
.Y(n_2422)
);

INVx2_ASAP7_75t_SL g2423 ( 
.A(n_2297),
.Y(n_2423)
);

OR2x2_ASAP7_75t_L g2424 ( 
.A(n_2255),
.B(n_2149),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2243),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2247),
.Y(n_2426)
);

INVx2_ASAP7_75t_SL g2427 ( 
.A(n_2361),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2347),
.B(n_2156),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2332),
.Y(n_2429)
);

INVx3_ASAP7_75t_L g2430 ( 
.A(n_2336),
.Y(n_2430)
);

INVx3_ASAP7_75t_L g2431 ( 
.A(n_2365),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2273),
.Y(n_2432)
);

OR2x2_ASAP7_75t_L g2433 ( 
.A(n_2355),
.B(n_2202),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2356),
.Y(n_2434)
);

HB1xp67_ASAP7_75t_L g2435 ( 
.A(n_2292),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2292),
.Y(n_2436)
);

INVx2_ASAP7_75t_L g2437 ( 
.A(n_2269),
.Y(n_2437)
);

NOR2x1_ASAP7_75t_L g2438 ( 
.A(n_2309),
.B(n_2176),
.Y(n_2438)
);

AOI22xp33_ASAP7_75t_L g2439 ( 
.A1(n_2250),
.A2(n_2211),
.B1(n_2220),
.B2(n_2225),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2358),
.B(n_2077),
.Y(n_2440)
);

NOR2x1_ASAP7_75t_L g2441 ( 
.A(n_2349),
.B(n_2207),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2250),
.A2(n_2211),
.B1(n_2220),
.B2(n_2225),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2359),
.Y(n_2443)
);

OR2x2_ASAP7_75t_L g2444 ( 
.A(n_2277),
.B(n_2077),
.Y(n_2444)
);

AND2x2_ASAP7_75t_L g2445 ( 
.A(n_2256),
.B(n_2177),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2353),
.Y(n_2446)
);

INVxp67_ASAP7_75t_SL g2447 ( 
.A(n_2266),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2266),
.B(n_2078),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2249),
.A2(n_2220),
.B1(n_2225),
.B2(n_2203),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2302),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2349),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_2290),
.B(n_2156),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2310),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2321),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_2308),
.B(n_2163),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2321),
.Y(n_2456)
);

NAND3xp33_ASAP7_75t_L g2457 ( 
.A(n_2305),
.B(n_2215),
.C(n_2186),
.Y(n_2457)
);

AND2x2_ASAP7_75t_L g2458 ( 
.A(n_2244),
.B(n_2155),
.Y(n_2458)
);

OR2x2_ASAP7_75t_L g2459 ( 
.A(n_2282),
.B(n_2078),
.Y(n_2459)
);

BUFx2_ASAP7_75t_L g2460 ( 
.A(n_2282),
.Y(n_2460)
);

NAND2xp5_ASAP7_75t_L g2461 ( 
.A(n_2267),
.B(n_2163),
.Y(n_2461)
);

AND2x2_ASAP7_75t_L g2462 ( 
.A(n_2357),
.B(n_2155),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2287),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2360),
.B(n_2155),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2270),
.B(n_2181),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2258),
.B(n_2171),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2287),
.Y(n_2467)
);

INVxp67_ASAP7_75t_SL g2468 ( 
.A(n_2265),
.Y(n_2468)
);

AOI21xp33_ASAP7_75t_L g2469 ( 
.A1(n_2300),
.A2(n_2215),
.B(n_2181),
.Y(n_2469)
);

AOI22xp33_ASAP7_75t_L g2470 ( 
.A1(n_2249),
.A2(n_2214),
.B1(n_2215),
.B2(n_2146),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2343),
.B(n_2170),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2287),
.B(n_2079),
.Y(n_2472)
);

AND2x2_ASAP7_75t_L g2473 ( 
.A(n_2344),
.B(n_2171),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2303),
.Y(n_2474)
);

AND2x4_ASAP7_75t_SL g2475 ( 
.A(n_2278),
.B(n_2188),
.Y(n_2475)
);

HB1xp67_ASAP7_75t_L g2476 ( 
.A(n_2338),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2274),
.Y(n_2477)
);

INVx1_ASAP7_75t_L g2478 ( 
.A(n_2307),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2379),
.Y(n_2479)
);

AOI31xp33_ASAP7_75t_L g2480 ( 
.A1(n_2422),
.A2(n_2354),
.A3(n_2327),
.B(n_2334),
.Y(n_2480)
);

AOI22xp33_ASAP7_75t_L g2481 ( 
.A1(n_2457),
.A2(n_2305),
.B1(n_2254),
.B2(n_2253),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2384),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2385),
.Y(n_2483)
);

OAI211xp5_ASAP7_75t_L g2484 ( 
.A1(n_2399),
.A2(n_2382),
.B(n_2442),
.C(n_2439),
.Y(n_2484)
);

OAI31xp33_ASAP7_75t_SL g2485 ( 
.A1(n_2447),
.A2(n_2314),
.A3(n_2334),
.B(n_2354),
.Y(n_2485)
);

OAI22xp33_ASAP7_75t_L g2486 ( 
.A1(n_2414),
.A2(n_2362),
.B1(n_2274),
.B2(n_2188),
.Y(n_2486)
);

OAI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2382),
.A2(n_2362),
.B1(n_2283),
.B2(n_2331),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2376),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_2376),
.Y(n_2489)
);

NAND3xp33_ASAP7_75t_L g2490 ( 
.A(n_2399),
.B(n_2331),
.C(n_2327),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2387),
.Y(n_2491)
);

OAI21xp5_ASAP7_75t_L g2492 ( 
.A1(n_2447),
.A2(n_2281),
.B(n_2294),
.Y(n_2492)
);

OAI211xp5_ASAP7_75t_L g2493 ( 
.A1(n_2439),
.A2(n_2442),
.B(n_2470),
.C(n_2378),
.Y(n_2493)
);

OR2x2_ASAP7_75t_L g2494 ( 
.A(n_2444),
.B(n_2170),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2388),
.Y(n_2495)
);

OAI22xp5_ASAP7_75t_L g2496 ( 
.A1(n_2470),
.A2(n_2268),
.B1(n_2307),
.B2(n_2346),
.Y(n_2496)
);

INVxp67_ASAP7_75t_SL g2497 ( 
.A(n_2441),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2391),
.Y(n_2498)
);

OAI21x1_ASAP7_75t_L g2499 ( 
.A1(n_2438),
.A2(n_2087),
.B(n_2127),
.Y(n_2499)
);

AOI22xp33_ASAP7_75t_L g2500 ( 
.A1(n_2477),
.A2(n_2252),
.B1(n_2279),
.B2(n_2294),
.Y(n_2500)
);

OAI211xp5_ASAP7_75t_L g2501 ( 
.A1(n_2378),
.A2(n_2252),
.B(n_2293),
.C(n_2298),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2375),
.B(n_2085),
.Y(n_2502)
);

AOI222xp33_ASAP7_75t_L g2503 ( 
.A1(n_2477),
.A2(n_2351),
.B1(n_2263),
.B2(n_2301),
.C1(n_2262),
.C2(n_2304),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2375),
.B(n_2085),
.Y(n_2504)
);

NAND2xp5_ASAP7_75t_L g2505 ( 
.A(n_2478),
.B(n_2101),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2373),
.B(n_2174),
.Y(n_2506)
);

AOI22xp33_ASAP7_75t_L g2507 ( 
.A1(n_2460),
.A2(n_2469),
.B1(n_2398),
.B2(n_2408),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2383),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2392),
.Y(n_2509)
);

AO21x2_ASAP7_75t_L g2510 ( 
.A1(n_2412),
.A2(n_2263),
.B(n_2301),
.Y(n_2510)
);

NOR2xp67_ASAP7_75t_L g2511 ( 
.A(n_2371),
.B(n_2182),
.Y(n_2511)
);

INVx2_ASAP7_75t_SL g2512 ( 
.A(n_2410),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_2400),
.B(n_2214),
.Y(n_2513)
);

INVx3_ASAP7_75t_L g2514 ( 
.A(n_2383),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2393),
.Y(n_2515)
);

INVx5_ASAP7_75t_SL g2516 ( 
.A(n_2377),
.Y(n_2516)
);

NAND2xp33_ASAP7_75t_R g2517 ( 
.A(n_2473),
.B(n_2171),
.Y(n_2517)
);

AOI22xp33_ASAP7_75t_L g2518 ( 
.A1(n_2433),
.A2(n_2262),
.B1(n_2215),
.B2(n_2174),
.Y(n_2518)
);

AOI222xp33_ASAP7_75t_L g2519 ( 
.A1(n_2389),
.A2(n_2126),
.B1(n_2323),
.B2(n_2135),
.C1(n_2079),
.C2(n_2157),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2423),
.Y(n_2520)
);

AOI22xp33_ASAP7_75t_L g2521 ( 
.A1(n_2475),
.A2(n_2461),
.B1(n_2420),
.B2(n_2419),
.Y(n_2521)
);

AOI21xp5_ASAP7_75t_L g2522 ( 
.A1(n_2370),
.A2(n_2215),
.B(n_2157),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2371),
.B(n_2101),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2396),
.B(n_2173),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2369),
.B(n_2173),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_2466),
.Y(n_2526)
);

AOI222xp33_ASAP7_75t_L g2527 ( 
.A1(n_2475),
.A2(n_2126),
.B1(n_2135),
.B2(n_2157),
.C1(n_2192),
.C2(n_2183),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2403),
.Y(n_2528)
);

AOI21xp5_ASAP7_75t_L g2529 ( 
.A1(n_2455),
.A2(n_2157),
.B(n_2208),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_L g2530 ( 
.A(n_2434),
.B(n_2121),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2432),
.B(n_2102),
.Y(n_2531)
);

AO21x2_ASAP7_75t_L g2532 ( 
.A1(n_2412),
.A2(n_2136),
.B(n_2151),
.Y(n_2532)
);

OAI31xp33_ASAP7_75t_L g2533 ( 
.A1(n_2449),
.A2(n_2198),
.A3(n_2208),
.B(n_2105),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2443),
.B(n_2102),
.Y(n_2534)
);

BUFx2_ASAP7_75t_L g2535 ( 
.A(n_2427),
.Y(n_2535)
);

BUFx2_ASAP7_75t_L g2536 ( 
.A(n_2427),
.Y(n_2536)
);

INVxp67_ASAP7_75t_SL g2537 ( 
.A(n_2474),
.Y(n_2537)
);

INVx1_ASAP7_75t_L g2538 ( 
.A(n_2415),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_SL g2539 ( 
.A1(n_2474),
.A2(n_2097),
.B1(n_2166),
.B2(n_2206),
.Y(n_2539)
);

AO21x2_ASAP7_75t_L g2540 ( 
.A1(n_2468),
.A2(n_2136),
.B(n_2151),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2417),
.Y(n_2541)
);

AOI22xp33_ASAP7_75t_L g2542 ( 
.A1(n_2449),
.A2(n_2188),
.B1(n_2317),
.B2(n_2210),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2423),
.Y(n_2543)
);

AOI22xp33_ASAP7_75t_L g2544 ( 
.A1(n_2424),
.A2(n_2188),
.B1(n_2210),
.B2(n_2311),
.Y(n_2544)
);

NAND2xp33_ASAP7_75t_R g2545 ( 
.A(n_2374),
.B(n_2437),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2418),
.Y(n_2546)
);

AND2x2_ASAP7_75t_L g2547 ( 
.A(n_2458),
.B(n_2173),
.Y(n_2547)
);

INVxp67_ASAP7_75t_L g2548 ( 
.A(n_2437),
.Y(n_2548)
);

OAI22xp5_ASAP7_75t_SL g2549 ( 
.A1(n_2468),
.A2(n_2451),
.B1(n_2471),
.B2(n_2390),
.Y(n_2549)
);

AOI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2453),
.A2(n_2210),
.B1(n_2103),
.B2(n_2166),
.Y(n_2550)
);

NAND2xp33_ASAP7_75t_R g2551 ( 
.A(n_2451),
.B(n_62),
.Y(n_2551)
);

INVx1_ASAP7_75t_SL g2552 ( 
.A(n_2410),
.Y(n_2552)
);

OAI22xp5_ASAP7_75t_L g2553 ( 
.A1(n_2446),
.A2(n_2137),
.B1(n_2206),
.B2(n_2194),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2440),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2394),
.B(n_2097),
.Y(n_2555)
);

AND2x2_ASAP7_75t_L g2556 ( 
.A(n_2386),
.B(n_2145),
.Y(n_2556)
);

OAI221xp5_ASAP7_75t_L g2557 ( 
.A1(n_2380),
.A2(n_2459),
.B1(n_2448),
.B2(n_2407),
.C(n_2395),
.Y(n_2557)
);

OAI221xp5_ASAP7_75t_L g2558 ( 
.A1(n_2428),
.A2(n_2198),
.B1(n_2194),
.B2(n_2197),
.C(n_2166),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2402),
.B(n_2097),
.Y(n_2559)
);

BUFx3_ASAP7_75t_L g2560 ( 
.A(n_2405),
.Y(n_2560)
);

NOR2xp33_ASAP7_75t_R g2561 ( 
.A(n_2452),
.B(n_2097),
.Y(n_2561)
);

NOR2x1p5_ASAP7_75t_L g2562 ( 
.A(n_2409),
.B(n_2166),
.Y(n_2562)
);

OR2x2_ASAP7_75t_L g2563 ( 
.A(n_2368),
.B(n_2366),
.Y(n_2563)
);

OAI211xp5_ASAP7_75t_SL g2564 ( 
.A1(n_2425),
.A2(n_2152),
.B(n_2197),
.C(n_2154),
.Y(n_2564)
);

BUFx3_ASAP7_75t_L g2565 ( 
.A(n_2406),
.Y(n_2565)
);

NAND3xp33_ASAP7_75t_L g2566 ( 
.A(n_2450),
.B(n_2200),
.C(n_2103),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2480),
.B(n_2445),
.Y(n_2567)
);

INVx2_ASAP7_75t_L g2568 ( 
.A(n_2508),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2494),
.B(n_2366),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2508),
.B(n_2377),
.Y(n_2570)
);

BUFx2_ASAP7_75t_L g2571 ( 
.A(n_2497),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2479),
.Y(n_2572)
);

AND2x2_ASAP7_75t_L g2573 ( 
.A(n_2514),
.B(n_2377),
.Y(n_2573)
);

AOI22xp5_ASAP7_75t_L g2574 ( 
.A1(n_2487),
.A2(n_2462),
.B1(n_2464),
.B2(n_2435),
.Y(n_2574)
);

NAND3xp33_ASAP7_75t_L g2575 ( 
.A(n_2484),
.B(n_2435),
.C(n_2436),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2482),
.Y(n_2576)
);

AOI211xp5_ASAP7_75t_L g2577 ( 
.A1(n_2490),
.A2(n_2465),
.B(n_2404),
.C(n_2397),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_SL g2578 ( 
.A(n_2485),
.B(n_2465),
.Y(n_2578)
);

NAND3xp33_ASAP7_75t_L g2579 ( 
.A(n_2493),
.B(n_2436),
.C(n_2476),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2514),
.B(n_2552),
.Y(n_2580)
);

NAND4xp75_ASAP7_75t_L g2581 ( 
.A(n_2492),
.B(n_2416),
.C(n_2467),
.D(n_2463),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2481),
.B(n_2476),
.C(n_2426),
.Y(n_2582)
);

INVxp67_ASAP7_75t_SL g2583 ( 
.A(n_2545),
.Y(n_2583)
);

OR2x2_ASAP7_75t_L g2584 ( 
.A(n_2548),
.B(n_2367),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2565),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2483),
.Y(n_2586)
);

INVxp67_ASAP7_75t_L g2587 ( 
.A(n_2551),
.Y(n_2587)
);

AND2x2_ASAP7_75t_L g2588 ( 
.A(n_2512),
.B(n_2416),
.Y(n_2588)
);

NAND4xp25_ASAP7_75t_L g2589 ( 
.A(n_2507),
.B(n_2465),
.C(n_2411),
.D(n_2404),
.Y(n_2589)
);

NOR3xp33_ASAP7_75t_L g2590 ( 
.A(n_2549),
.B(n_2501),
.C(n_2492),
.Y(n_2590)
);

NOR2x1_ASAP7_75t_R g2591 ( 
.A(n_2526),
.B(n_2166),
.Y(n_2591)
);

INVx2_ASAP7_75t_L g2592 ( 
.A(n_2516),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2525),
.B(n_2411),
.Y(n_2593)
);

AND2x4_ASAP7_75t_L g2594 ( 
.A(n_2511),
.B(n_2535),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2487),
.A2(n_2510),
.B1(n_2486),
.B2(n_2500),
.Y(n_2595)
);

BUFx6f_ASAP7_75t_L g2596 ( 
.A(n_2536),
.Y(n_2596)
);

NOR3xp33_ASAP7_75t_L g2597 ( 
.A(n_2557),
.B(n_2411),
.C(n_2429),
.Y(n_2597)
);

AND2x2_ASAP7_75t_L g2598 ( 
.A(n_2516),
.B(n_2397),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2513),
.B(n_2429),
.Y(n_2599)
);

INVxp67_ASAP7_75t_L g2600 ( 
.A(n_2517),
.Y(n_2600)
);

OR2x2_ASAP7_75t_L g2601 ( 
.A(n_2563),
.B(n_2367),
.Y(n_2601)
);

NOR3xp33_ASAP7_75t_L g2602 ( 
.A(n_2537),
.B(n_2381),
.C(n_2372),
.Y(n_2602)
);

OAI211xp5_ASAP7_75t_L g2603 ( 
.A1(n_2533),
.A2(n_2521),
.B(n_2503),
.C(n_2542),
.Y(n_2603)
);

INVx3_ASAP7_75t_L g2604 ( 
.A(n_2516),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2520),
.B(n_2372),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2510),
.A2(n_2404),
.B1(n_2397),
.B2(n_2413),
.Y(n_2606)
);

AOI22xp33_ASAP7_75t_SL g2607 ( 
.A1(n_2496),
.A2(n_2430),
.B1(n_2431),
.B2(n_2103),
.Y(n_2607)
);

OAI211xp5_ASAP7_75t_SL g2608 ( 
.A1(n_2518),
.A2(n_2401),
.B(n_2381),
.C(n_2413),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2491),
.Y(n_2609)
);

AOI22xp33_ASAP7_75t_L g2610 ( 
.A1(n_2560),
.A2(n_2421),
.B1(n_2401),
.B2(n_2430),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2519),
.A2(n_2421),
.B1(n_2431),
.B2(n_2430),
.Y(n_2611)
);

NAND3xp33_ASAP7_75t_L g2612 ( 
.A(n_2496),
.B(n_2456),
.C(n_2454),
.Y(n_2612)
);

AO21x2_ASAP7_75t_L g2613 ( 
.A1(n_2540),
.A2(n_2456),
.B(n_2454),
.Y(n_2613)
);

OR2x2_ASAP7_75t_L g2614 ( 
.A(n_2530),
.B(n_2472),
.Y(n_2614)
);

NAND3xp33_ASAP7_75t_L g2615 ( 
.A(n_2543),
.B(n_2431),
.C(n_2200),
.Y(n_2615)
);

NAND4xp75_ASAP7_75t_L g2616 ( 
.A(n_2522),
.B(n_2103),
.C(n_2169),
.D(n_2192),
.Y(n_2616)
);

OR2x2_ASAP7_75t_L g2617 ( 
.A(n_2530),
.B(n_2090),
.Y(n_2617)
);

NAND3xp33_ASAP7_75t_L g2618 ( 
.A(n_2566),
.B(n_2210),
.C(n_2110),
.Y(n_2618)
);

NAND4xp75_ASAP7_75t_L g2619 ( 
.A(n_2529),
.B(n_2169),
.C(n_2183),
.D(n_2152),
.Y(n_2619)
);

NAND4xp75_ASAP7_75t_L g2620 ( 
.A(n_2488),
.B(n_2134),
.C(n_2131),
.D(n_2154),
.Y(n_2620)
);

NAND3xp33_ASAP7_75t_L g2621 ( 
.A(n_2550),
.B(n_2210),
.C(n_2110),
.Y(n_2621)
);

AOI211x1_ASAP7_75t_L g2622 ( 
.A1(n_2558),
.A2(n_2505),
.B(n_2553),
.C(n_2504),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2554),
.B(n_2505),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2495),
.Y(n_2624)
);

NAND3xp33_ASAP7_75t_L g2625 ( 
.A(n_2544),
.B(n_2090),
.C(n_2131),
.Y(n_2625)
);

NAND3xp33_ASAP7_75t_L g2626 ( 
.A(n_2498),
.B(n_2134),
.C(n_2114),
.Y(n_2626)
);

NOR3xp33_ASAP7_75t_L g2627 ( 
.A(n_2539),
.B(n_2236),
.C(n_2087),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2547),
.B(n_2559),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2509),
.Y(n_2629)
);

OR2x2_ASAP7_75t_L g2630 ( 
.A(n_2506),
.B(n_2124),
.Y(n_2630)
);

AOI221xp5_ASAP7_75t_L g2631 ( 
.A1(n_2515),
.A2(n_2114),
.B1(n_2113),
.B2(n_2124),
.C(n_2142),
.Y(n_2631)
);

AO21x2_ASAP7_75t_L g2632 ( 
.A1(n_2540),
.A2(n_2129),
.B(n_2236),
.Y(n_2632)
);

AND2x2_ASAP7_75t_L g2633 ( 
.A(n_2524),
.B(n_2153),
.Y(n_2633)
);

AND4x1_ASAP7_75t_L g2634 ( 
.A(n_2555),
.B(n_2527),
.C(n_2538),
.D(n_2528),
.Y(n_2634)
);

NOR3xp33_ASAP7_75t_L g2635 ( 
.A(n_2489),
.B(n_2546),
.C(n_2541),
.Y(n_2635)
);

NOR2x1_ASAP7_75t_L g2636 ( 
.A(n_2532),
.B(n_2562),
.Y(n_2636)
);

AOI211x1_ASAP7_75t_L g2637 ( 
.A1(n_2553),
.A2(n_2129),
.B(n_2099),
.C(n_2185),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2556),
.B(n_2531),
.Y(n_2638)
);

XNOR2x1_ASAP7_75t_L g2639 ( 
.A(n_2499),
.B(n_63),
.Y(n_2639)
);

NAND3xp33_ASAP7_75t_L g2640 ( 
.A(n_2502),
.B(n_2113),
.C(n_2142),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2531),
.B(n_2089),
.Y(n_2641)
);

AND2x4_ASAP7_75t_L g2642 ( 
.A(n_2532),
.B(n_2105),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2561),
.B(n_2153),
.Y(n_2643)
);

NAND3xp33_ASAP7_75t_L g2644 ( 
.A(n_2502),
.B(n_2086),
.C(n_2089),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2504),
.B(n_2153),
.Y(n_2645)
);

NOR2xp33_ASAP7_75t_L g2646 ( 
.A(n_2534),
.B(n_2092),
.Y(n_2646)
);

NAND3xp33_ASAP7_75t_L g2647 ( 
.A(n_2534),
.B(n_2086),
.C(n_2092),
.Y(n_2647)
);

OR2x2_ASAP7_75t_L g2648 ( 
.A(n_2523),
.B(n_2100),
.Y(n_2648)
);

OAI31xp33_ASAP7_75t_L g2649 ( 
.A1(n_2590),
.A2(n_2564),
.A3(n_2523),
.B(n_2137),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2596),
.Y(n_2650)
);

BUFx2_ASAP7_75t_L g2651 ( 
.A(n_2596),
.Y(n_2651)
);

OAI33xp33_ASAP7_75t_L g2652 ( 
.A1(n_2575),
.A2(n_2579),
.A3(n_2567),
.B1(n_2578),
.B2(n_2582),
.B3(n_2612),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2596),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2572),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2587),
.B(n_2100),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2576),
.Y(n_2656)
);

NAND2xp33_ASAP7_75t_L g2657 ( 
.A(n_2595),
.B(n_2137),
.Y(n_2657)
);

CKINVDCx16_ASAP7_75t_R g2658 ( 
.A(n_2580),
.Y(n_2658)
);

OAI221xp5_ASAP7_75t_L g2659 ( 
.A1(n_2634),
.A2(n_2106),
.B1(n_2108),
.B2(n_2185),
.C(n_2099),
.Y(n_2659)
);

INVx4_ASAP7_75t_L g2660 ( 
.A(n_2604),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2570),
.B(n_2106),
.Y(n_2661)
);

INVx4_ASAP7_75t_L g2662 ( 
.A(n_2604),
.Y(n_2662)
);

OAI33xp33_ASAP7_75t_L g2663 ( 
.A1(n_2586),
.A2(n_2629),
.A3(n_2624),
.B1(n_2609),
.B2(n_2623),
.B3(n_2605),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2569),
.Y(n_2664)
);

BUFx2_ASAP7_75t_L g2665 ( 
.A(n_2594),
.Y(n_2665)
);

OA211x2_ASAP7_75t_L g2666 ( 
.A1(n_2600),
.A2(n_66),
.B(n_64),
.C(n_65),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2584),
.Y(n_2667)
);

INVxp67_ASAP7_75t_L g2668 ( 
.A(n_2571),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2573),
.B(n_2108),
.Y(n_2669)
);

AND2x4_ASAP7_75t_L g2670 ( 
.A(n_2594),
.B(n_2098),
.Y(n_2670)
);

AND2x4_ASAP7_75t_SL g2671 ( 
.A(n_2568),
.B(n_1452),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2613),
.Y(n_2672)
);

OAI211xp5_ASAP7_75t_L g2673 ( 
.A1(n_2622),
.A2(n_2574),
.B(n_2603),
.C(n_2606),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2628),
.B(n_2098),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2588),
.B(n_2082),
.Y(n_2675)
);

OR2x2_ASAP7_75t_L g2676 ( 
.A(n_2638),
.B(n_2168),
.Y(n_2676)
);

NOR3xp33_ASAP7_75t_L g2677 ( 
.A(n_2581),
.B(n_66),
.C(n_67),
.Y(n_2677)
);

AOI22xp33_ASAP7_75t_SL g2678 ( 
.A1(n_2583),
.A2(n_2639),
.B1(n_2634),
.B2(n_2599),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2601),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2613),
.Y(n_2680)
);

NAND3xp33_ASAP7_75t_SL g2681 ( 
.A(n_2574),
.B(n_68),
.C(n_69),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2642),
.Y(n_2682)
);

OAI33xp33_ASAP7_75t_L g2683 ( 
.A1(n_2614),
.A2(n_69),
.A3(n_70),
.B1(n_71),
.B2(n_72),
.B3(n_75),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2598),
.B(n_2082),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2648),
.Y(n_2685)
);

OAI31xp33_ASAP7_75t_L g2686 ( 
.A1(n_2589),
.A2(n_72),
.A3(n_70),
.B(n_71),
.Y(n_2686)
);

AND2x4_ASAP7_75t_SL g2687 ( 
.A(n_2592),
.B(n_1452),
.Y(n_2687)
);

OR2x2_ASAP7_75t_L g2688 ( 
.A(n_2585),
.B(n_2168),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2641),
.Y(n_2689)
);

NAND4xp25_ASAP7_75t_L g2690 ( 
.A(n_2622),
.B(n_79),
.C(n_77),
.D(n_78),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2642),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2646),
.Y(n_2692)
);

AND2x2_ASAP7_75t_L g2693 ( 
.A(n_2593),
.B(n_2643),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2602),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2635),
.Y(n_2695)
);

OR2x6_ASAP7_75t_L g2696 ( 
.A(n_2636),
.B(n_2112),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2640),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2632),
.Y(n_2698)
);

AOI221xp5_ASAP7_75t_L g2699 ( 
.A1(n_2611),
.A2(n_2168),
.B1(n_80),
.B2(n_81),
.C(n_82),
.Y(n_2699)
);

NAND3xp33_ASAP7_75t_L g2700 ( 
.A(n_2607),
.B(n_78),
.C(n_81),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2632),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2620),
.Y(n_2702)
);

AOI211xp5_ASAP7_75t_L g2703 ( 
.A1(n_2597),
.A2(n_2591),
.B(n_2577),
.C(n_2608),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2633),
.B(n_2130),
.Y(n_2704)
);

OAI22xp5_ASAP7_75t_L g2705 ( 
.A1(n_2619),
.A2(n_2130),
.B1(n_2150),
.B2(n_2112),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2610),
.B(n_83),
.Y(n_2706)
);

INVx4_ASAP7_75t_L g2707 ( 
.A(n_2591),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2616),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2645),
.B(n_2130),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2617),
.B(n_2150),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2658),
.B(n_2678),
.Y(n_2711)
);

AND2x4_ASAP7_75t_L g2712 ( 
.A(n_2665),
.B(n_2615),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2678),
.B(n_2627),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2672),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2672),
.Y(n_2715)
);

AND2x2_ASAP7_75t_L g2716 ( 
.A(n_2693),
.B(n_2630),
.Y(n_2716)
);

OAI31xp33_ASAP7_75t_L g2717 ( 
.A1(n_2673),
.A2(n_2621),
.A3(n_2618),
.B(n_2625),
.Y(n_2717)
);

XNOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2666),
.B(n_85),
.Y(n_2718)
);

NOR2x1_ASAP7_75t_L g2719 ( 
.A(n_2690),
.B(n_2626),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2653),
.B(n_2631),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2700),
.A2(n_2637),
.B1(n_2644),
.B2(n_2647),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2680),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2680),
.Y(n_2723)
);

INVxp67_ASAP7_75t_SL g2724 ( 
.A(n_2668),
.Y(n_2724)
);

AO22x1_ASAP7_75t_L g2725 ( 
.A1(n_2677),
.A2(n_2637),
.B1(n_87),
.B2(n_85),
.Y(n_2725)
);

AOI32xp33_ASAP7_75t_L g2726 ( 
.A1(n_2677),
.A2(n_2162),
.A3(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2668),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2650),
.Y(n_2728)
);

OAI211xp5_ASAP7_75t_SL g2729 ( 
.A1(n_2703),
.A2(n_91),
.B(n_86),
.C(n_90),
.Y(n_2729)
);

A2O1A1Ixp33_ASAP7_75t_L g2730 ( 
.A1(n_2686),
.A2(n_2196),
.B(n_2162),
.C(n_2128),
.Y(n_2730)
);

OR2x2_ASAP7_75t_L g2731 ( 
.A(n_2681),
.B(n_86),
.Y(n_2731)
);

OAI322xp33_ASAP7_75t_L g2732 ( 
.A1(n_2659),
.A2(n_91),
.A3(n_92),
.B1(n_95),
.B2(n_96),
.C1(n_98),
.C2(n_99),
.Y(n_2732)
);

INVx1_ASAP7_75t_L g2733 ( 
.A(n_2651),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2679),
.Y(n_2734)
);

XNOR2x1_ASAP7_75t_L g2735 ( 
.A(n_2695),
.B(n_92),
.Y(n_2735)
);

OAI332xp33_ASAP7_75t_L g2736 ( 
.A1(n_2708),
.A2(n_95),
.A3(n_99),
.B1(n_101),
.B2(n_104),
.B3(n_108),
.C1(n_110),
.C2(n_112),
.Y(n_2736)
);

AND2x4_ASAP7_75t_L g2737 ( 
.A(n_2653),
.B(n_2150),
.Y(n_2737)
);

AND2x4_ASAP7_75t_L g2738 ( 
.A(n_2662),
.B(n_101),
.Y(n_2738)
);

AOI32xp33_ASAP7_75t_L g2739 ( 
.A1(n_2699),
.A2(n_110),
.A3(n_113),
.B1(n_115),
.B2(n_116),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2660),
.B(n_113),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2667),
.Y(n_2741)
);

AND2x2_ASAP7_75t_L g2742 ( 
.A(n_2660),
.B(n_117),
.Y(n_2742)
);

AOI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2652),
.A2(n_2196),
.B1(n_2128),
.B2(n_119),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_L g2744 ( 
.A(n_2694),
.B(n_117),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2664),
.B(n_2662),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2662),
.B(n_118),
.Y(n_2746)
);

INVx2_ASAP7_75t_SL g2747 ( 
.A(n_2682),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2682),
.Y(n_2748)
);

OAI222xp33_ASAP7_75t_L g2749 ( 
.A1(n_2708),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.C1(n_123),
.C2(n_125),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2685),
.B(n_2692),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2655),
.Y(n_2751)
);

INVxp67_ASAP7_75t_L g2752 ( 
.A(n_2706),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2707),
.B(n_120),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2691),
.B(n_123),
.Y(n_2754)
);

XNOR2x2_ASAP7_75t_L g2755 ( 
.A(n_2652),
.B(n_125),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2691),
.Y(n_2756)
);

OR2x6_ASAP7_75t_L g2757 ( 
.A(n_2707),
.B(n_126),
.Y(n_2757)
);

OR2x2_ASAP7_75t_L g2758 ( 
.A(n_2728),
.B(n_2697),
.Y(n_2758)
);

OR2x2_ASAP7_75t_L g2759 ( 
.A(n_2733),
.B(n_2689),
.Y(n_2759)
);

INVx1_ASAP7_75t_SL g2760 ( 
.A(n_2712),
.Y(n_2760)
);

AND2x2_ASAP7_75t_L g2761 ( 
.A(n_2716),
.B(n_2702),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2724),
.B(n_2687),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2756),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2748),
.Y(n_2764)
);

NOR2xp67_ASAP7_75t_L g2765 ( 
.A(n_2747),
.B(n_2702),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2712),
.Y(n_2766)
);

INVx3_ASAP7_75t_L g2767 ( 
.A(n_2738),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2725),
.B(n_2687),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2714),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2711),
.B(n_2663),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2753),
.B(n_2669),
.Y(n_2771)
);

HB1xp67_ASAP7_75t_L g2772 ( 
.A(n_2757),
.Y(n_2772)
);

OAI31xp33_ASAP7_75t_L g2773 ( 
.A1(n_2729),
.A2(n_2649),
.A3(n_2705),
.B(n_2701),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2715),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2726),
.B(n_2698),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2727),
.B(n_2671),
.Y(n_2776)
);

INVx1_ASAP7_75t_SL g2777 ( 
.A(n_2718),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2722),
.Y(n_2778)
);

NAND2xp33_ASAP7_75t_R g2779 ( 
.A(n_2757),
.B(n_2696),
.Y(n_2779)
);

INVxp67_ASAP7_75t_L g2780 ( 
.A(n_2740),
.Y(n_2780)
);

NAND2xp33_ASAP7_75t_SL g2781 ( 
.A(n_2713),
.B(n_2698),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2738),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2745),
.B(n_2663),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2723),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2746),
.Y(n_2785)
);

HB1xp67_ASAP7_75t_L g2786 ( 
.A(n_2742),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2754),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2726),
.B(n_2654),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2741),
.B(n_2734),
.Y(n_2789)
);

OR2x2_ASAP7_75t_L g2790 ( 
.A(n_2720),
.B(n_2656),
.Y(n_2790)
);

INVx3_ASAP7_75t_L g2791 ( 
.A(n_2755),
.Y(n_2791)
);

AOI211xp5_ASAP7_75t_L g2792 ( 
.A1(n_2732),
.A2(n_2657),
.B(n_2683),
.C(n_2701),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2750),
.Y(n_2793)
);

AND2x4_ASAP7_75t_SL g2794 ( 
.A(n_2751),
.B(n_2670),
.Y(n_2794)
);

NOR2xp33_ASAP7_75t_SL g2795 ( 
.A(n_2749),
.B(n_2683),
.Y(n_2795)
);

OAI221xp5_ASAP7_75t_L g2796 ( 
.A1(n_2770),
.A2(n_2717),
.B1(n_2743),
.B2(n_2739),
.C(n_2657),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2767),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2760),
.B(n_2719),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2767),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2786),
.Y(n_2800)
);

OR2x2_ASAP7_75t_L g2801 ( 
.A(n_2777),
.B(n_2744),
.Y(n_2801)
);

OAI21xp33_ASAP7_75t_L g2802 ( 
.A1(n_2770),
.A2(n_2719),
.B(n_2752),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2772),
.Y(n_2803)
);

NAND2x1_ASAP7_75t_L g2804 ( 
.A(n_2767),
.B(n_2670),
.Y(n_2804)
);

INVxp67_ASAP7_75t_L g2805 ( 
.A(n_2779),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2791),
.B(n_2735),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2766),
.B(n_2731),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2791),
.B(n_2739),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2794),
.Y(n_2809)
);

NOR3xp33_ASAP7_75t_L g2810 ( 
.A(n_2791),
.B(n_2736),
.C(n_2721),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2761),
.B(n_2661),
.Y(n_2811)
);

NOR2x1_ASAP7_75t_L g2812 ( 
.A(n_2775),
.B(n_2696),
.Y(n_2812)
);

NOR2x1_ASAP7_75t_L g2813 ( 
.A(n_2775),
.B(n_2696),
.Y(n_2813)
);

INVx2_ASAP7_75t_L g2814 ( 
.A(n_2766),
.Y(n_2814)
);

AND2x2_ASAP7_75t_L g2815 ( 
.A(n_2771),
.B(n_2671),
.Y(n_2815)
);

NOR4xp25_ASAP7_75t_L g2816 ( 
.A(n_2783),
.B(n_2730),
.C(n_2688),
.D(n_2709),
.Y(n_2816)
);

NAND3xp33_ASAP7_75t_L g2817 ( 
.A(n_2781),
.B(n_2676),
.C(n_2737),
.Y(n_2817)
);

INVxp67_ASAP7_75t_L g2818 ( 
.A(n_2779),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2785),
.B(n_2684),
.Y(n_2819)
);

OAI21xp33_ASAP7_75t_L g2820 ( 
.A1(n_2795),
.A2(n_2670),
.B(n_2675),
.Y(n_2820)
);

INVx2_ASAP7_75t_SL g2821 ( 
.A(n_2794),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2782),
.Y(n_2822)
);

NAND2x1p5_ASAP7_75t_L g2823 ( 
.A(n_2782),
.B(n_2737),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2788),
.B(n_2674),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2765),
.B(n_2704),
.Y(n_2825)
);

NOR4xp25_ASAP7_75t_L g2826 ( 
.A(n_2783),
.B(n_2710),
.C(n_129),
.D(n_127),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2758),
.Y(n_2827)
);

A2O1A1Ixp33_ASAP7_75t_L g2828 ( 
.A1(n_2810),
.A2(n_2792),
.B(n_2773),
.C(n_2781),
.Y(n_2828)
);

AND2x2_ASAP7_75t_L g2829 ( 
.A(n_2811),
.B(n_2780),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2797),
.Y(n_2830)
);

O2A1O1Ixp33_ASAP7_75t_SL g2831 ( 
.A1(n_2808),
.A2(n_2804),
.B(n_2806),
.C(n_2768),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2799),
.Y(n_2832)
);

OAI21xp33_ASAP7_75t_L g2833 ( 
.A1(n_2806),
.A2(n_2762),
.B(n_2776),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2798),
.B(n_2776),
.Y(n_2834)
);

INVx2_ASAP7_75t_SL g2835 ( 
.A(n_2809),
.Y(n_2835)
);

AOI222xp33_ASAP7_75t_L g2836 ( 
.A1(n_2796),
.A2(n_2802),
.B1(n_2808),
.B2(n_2818),
.C1(n_2805),
.C2(n_2812),
.Y(n_2836)
);

OAI21xp5_ASAP7_75t_SL g2837 ( 
.A1(n_2803),
.A2(n_2793),
.B(n_2764),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2823),
.Y(n_2838)
);

AOI31xp33_ASAP7_75t_L g2839 ( 
.A1(n_2821),
.A2(n_2827),
.A3(n_2801),
.B(n_2800),
.Y(n_2839)
);

AND2x4_ASAP7_75t_SL g2840 ( 
.A(n_2815),
.B(n_2814),
.Y(n_2840)
);

AND2x4_ASAP7_75t_L g2841 ( 
.A(n_2822),
.B(n_2789),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2813),
.A2(n_2790),
.B1(n_2789),
.B2(n_2787),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2826),
.B(n_2819),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2826),
.B(n_2763),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2823),
.Y(n_2845)
);

OR2x2_ASAP7_75t_L g2846 ( 
.A(n_2807),
.B(n_2759),
.Y(n_2846)
);

OAI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_2824),
.A2(n_2774),
.B1(n_2778),
.B2(n_2769),
.Y(n_2847)
);

AOI211xp5_ASAP7_75t_L g2848 ( 
.A1(n_2816),
.A2(n_2820),
.B(n_2825),
.C(n_2817),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2817),
.Y(n_2849)
);

NAND2x1_ASAP7_75t_L g2850 ( 
.A(n_2816),
.B(n_2784),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2797),
.B(n_128),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2797),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2835),
.Y(n_2853)
);

A2O1A1Ixp33_ASAP7_75t_L g2854 ( 
.A1(n_2850),
.A2(n_130),
.B(n_128),
.C(n_129),
.Y(n_2854)
);

XNOR2x1_ASAP7_75t_L g2855 ( 
.A(n_2834),
.B(n_130),
.Y(n_2855)
);

INVx1_ASAP7_75t_SL g2856 ( 
.A(n_2846),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2841),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2841),
.Y(n_2858)
);

OAI21xp33_ASAP7_75t_L g2859 ( 
.A1(n_2828),
.A2(n_132),
.B(n_133),
.Y(n_2859)
);

AND2x2_ASAP7_75t_L g2860 ( 
.A(n_2840),
.B(n_2829),
.Y(n_2860)
);

AOI321xp33_ASAP7_75t_L g2861 ( 
.A1(n_2848),
.A2(n_133),
.A3(n_135),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2839),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2830),
.Y(n_2863)
);

AO21x1_ASAP7_75t_L g2864 ( 
.A1(n_2849),
.A2(n_136),
.B(n_139),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2832),
.B(n_140),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2852),
.Y(n_2866)
);

OAI32xp33_ASAP7_75t_L g2867 ( 
.A1(n_2844),
.A2(n_2843),
.A3(n_2845),
.B1(n_2838),
.B2(n_2833),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2851),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2847),
.Y(n_2869)
);

XNOR2xp5_ASAP7_75t_L g2870 ( 
.A(n_2842),
.B(n_142),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_SL g2871 ( 
.A(n_2842),
.B(n_142),
.Y(n_2871)
);

BUFx2_ASAP7_75t_L g2872 ( 
.A(n_2857),
.Y(n_2872)
);

NOR2x1_ASAP7_75t_L g2873 ( 
.A(n_2858),
.B(n_2837),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2860),
.B(n_2836),
.Y(n_2874)
);

BUFx2_ASAP7_75t_R g2875 ( 
.A(n_2862),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_2856),
.Y(n_2876)
);

OAI221xp5_ASAP7_75t_L g2877 ( 
.A1(n_2861),
.A2(n_2831),
.B1(n_144),
.B2(n_145),
.C(n_146),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_SL g2878 ( 
.A(n_2856),
.B(n_1455),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2864),
.Y(n_2879)
);

NOR3x1_ASAP7_75t_L g2880 ( 
.A(n_2869),
.B(n_143),
.C(n_145),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2853),
.Y(n_2881)
);

INVx2_ASAP7_75t_SL g2882 ( 
.A(n_2865),
.Y(n_2882)
);

NAND2xp5_ASAP7_75t_L g2883 ( 
.A(n_2854),
.B(n_2870),
.Y(n_2883)
);

AOI211xp5_ASAP7_75t_L g2884 ( 
.A1(n_2871),
.A2(n_149),
.B(n_147),
.C(n_148),
.Y(n_2884)
);

INVxp67_ASAP7_75t_L g2885 ( 
.A(n_2872),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2876),
.B(n_2855),
.Y(n_2886)
);

OA22x2_ASAP7_75t_L g2887 ( 
.A1(n_2879),
.A2(n_2859),
.B1(n_2871),
.B2(n_2866),
.Y(n_2887)
);

OAI21xp33_ASAP7_75t_L g2888 ( 
.A1(n_2875),
.A2(n_2867),
.B(n_2863),
.Y(n_2888)
);

NOR2x1_ASAP7_75t_L g2889 ( 
.A(n_2873),
.B(n_2868),
.Y(n_2889)
);

NOR3x1_ASAP7_75t_L g2890 ( 
.A(n_2877),
.B(n_2882),
.C(n_2883),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2874),
.B(n_2861),
.Y(n_2891)
);

OAI21xp33_ASAP7_75t_L g2892 ( 
.A1(n_2881),
.A2(n_147),
.B(n_150),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2880),
.Y(n_2893)
);

AOI211xp5_ASAP7_75t_L g2894 ( 
.A1(n_2884),
.A2(n_150),
.B(n_151),
.C(n_152),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2884),
.B(n_151),
.Y(n_2895)
);

NOR2xp67_ASAP7_75t_L g2896 ( 
.A(n_2878),
.B(n_153),
.Y(n_2896)
);

OAI21xp33_ASAP7_75t_L g2897 ( 
.A1(n_2875),
.A2(n_154),
.B(n_156),
.Y(n_2897)
);

AOI211xp5_ASAP7_75t_SL g2898 ( 
.A1(n_2888),
.A2(n_159),
.B(n_161),
.C(n_162),
.Y(n_2898)
);

OR2x2_ASAP7_75t_L g2899 ( 
.A(n_2891),
.B(n_159),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2885),
.B(n_162),
.Y(n_2900)
);

OAI21xp5_ASAP7_75t_SL g2901 ( 
.A1(n_2889),
.A2(n_163),
.B(n_164),
.Y(n_2901)
);

INVxp67_ASAP7_75t_L g2902 ( 
.A(n_2895),
.Y(n_2902)
);

XOR2xp5_ASAP7_75t_L g2903 ( 
.A(n_2886),
.B(n_163),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2887),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_2893),
.B(n_165),
.Y(n_2905)
);

AND2x2_ASAP7_75t_L g2906 ( 
.A(n_2890),
.B(n_166),
.Y(n_2906)
);

INVxp67_ASAP7_75t_L g2907 ( 
.A(n_2897),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2892),
.Y(n_2908)
);

OR2x2_ASAP7_75t_L g2909 ( 
.A(n_2896),
.B(n_2894),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_SL g2910 ( 
.A(n_2889),
.B(n_1455),
.Y(n_2910)
);

NAND4xp25_ASAP7_75t_L g2911 ( 
.A(n_2888),
.B(n_167),
.C(n_169),
.D(n_170),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2885),
.B(n_171),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2885),
.B(n_172),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2885),
.B(n_172),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2903),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_2911),
.B(n_173),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_SL g2917 ( 
.A1(n_2904),
.A2(n_2907),
.B1(n_2908),
.B2(n_2909),
.Y(n_2917)
);

OAI31xp33_ASAP7_75t_L g2918 ( 
.A1(n_2901),
.A2(n_173),
.A3(n_174),
.B(n_175),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2906),
.Y(n_2919)
);

AO22x2_ASAP7_75t_L g2920 ( 
.A1(n_2899),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_2920)
);

NOR2xp33_ASAP7_75t_L g2921 ( 
.A(n_2911),
.B(n_176),
.Y(n_2921)
);

OAI22xp5_ASAP7_75t_L g2922 ( 
.A1(n_2905),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_2922)
);

INVx2_ASAP7_75t_L g2923 ( 
.A(n_2913),
.Y(n_2923)
);

AOI22xp5_ASAP7_75t_L g2924 ( 
.A1(n_2914),
.A2(n_1455),
.B1(n_1459),
.B2(n_1467),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2900),
.Y(n_2925)
);

AO22x2_ASAP7_75t_L g2926 ( 
.A1(n_2912),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_2926)
);

AOI22xp5_ASAP7_75t_L g2927 ( 
.A1(n_2902),
.A2(n_2910),
.B1(n_2898),
.B2(n_1467),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2903),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2903),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2920),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2926),
.Y(n_2931)
);

OAI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2919),
.A2(n_1459),
.B1(n_1467),
.B2(n_186),
.Y(n_2932)
);

AOI322xp5_ASAP7_75t_L g2933 ( 
.A1(n_2915),
.A2(n_181),
.A3(n_182),
.B1(n_188),
.B2(n_189),
.C1(n_192),
.C2(n_193),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_2923),
.Y(n_2934)
);

INVxp67_ASAP7_75t_L g2935 ( 
.A(n_2916),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2921),
.Y(n_2936)
);

AO22x2_ASAP7_75t_L g2937 ( 
.A1(n_2928),
.A2(n_182),
.B1(n_189),
.B2(n_193),
.Y(n_2937)
);

AOI22x1_ASAP7_75t_L g2938 ( 
.A1(n_2929),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_2938)
);

NAND2xp33_ASAP7_75t_L g2939 ( 
.A(n_2917),
.B(n_1459),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2922),
.Y(n_2940)
);

AOI221xp5_ASAP7_75t_L g2941 ( 
.A1(n_2925),
.A2(n_196),
.B1(n_904),
.B2(n_867),
.C(n_876),
.Y(n_2941)
);

NAND4xp75_ASAP7_75t_L g2942 ( 
.A(n_2930),
.B(n_2918),
.C(n_2927),
.D(n_2924),
.Y(n_2942)
);

XNOR2xp5_ASAP7_75t_L g2943 ( 
.A(n_2938),
.B(n_200),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2937),
.Y(n_2944)
);

OR2x2_ASAP7_75t_L g2945 ( 
.A(n_2931),
.B(n_201),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2937),
.Y(n_2946)
);

NOR2x1p5_ASAP7_75t_L g2947 ( 
.A(n_2936),
.B(n_904),
.Y(n_2947)
);

OAI22x1_ASAP7_75t_L g2948 ( 
.A1(n_2934),
.A2(n_2935),
.B1(n_2940),
.B2(n_2939),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2932),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2941),
.Y(n_2950)
);

NOR2x1_ASAP7_75t_L g2951 ( 
.A(n_2933),
.B(n_1195),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2930),
.Y(n_2952)
);

NOR2xp33_ASAP7_75t_L g2953 ( 
.A(n_2952),
.B(n_202),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2946),
.Y(n_2954)
);

AOI211xp5_ASAP7_75t_SL g2955 ( 
.A1(n_2950),
.A2(n_204),
.B(n_206),
.C(n_210),
.Y(n_2955)
);

INVxp67_ASAP7_75t_SL g2956 ( 
.A(n_2944),
.Y(n_2956)
);

AOI22xp5_ASAP7_75t_L g2957 ( 
.A1(n_2942),
.A2(n_1423),
.B1(n_1388),
.B2(n_1483),
.Y(n_2957)
);

A2O1A1Ixp33_ASAP7_75t_L g2958 ( 
.A1(n_2945),
.A2(n_904),
.B(n_1282),
.C(n_1313),
.Y(n_2958)
);

AOI22xp5_ASAP7_75t_L g2959 ( 
.A1(n_2948),
.A2(n_1423),
.B1(n_1388),
.B2(n_1483),
.Y(n_2959)
);

OAI21xp5_ASAP7_75t_SL g2960 ( 
.A1(n_2943),
.A2(n_904),
.B(n_1311),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2949),
.B(n_212),
.Y(n_2961)
);

AOI211xp5_ASAP7_75t_L g2962 ( 
.A1(n_2951),
.A2(n_219),
.B(n_222),
.C(n_230),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2947),
.Y(n_2963)
);

OAI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2952),
.A2(n_1331),
.B1(n_1304),
.B2(n_1307),
.Y(n_2964)
);

AND2x4_ASAP7_75t_L g2965 ( 
.A(n_2952),
.B(n_236),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2956),
.Y(n_2966)
);

OR2x2_ASAP7_75t_L g2967 ( 
.A(n_2954),
.B(n_240),
.Y(n_2967)
);

NOR2xp67_ASAP7_75t_L g2968 ( 
.A(n_2953),
.B(n_241),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2961),
.B(n_242),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2965),
.Y(n_2970)
);

HB1xp67_ASAP7_75t_L g2971 ( 
.A(n_2955),
.Y(n_2971)
);

NAND2xp33_ASAP7_75t_L g2972 ( 
.A(n_2963),
.B(n_1326),
.Y(n_2972)
);

INVx1_ASAP7_75t_SL g2973 ( 
.A(n_2957),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2960),
.Y(n_2974)
);

NAND3x1_ASAP7_75t_L g2975 ( 
.A(n_2959),
.B(n_244),
.C(n_245),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2964),
.Y(n_2976)
);

AOI221xp5_ASAP7_75t_L g2977 ( 
.A1(n_2966),
.A2(n_2962),
.B1(n_2958),
.B2(n_1326),
.C(n_874),
.Y(n_2977)
);

NAND4xp25_ASAP7_75t_L g2978 ( 
.A(n_2968),
.B(n_1324),
.C(n_1267),
.D(n_1264),
.Y(n_2978)
);

CKINVDCx5p33_ASAP7_75t_R g2979 ( 
.A(n_2970),
.Y(n_2979)
);

HB1xp67_ASAP7_75t_L g2980 ( 
.A(n_2967),
.Y(n_2980)
);

CKINVDCx16_ASAP7_75t_R g2981 ( 
.A(n_2971),
.Y(n_2981)
);

O2A1O1Ixp33_ASAP7_75t_L g2982 ( 
.A1(n_2972),
.A2(n_1230),
.B(n_1222),
.C(n_1201),
.Y(n_2982)
);

NOR2x1p5_ASAP7_75t_L g2983 ( 
.A(n_2969),
.B(n_250),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2975),
.B(n_254),
.Y(n_2984)
);

BUFx2_ASAP7_75t_L g2985 ( 
.A(n_2974),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2976),
.Y(n_2986)
);

AOI21xp5_ASAP7_75t_L g2987 ( 
.A1(n_2973),
.A2(n_930),
.B(n_1320),
.Y(n_2987)
);

XNOR2xp5_ASAP7_75t_SL g2988 ( 
.A(n_2971),
.B(n_255),
.Y(n_2988)
);

NOR3xp33_ASAP7_75t_SL g2989 ( 
.A(n_2966),
.B(n_257),
.C(n_260),
.Y(n_2989)
);

CKINVDCx5p33_ASAP7_75t_R g2990 ( 
.A(n_2966),
.Y(n_2990)
);

CKINVDCx5p33_ASAP7_75t_R g2991 ( 
.A(n_2966),
.Y(n_2991)
);

NOR4xp75_ASAP7_75t_L g2992 ( 
.A(n_2975),
.B(n_264),
.C(n_265),
.D(n_266),
.Y(n_2992)
);

CKINVDCx16_ASAP7_75t_R g2993 ( 
.A(n_2971),
.Y(n_2993)
);

OR2x2_ASAP7_75t_L g2994 ( 
.A(n_2967),
.B(n_268),
.Y(n_2994)
);

OAI21x1_ASAP7_75t_SL g2995 ( 
.A1(n_2966),
.A2(n_272),
.B(n_277),
.Y(n_2995)
);

NAND3xp33_ASAP7_75t_L g2996 ( 
.A(n_2966),
.B(n_876),
.C(n_869),
.Y(n_2996)
);

OAI211xp5_ASAP7_75t_SL g2997 ( 
.A1(n_2966),
.A2(n_278),
.B(n_280),
.C(n_285),
.Y(n_2997)
);

CKINVDCx5p33_ASAP7_75t_R g2998 ( 
.A(n_2966),
.Y(n_2998)
);

AOI22xp33_ASAP7_75t_L g2999 ( 
.A1(n_2966),
.A2(n_867),
.B1(n_869),
.B2(n_874),
.Y(n_2999)
);

INVx2_ASAP7_75t_L g3000 ( 
.A(n_2967),
.Y(n_3000)
);

OAI22xp5_ASAP7_75t_SL g3001 ( 
.A1(n_2966),
.A2(n_1282),
.B1(n_1284),
.B2(n_1285),
.Y(n_3001)
);

NOR2x1p5_ASAP7_75t_L g3002 ( 
.A(n_2966),
.B(n_287),
.Y(n_3002)
);

AO22x2_ASAP7_75t_L g3003 ( 
.A1(n_2986),
.A2(n_293),
.B1(n_295),
.B2(n_297),
.Y(n_3003)
);

NAND3xp33_ASAP7_75t_L g3004 ( 
.A(n_2979),
.B(n_867),
.C(n_869),
.Y(n_3004)
);

AOI21xp5_ASAP7_75t_L g3005 ( 
.A1(n_2984),
.A2(n_930),
.B(n_869),
.Y(n_3005)
);

OAI22xp5_ASAP7_75t_L g3006 ( 
.A1(n_2981),
.A2(n_1312),
.B1(n_1331),
.B2(n_1304),
.Y(n_3006)
);

XOR2x1_ASAP7_75t_L g3007 ( 
.A(n_3002),
.B(n_299),
.Y(n_3007)
);

OR2x2_ASAP7_75t_L g3008 ( 
.A(n_2994),
.B(n_300),
.Y(n_3008)
);

OAI22x1_ASAP7_75t_L g3009 ( 
.A1(n_2983),
.A2(n_305),
.B1(n_306),
.B2(n_307),
.Y(n_3009)
);

NOR2xp33_ASAP7_75t_L g3010 ( 
.A(n_2993),
.B(n_313),
.Y(n_3010)
);

OA22x2_ASAP7_75t_L g3011 ( 
.A1(n_2995),
.A2(n_1286),
.B1(n_1307),
.B2(n_1312),
.Y(n_3011)
);

NAND3xp33_ASAP7_75t_L g3012 ( 
.A(n_2990),
.B(n_867),
.C(n_869),
.Y(n_3012)
);

CKINVDCx20_ASAP7_75t_R g3013 ( 
.A(n_2991),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2989),
.B(n_315),
.Y(n_3014)
);

OAI21xp5_ASAP7_75t_L g3015 ( 
.A1(n_2988),
.A2(n_1320),
.B(n_1317),
.Y(n_3015)
);

AND2x2_ASAP7_75t_L g3016 ( 
.A(n_2980),
.B(n_323),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_3000),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2998),
.Y(n_3018)
);

BUFx2_ASAP7_75t_L g3019 ( 
.A(n_2985),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2992),
.Y(n_3020)
);

INVx2_ASAP7_75t_SL g3021 ( 
.A(n_2996),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_3001),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2978),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2977),
.Y(n_3024)
);

AOI221xp5_ASAP7_75t_L g3025 ( 
.A1(n_2987),
.A2(n_874),
.B1(n_876),
.B2(n_930),
.C(n_1132),
.Y(n_3025)
);

HB1xp67_ASAP7_75t_L g3026 ( 
.A(n_2999),
.Y(n_3026)
);

AOI21xp33_ASAP7_75t_SL g3027 ( 
.A1(n_2982),
.A2(n_329),
.B(n_331),
.Y(n_3027)
);

OA21x2_ASAP7_75t_L g3028 ( 
.A1(n_2997),
.A2(n_1325),
.B(n_1286),
.Y(n_3028)
);

AOI21xp5_ASAP7_75t_L g3029 ( 
.A1(n_2986),
.A2(n_930),
.B(n_874),
.Y(n_3029)
);

CKINVDCx20_ASAP7_75t_R g3030 ( 
.A(n_2979),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2988),
.Y(n_3031)
);

NOR3xp33_ASAP7_75t_L g3032 ( 
.A(n_2981),
.B(n_333),
.C(n_335),
.Y(n_3032)
);

NOR2xp67_ASAP7_75t_L g3033 ( 
.A(n_2984),
.B(n_341),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2983),
.B(n_343),
.Y(n_3034)
);

OAI211xp5_ASAP7_75t_L g3035 ( 
.A1(n_2984),
.A2(n_345),
.B(n_351),
.C(n_352),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2988),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2985),
.A2(n_874),
.B1(n_876),
.B2(n_1423),
.Y(n_3037)
);

OR5x1_ASAP7_75t_L g3038 ( 
.A(n_2978),
.B(n_353),
.C(n_357),
.D(n_359),
.E(n_360),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_3019),
.B(n_363),
.Y(n_3039)
);

NAND4xp75_ASAP7_75t_L g3040 ( 
.A(n_3010),
.B(n_365),
.C(n_366),
.D(n_371),
.Y(n_3040)
);

NOR2x2_ASAP7_75t_L g3041 ( 
.A(n_3017),
.B(n_3022),
.Y(n_3041)
);

NOR2x1_ASAP7_75t_L g3042 ( 
.A(n_3030),
.B(n_3016),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_3034),
.Y(n_3043)
);

NOR3x1_ASAP7_75t_L g3044 ( 
.A(n_3035),
.B(n_372),
.C(n_374),
.Y(n_3044)
);

NOR2xp67_ASAP7_75t_L g3045 ( 
.A(n_3009),
.B(n_375),
.Y(n_3045)
);

OAI221xp5_ASAP7_75t_L g3046 ( 
.A1(n_3014),
.A2(n_3018),
.B1(n_3015),
.B2(n_3020),
.C(n_3033),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_3007),
.Y(n_3047)
);

NAND3xp33_ASAP7_75t_L g3048 ( 
.A(n_3032),
.B(n_876),
.C(n_1113),
.Y(n_3048)
);

AOI22xp5_ASAP7_75t_L g3049 ( 
.A1(n_3013),
.A2(n_1320),
.B1(n_1317),
.B2(n_1325),
.Y(n_3049)
);

NOR3xp33_ASAP7_75t_L g3050 ( 
.A(n_3031),
.B(n_376),
.C(n_377),
.Y(n_3050)
);

AND3x4_ASAP7_75t_L g3051 ( 
.A(n_3038),
.B(n_378),
.C(n_379),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_3008),
.Y(n_3052)
);

OR2x6_ASAP7_75t_L g3053 ( 
.A(n_3036),
.B(n_3024),
.Y(n_3053)
);

NOR2x1p5_ASAP7_75t_L g3054 ( 
.A(n_3023),
.B(n_380),
.Y(n_3054)
);

XNOR2xp5_ASAP7_75t_L g3055 ( 
.A(n_3011),
.B(n_381),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_3026),
.Y(n_3056)
);

AND4x1_ASAP7_75t_L g3057 ( 
.A(n_3005),
.B(n_3004),
.C(n_3012),
.D(n_3029),
.Y(n_3057)
);

NAND3xp33_ASAP7_75t_SL g3058 ( 
.A(n_3025),
.B(n_382),
.C(n_388),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_3028),
.Y(n_3059)
);

NOR4xp25_ASAP7_75t_L g3060 ( 
.A(n_3021),
.B(n_391),
.C(n_392),
.D(n_393),
.Y(n_3060)
);

AO22x2_ASAP7_75t_L g3061 ( 
.A1(n_3006),
.A2(n_394),
.B1(n_398),
.B2(n_404),
.Y(n_3061)
);

INVx1_ASAP7_75t_L g3062 ( 
.A(n_3028),
.Y(n_3062)
);

OAI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_3027),
.A2(n_1313),
.B1(n_1329),
.B2(n_1224),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_3003),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_3003),
.Y(n_3065)
);

NAND2xp5_ASAP7_75t_L g3066 ( 
.A(n_3037),
.B(n_406),
.Y(n_3066)
);

AOI22xp5_ASAP7_75t_L g3067 ( 
.A1(n_3030),
.A2(n_1388),
.B1(n_1423),
.B2(n_1224),
.Y(n_3067)
);

OAI211xp5_ASAP7_75t_SL g3068 ( 
.A1(n_3018),
.A2(n_408),
.B(n_409),
.C(n_413),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_SL g3069 ( 
.A1(n_3030),
.A2(n_415),
.B1(n_1142),
.B2(n_1132),
.Y(n_3069)
);

NOR3xp33_ASAP7_75t_L g3070 ( 
.A(n_3019),
.B(n_969),
.C(n_980),
.Y(n_3070)
);

XNOR2x1_ASAP7_75t_L g3071 ( 
.A(n_3007),
.B(n_1092),
.Y(n_3071)
);

NAND3xp33_ASAP7_75t_SL g3072 ( 
.A(n_3030),
.B(n_1298),
.C(n_1293),
.Y(n_3072)
);

NAND4xp25_ASAP7_75t_L g3073 ( 
.A(n_3019),
.B(n_1225),
.C(n_1285),
.D(n_1284),
.Y(n_3073)
);

AO22x2_ASAP7_75t_L g3074 ( 
.A1(n_3017),
.A2(n_1225),
.B1(n_1285),
.B2(n_1284),
.Y(n_3074)
);

AO22x1_ASAP7_75t_L g3075 ( 
.A1(n_3010),
.A2(n_1142),
.B1(n_1092),
.B2(n_1113),
.Y(n_3075)
);

INVx2_ASAP7_75t_L g3076 ( 
.A(n_3008),
.Y(n_3076)
);

HB1xp67_ASAP7_75t_L g3077 ( 
.A(n_3054),
.Y(n_3077)
);

INVxp67_ASAP7_75t_L g3078 ( 
.A(n_3039),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_3055),
.Y(n_3079)
);

AOI221x1_ASAP7_75t_L g3080 ( 
.A1(n_3056),
.A2(n_1113),
.B1(n_1132),
.B2(n_1128),
.C(n_1092),
.Y(n_3080)
);

INVx3_ASAP7_75t_L g3081 ( 
.A(n_3064),
.Y(n_3081)
);

OAI22xp5_ASAP7_75t_L g3082 ( 
.A1(n_3051),
.A2(n_3045),
.B1(n_3047),
.B2(n_3042),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3065),
.Y(n_3083)
);

OAI21xp5_ASAP7_75t_L g3084 ( 
.A1(n_3052),
.A2(n_1195),
.B(n_1329),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_3076),
.B(n_1128),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_3071),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_3044),
.Y(n_3087)
);

A2O1A1Ixp33_ASAP7_75t_L g3088 ( 
.A1(n_3048),
.A2(n_1132),
.B(n_1091),
.C(n_1092),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_L g3089 ( 
.A(n_3043),
.B(n_1142),
.Y(n_3089)
);

AOI21xp33_ASAP7_75t_SL g3090 ( 
.A1(n_3050),
.A2(n_1269),
.B(n_1291),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_3040),
.Y(n_3091)
);

OAI22x1_ASAP7_75t_L g3092 ( 
.A1(n_3059),
.A2(n_1224),
.B1(n_1329),
.B2(n_1267),
.Y(n_3092)
);

AOI221xp5_ASAP7_75t_L g3093 ( 
.A1(n_3063),
.A2(n_1128),
.B1(n_1142),
.B2(n_1113),
.C(n_1267),
.Y(n_3093)
);

OAI22xp5_ASAP7_75t_L g3094 ( 
.A1(n_3053),
.A2(n_1253),
.B1(n_1195),
.B2(n_1264),
.Y(n_3094)
);

OAI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_3053),
.A2(n_1253),
.B1(n_1264),
.B2(n_1128),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_3062),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_3046),
.Y(n_3097)
);

NAND2xp33_ASAP7_75t_SL g3098 ( 
.A(n_3069),
.B(n_1253),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_3081),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_3077),
.Y(n_3100)
);

AND3x1_ASAP7_75t_L g3101 ( 
.A(n_3081),
.B(n_3060),
.C(n_3070),
.Y(n_3101)
);

CKINVDCx20_ASAP7_75t_R g3102 ( 
.A(n_3082),
.Y(n_3102)
);

CKINVDCx20_ASAP7_75t_R g3103 ( 
.A(n_3079),
.Y(n_3103)
);

CKINVDCx20_ASAP7_75t_R g3104 ( 
.A(n_3097),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_3083),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_L g3106 ( 
.A(n_3087),
.B(n_3075),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_3085),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_3091),
.Y(n_3108)
);

HB1xp67_ASAP7_75t_L g3109 ( 
.A(n_3096),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_3078),
.B(n_3057),
.Y(n_3110)
);

NAND2x1p5_ASAP7_75t_L g3111 ( 
.A(n_3086),
.B(n_3041),
.Y(n_3111)
);

AOI21x1_ASAP7_75t_L g3112 ( 
.A1(n_3109),
.A2(n_3105),
.B(n_3099),
.Y(n_3112)
);

AOI21x1_ASAP7_75t_L g3113 ( 
.A1(n_3100),
.A2(n_3089),
.B(n_3080),
.Y(n_3113)
);

XOR2xp5_ASAP7_75t_L g3114 ( 
.A(n_3104),
.B(n_3072),
.Y(n_3114)
);

OA22x2_ASAP7_75t_L g3115 ( 
.A1(n_3108),
.A2(n_3084),
.B1(n_3049),
.B2(n_3066),
.Y(n_3115)
);

OAI21xp5_ASAP7_75t_L g3116 ( 
.A1(n_3111),
.A2(n_3058),
.B(n_3094),
.Y(n_3116)
);

AOI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_3106),
.A2(n_3101),
.B(n_3102),
.Y(n_3117)
);

OAI22xp5_ASAP7_75t_L g3118 ( 
.A1(n_3103),
.A2(n_3090),
.B1(n_3061),
.B2(n_3088),
.Y(n_3118)
);

AOI21xp5_ASAP7_75t_L g3119 ( 
.A1(n_3110),
.A2(n_3098),
.B(n_3093),
.Y(n_3119)
);

OA21x2_ASAP7_75t_L g3120 ( 
.A1(n_3107),
.A2(n_3073),
.B(n_3092),
.Y(n_3120)
);

AOI222xp33_ASAP7_75t_SL g3121 ( 
.A1(n_3105),
.A2(n_3068),
.B1(n_3095),
.B2(n_3074),
.C1(n_3067),
.C2(n_1388),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3112),
.Y(n_3122)
);

OAI22xp5_ASAP7_75t_L g3123 ( 
.A1(n_3117),
.A2(n_3074),
.B1(n_875),
.B2(n_908),
.Y(n_3123)
);

INVx1_ASAP7_75t_L g3124 ( 
.A(n_3113),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_3115),
.Y(n_3125)
);

BUFx2_ASAP7_75t_L g3126 ( 
.A(n_3122),
.Y(n_3126)
);

OAI22xp5_ASAP7_75t_SL g3127 ( 
.A1(n_3125),
.A2(n_3114),
.B1(n_3116),
.B2(n_3120),
.Y(n_3127)
);

OAI221xp5_ASAP7_75t_R g3128 ( 
.A1(n_3127),
.A2(n_3124),
.B1(n_3118),
.B2(n_3121),
.C(n_3119),
.Y(n_3128)
);

INVx1_ASAP7_75t_SL g3129 ( 
.A(n_3128),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_3129),
.A2(n_3126),
.B(n_3123),
.Y(n_3130)
);

AOI211xp5_ASAP7_75t_L g3131 ( 
.A1(n_3130),
.A2(n_1149),
.B(n_948),
.C(n_969),
.Y(n_3131)
);


endmodule