module real_jpeg_5981_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_0),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g163 ( 
.A(n_0),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g174 ( 
.A(n_0),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_0),
.B(n_258),
.Y(n_257)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_2),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_2),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_2),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_2),
.B(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_2),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_2),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_2),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_2),
.B(n_347),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_4),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_4),
.B(n_32),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_4),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_4),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_4),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_4),
.B(n_242),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_5),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_5),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_5),
.B(n_117),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_5),
.B(n_90),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g428 ( 
.A(n_5),
.B(n_111),
.Y(n_428)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_7),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_8),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_8),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_8),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_8),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_8),
.B(n_460),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_9),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_9),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_9),
.B(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_9),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_9),
.B(n_372),
.Y(n_371)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_11),
.Y(n_70)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g441 ( 
.A(n_11),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_12),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_12),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_13),
.B(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_13),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_13),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_13),
.B(n_115),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_13),
.B(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_14),
.Y(n_122)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_14),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_14),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_15),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_15),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_15),
.B(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_15),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_15),
.B(n_366),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_448),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_419),
.B(n_447),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_303),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_219),
.B(n_262),
.C(n_263),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_189),
.B(n_218),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_22),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_156),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_23),
.B(n_156),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_106),
.C(n_140),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_24),
.B(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_71),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_25),
.B(n_72),
.C(n_87),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_47),
.C(n_61),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_26),
.B(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_41),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_35),
.B2(n_40),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_28),
.A2(n_29),
.B1(n_426),
.B2(n_427),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_28),
.A2(n_29),
.B1(n_73),
.B2(n_74),
.Y(n_469)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_29),
.B(n_35),
.C(n_41),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_29),
.B(n_198),
.C(n_428),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g74 ( 
.A(n_30),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_30),
.B(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_33),
.B(n_102),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_34),
.Y(n_359)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_38),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_38),
.Y(n_444)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_39),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_39),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_39),
.Y(n_301)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g315 ( 
.A(n_46),
.Y(n_315)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_46),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_47),
.A2(n_61),
.B1(n_62),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_47),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_55),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_48),
.A2(n_55),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_48),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_48),
.A2(n_198),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_48),
.A2(n_198),
.B1(n_428),
.B2(n_429),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_48),
.B(n_129),
.C(n_272),
.Y(n_432)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_52),
.B(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_54),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_55),
.Y(n_199)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_59),
.Y(n_211)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_60),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_63),
.A2(n_173),
.B1(n_174),
.B2(n_176),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_63),
.A2(n_67),
.B1(n_68),
.B2(n_176),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_63),
.B(n_174),
.C(n_177),
.Y(n_260)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_66),
.Y(n_369)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_70),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_87),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_74),
.B(n_80),
.C(n_85),
.Y(n_188)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_84),
.B2(n_85),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_81),
.B(n_129),
.Y(n_319)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_83),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_83),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_96),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_89),
.B(n_92),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_88),
.B(n_97),
.C(n_101),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_91),
.Y(n_186)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_106),
.B(n_140),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_124),
.C(n_126),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_107),
.A2(n_124),
.B1(n_125),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_114),
.C(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_109),
.B(n_377),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_109),
.B(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_111),
.Y(n_110)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_118),
.B1(n_119),
.B2(n_123),
.Y(n_113)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_118),
.A2(n_119),
.B1(n_240),
.B2(n_244),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_119),
.B(n_174),
.C(n_241),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_121),
.Y(n_119)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_121),
.Y(n_167)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_121),
.Y(n_318)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_122),
.Y(n_361)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_126),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.C(n_136),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_127),
.A2(n_128),
.B1(n_406),
.B2(n_407),
.Y(n_405)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_129),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_129),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_129),
.A2(n_228),
.B1(n_272),
.B2(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_129),
.B(n_231),
.C(n_238),
.Y(n_277)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_132),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_133),
.A2(n_134),
.B1(n_136),
.B2(n_137),
.Y(n_407)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_155),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_142),
.B(n_143),
.C(n_155),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_150),
.C(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_150),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_157),
.B(n_159),
.C(n_179),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_179),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_170),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_162),
.C(n_170),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_163),
.Y(n_226)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_166),
.B(n_168),
.C(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_174),
.B1(n_241),
.B2(n_243),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_173),
.A2(n_174),
.B1(n_311),
.B2(n_312),
.Y(n_348)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_174),
.B(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_177),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_177),
.A2(n_178),
.B1(n_443),
.B2(n_445),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_178),
.B(n_438),
.C(n_443),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_180),
.B(n_182),
.C(n_183),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_185),
.B(n_187),
.C(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_188),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_216),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_190),
.B(n_216),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_195),
.C(n_213),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_191),
.A2(n_192),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_195),
.B(n_213),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.C(n_212),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_196),
.B(n_401),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_200),
.B(n_212),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.C(n_207),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_201),
.A2(n_202),
.B1(n_207),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_206),
.B(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_207),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_208),
.B(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_208),
.B(n_380),
.Y(n_379)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_220),
.B(n_264),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_222),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_265),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_222),
.B(n_265),
.Y(n_418)
);

FAx1_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_245),
.CI(n_261),
.CON(n_222),
.SN(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_239),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_225),
.B(n_227),
.C(n_239),
.Y(n_290)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_238),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_235),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_235),
.A2(n_238),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_260),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_257),
.B2(n_259),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_257),
.C(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_257),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_257),
.A2(n_259),
.B1(n_299),
.B2(n_302),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_259),
.B(n_295),
.C(n_302),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_266),
.B(n_268),
.C(n_288),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_288),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_276),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_269),
.B(n_277),
.C(n_278),
.Y(n_446)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

INVx8_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_287),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_433)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_282),
.Y(n_285)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_289),
.B(n_293),
.C(n_294),
.Y(n_422)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

AO22x1_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_299),
.Y(n_302)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI31xp33_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_415),
.A3(n_416),
.B(n_418),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_409),
.B(n_414),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_396),
.B(n_408),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_349),
.B(n_395),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_335),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_308),
.B(n_335),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_321),
.C(n_332),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_310),
.B(n_316),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_310),
.B(n_317),
.C(n_319),
.Y(n_404)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_332),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.C(n_327),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_322),
.B(n_337),
.Y(n_336)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_325),
.A2(n_326),
.B1(n_327),
.B2(n_328),
.Y(n_337)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.C(n_348),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_392),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_338),
.A2(n_339),
.B1(n_348),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_345),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_340),
.A2(n_341),
.B1(n_345),
.B2(n_346),
.Y(n_362)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_389),
.B(n_394),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_374),
.B(n_388),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_363),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_363),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_362),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_360),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_360),
.C(n_362),
.Y(n_390)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx5_ASAP7_75t_SL g356 ( 
.A(n_357),
.Y(n_356)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx4_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_370),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_364),
.A2(n_365),
.B1(n_370),
.B2(n_371),
.Y(n_386)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx6_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx8_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_382),
.B(n_387),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_379),
.Y(n_375)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_383),
.B(n_386),
.Y(n_387)
);

INVx4_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_390),
.B(n_391),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_398),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_399),
.A2(n_400),
.B1(n_402),
.B2(n_403),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_399),
.B(n_404),
.C(n_405),
.Y(n_413)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_410),
.B(n_413),
.Y(n_414)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_411),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_421),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g472 ( 
.A(n_421),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_423),
.CI(n_434),
.CON(n_421),
.SN(n_421)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_423),
.C(n_434),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_425),
.B1(n_430),
.B2(n_431),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_424),
.B(n_432),
.C(n_433),
.Y(n_454)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_428),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_435),
.B(n_446),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_437),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_437),
.C(n_446),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_443),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_470),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_450),
.B(n_451),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_465),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_459),
.A2(n_462),
.B1(n_463),
.B2(n_464),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_459),
.Y(n_463)
);

INVx6_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_462),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);


endmodule