module fake_jpeg_5784_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_42),
.B(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_44),
.B(n_45),
.Y(n_82)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_46),
.B(n_54),
.Y(n_107)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_49),
.B(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_14),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_58),
.Y(n_88)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_56),
.A2(n_23),
.B1(n_37),
.B2(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_30),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_19),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_23),
.B1(n_35),
.B2(n_37),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_73),
.B1(n_18),
.B2(n_13),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_62),
.Y(n_125)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_72),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_29),
.B1(n_37),
.B2(n_15),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_79),
.B1(n_86),
.B2(n_105),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_68),
.B1(n_85),
.B2(n_100),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_29),
.B1(n_23),
.B2(n_31),
.Y(n_68)
);

AO22x1_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_31),
.B1(n_20),
.B2(n_34),
.Y(n_71)
);

OR2x4_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_12),
.Y(n_119)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_56),
.B1(n_27),
.B2(n_22),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_74),
.B(n_108),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_75),
.B(n_80),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_38),
.B1(n_22),
.B2(n_27),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_76),
.A2(n_84),
.B1(n_93),
.B2(n_103),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_36),
.B1(n_24),
.B2(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_83),
.B(n_94),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_46),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_39),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_36),
.B1(n_21),
.B2(n_20),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_45),
.Y(n_90)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_20),
.B1(n_30),
.B2(n_32),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_18),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_96),
.Y(n_133)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_57),
.A2(n_19),
.B1(n_18),
.B2(n_32),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_18),
.C(n_32),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_71),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_32),
.B1(n_30),
.B2(n_19),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_58),
.A2(n_18),
.B1(n_30),
.B2(n_3),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_109),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_111),
.B(n_112),
.Y(n_144)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_13),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_82),
.Y(n_163)
);

BUFx16f_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g116 ( 
.A1(n_64),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_74),
.B1(n_70),
.B2(n_99),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_69),
.A2(n_11),
.B1(n_9),
.B2(n_5),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_69),
.B1(n_87),
.B2(n_95),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_91),
.B(n_92),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_136),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_0),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_5),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_161),
.B(n_112),
.Y(n_184)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_146),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_133),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_151),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_95),
.B1(n_86),
.B2(n_99),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_145),
.A2(n_124),
.B1(n_116),
.B2(n_119),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_115),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_136),
.B(n_78),
.Y(n_149)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_150),
.Y(n_191)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_153),
.A2(n_147),
.B1(n_114),
.B2(n_109),
.Y(n_179)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_154),
.A2(n_155),
.B1(n_166),
.B2(n_171),
.Y(n_182)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_81),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_156),
.B(n_165),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g176 ( 
.A(n_157),
.Y(n_176)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_133),
.B(n_80),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_118),
.B(n_77),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_63),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_163),
.B(n_116),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_6),
.B(n_7),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_98),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_168),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_111),
.B(n_67),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_172),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_115),
.Y(n_170)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_111),
.B(n_67),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_123),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_173),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_125),
.B(n_106),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_178),
.A2(n_193),
.B1(n_208),
.B2(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_196),
.B1(n_202),
.B2(n_205),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_120),
.C(n_114),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_190),
.C(n_198),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_184),
.A2(n_173),
.B(n_155),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_150),
.B(n_120),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_187),
.B(n_204),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_167),
.B(n_185),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_135),
.C(n_117),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_147),
.A2(n_113),
.B1(n_127),
.B2(n_131),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_152),
.B(n_139),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_199),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_195),
.A2(n_164),
.B1(n_171),
.B2(n_141),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_144),
.A2(n_127),
.B1(n_131),
.B2(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_148),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_144),
.B(n_104),
.C(n_101),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_118),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_118),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_145),
.A2(n_77),
.B1(n_60),
.B2(n_65),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_143),
.B(n_6),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_165),
.A2(n_60),
.B1(n_65),
.B2(n_130),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_91),
.C(n_130),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_192),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_7),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_207),
.B(n_148),
.C(n_146),
.Y(n_227)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_161),
.B1(n_140),
.B2(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_209),
.B(n_211),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_185),
.A2(n_164),
.B(n_158),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_210),
.A2(n_229),
.B(n_230),
.Y(n_255)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_217),
.Y(n_237)
);

BUFx12f_ASAP7_75t_SL g213 ( 
.A(n_208),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_213),
.A2(n_218),
.B(n_221),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_219),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_202),
.B1(n_190),
.B2(n_178),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_179),
.A2(n_166),
.B1(n_154),
.B2(n_157),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_223),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_224),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_175),
.B(n_170),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_228),
.B(n_180),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_167),
.B(n_208),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_183),
.C(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_226),
.Y(n_266)
);

NAND3xp33_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_198),
.C(n_191),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g268 ( 
.A1(n_236),
.A2(n_210),
.B(n_217),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_213),
.Y(n_239)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_239),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_226),
.C(n_211),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_245),
.A2(n_216),
.B1(n_226),
.B2(n_233),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_251),
.Y(n_269)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_256),
.A2(n_209),
.B1(n_225),
.B2(n_221),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_257),
.A2(n_258),
.B1(n_248),
.B2(n_243),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_242),
.A2(n_216),
.B1(n_212),
.B2(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_263),
.B(n_247),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_242),
.A2(n_220),
.B1(n_230),
.B2(n_229),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_247),
.B1(n_256),
.B2(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_271),
.C(n_272),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_207),
.C(n_227),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_227),
.C(n_218),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_215),
.B(n_195),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_273),
.A2(n_255),
.B(n_237),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_283),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_276),
.B(n_278),
.Y(n_297)
);

AOI322xp5_ASAP7_75t_SL g276 ( 
.A1(n_268),
.A2(n_269),
.A3(n_272),
.B1(n_266),
.B2(n_271),
.C1(n_265),
.C2(n_261),
.Y(n_276)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_193),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_240),
.Y(n_281)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_281),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_287),
.B1(n_259),
.B2(n_264),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_245),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_260),
.B(n_228),
.Y(n_284)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_285),
.A2(n_238),
.B1(n_186),
.B2(n_241),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_240),
.B1(n_246),
.B2(n_252),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_290),
.A2(n_292),
.B(n_296),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_263),
.B1(n_270),
.B2(n_273),
.Y(n_291)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_291),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_279),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_258),
.C(n_231),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_294),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_253),
.B1(n_241),
.B2(n_195),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_298),
.A2(n_275),
.B1(n_201),
.B2(n_180),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_303),
.B(n_308),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_274),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_299),
.Y(n_312)
);

NOR2x1_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_281),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_203),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_203),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_307),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_201),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_293),
.C(n_286),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_312),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_296),
.B1(n_290),
.B2(n_291),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_302),
.B1(n_304),
.B2(n_306),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_311),
.B1(n_285),
.B2(n_300),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_313),
.A3(n_310),
.B1(n_283),
.B2(n_297),
.C1(n_316),
.C2(n_177),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_320),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_318),
.Y(n_323)
);


endmodule