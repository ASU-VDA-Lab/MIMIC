module real_jpeg_1214_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_84),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_84),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_1),
.A2(n_60),
.B1(n_64),
.B2(n_84),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_37),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_2),
.A2(n_37),
.B1(n_60),
.B2(n_64),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_44),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_44),
.B1(n_60),
.B2(n_64),
.Y(n_170)
);

BUFx4f_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_52),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_52),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_5),
.A2(n_52),
.B1(n_60),
.B2(n_64),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_41),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_6),
.B(n_53),
.Y(n_214)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_6),
.A2(n_7),
.B(n_25),
.C(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_6),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_6),
.B(n_30),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_6),
.B(n_60),
.C(n_63),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_227),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_6),
.B(n_113),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_6),
.B(n_58),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_7),
.A2(n_25),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_7),
.B(n_25),
.Y(n_29)
);

AO22x2_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_9),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_76),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_9),
.A2(n_60),
.B1(n_64),
.B2(n_76),
.Y(n_202)
);

BUFx16f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_123),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_123),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_12),
.A2(n_60),
.B1(n_64),
.B2(n_123),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_13),
.A2(n_41),
.B1(n_42),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_13),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_145),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_145),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_13),
.A2(n_60),
.B1(n_64),
.B2(n_145),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_15),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_177),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_177),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_15),
.A2(n_60),
.B1(n_64),
.B2(n_177),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_90),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_21),
.B(n_77),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_56),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_38),
.B1(n_54),
.B2(n_55),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_23),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_30),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_24),
.A2(n_30),
.B1(n_194),
.B2(n_211),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_25),
.A2(n_26),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

AOI32xp33_ASAP7_75t_L g197 ( 
.A1(n_25),
.A2(n_42),
.A3(n_47),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g199 ( 
.A(n_26),
.B(n_48),
.Y(n_199)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_30),
.B(n_174),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_31),
.A2(n_32),
.B1(n_62),
.B2(n_63),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_31),
.A2(n_34),
.B(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_32),
.B(n_272),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_36),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_45),
.B1(n_51),
.B2(n_53),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_40),
.A2(n_46),
.B1(n_74),
.B2(n_75),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_42),
.B1(n_47),
.B2(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

O2A1O1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_42),
.A2(n_74),
.B(n_227),
.C(n_236),
.Y(n_235)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_45),
.A2(n_53),
.B1(n_144),
.B2(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_74),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_46),
.A2(n_83),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_46),
.B(n_122),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_46),
.A2(n_120),
.B(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.C(n_73),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_69),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_82),
.C(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_65),
.B(n_67),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_58),
.A2(n_65),
.B1(n_118),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_58),
.A2(n_65),
.B1(n_139),
.B2(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_58),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_59),
.A2(n_68),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_59),
.A2(n_99),
.B1(n_100),
.B2(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_59),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_59),
.A2(n_243),
.B(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_59),
.A2(n_99),
.B1(n_220),
.B2(n_254),
.Y(n_265)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_60),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_60),
.B(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_65),
.A2(n_219),
.B(n_221),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_65),
.B(n_223),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_70),
.A2(n_72),
.B1(n_88),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_70),
.A2(n_72),
.B1(n_97),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_70),
.A2(n_193),
.B(n_195),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_70),
.A2(n_195),
.B(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_72),
.A2(n_141),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_72),
.A2(n_173),
.B(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_74),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_82),
.C(n_85),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_78),
.A2(n_82),
.B1(n_102),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_78),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_85),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AO21x1_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_153),
.B(n_324),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_148),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_124),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_93),
.B(n_124),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_101),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_96),
.B(n_98),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_101),
.C(n_105),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_99),
.A2(n_222),
.B(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_119),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_106),
.A2(n_107),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_108),
.A2(n_109),
.B1(n_119),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_113),
.B(n_114),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_110),
.A2(n_113),
.B1(n_136),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_110),
.A2(n_227),
.B(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_111),
.A2(n_112),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_111),
.A2(n_112),
.B1(n_202),
.B2(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_111),
.B(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_111),
.A2(n_258),
.B(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_111),
.A2(n_112),
.B1(n_258),
.B2(n_292),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_112),
.A2(n_217),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_112),
.B(n_231),
.Y(n_260)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_113),
.A2(n_230),
.B(n_287),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_116),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_119),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_131),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_140),
.C(n_142),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_133),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_134),
.A2(n_137),
.B1(n_138),
.B2(n_188),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_140),
.B(n_142),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_147),
.B(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_148),
.A2(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_149),
.B(n_152),
.Y(n_326)
);

AO21x1_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_178),
.B(n_323),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_155),
.B(n_158),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_164),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_162),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.C(n_175),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_166),
.B1(n_184),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_167),
.B(n_169),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_171),
.A2(n_172),
.B1(n_175),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_204),
.B(n_322),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_180),
.B(n_182),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_183),
.B(n_187),
.Y(n_307)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_189),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_196),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_190),
.B(n_192),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_196),
.B(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI31xp33_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_304),
.A3(n_314),
.B(n_319),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_248),
.B(n_303),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_232),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_207),
.B(n_232),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_218),
.C(n_224),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_208),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_213),
.C(n_216),
.Y(n_247)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_218),
.B(n_224),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_225),
.B(n_228),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_244),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_233),
.B(n_245),
.C(n_247),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_298),
.B(n_302),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_267),
.B(n_297),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_261),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_261),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_257),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_279),
.B(n_296),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_275),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_273),
.Y(n_294)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_290),
.B(n_295),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_285),
.B(n_289),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_288),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_287),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_293),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_301),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g319 ( 
.A1(n_305),
.A2(n_320),
.B(n_321),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_308),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_316),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_318),
.Y(n_320)
);


endmodule