module fake_jpeg_20178_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_30),
.B1(n_22),
.B2(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_9),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_36),
.Y(n_49)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_67),
.B1(n_39),
.B2(n_37),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_52),
.B(n_55),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_23),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_39),
.B(n_27),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_17),
.B1(n_31),
.B2(n_30),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_38),
.B1(n_35),
.B2(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_56),
.A2(n_32),
.B1(n_20),
.B2(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_19),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_38),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_40),
.A2(n_32),
.B1(n_20),
.B2(n_22),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

AND2x4_ASAP7_75t_SL g67 ( 
.A(n_41),
.B(n_31),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_41),
.B1(n_43),
.B2(n_35),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_68),
.A2(n_90),
.B1(n_57),
.B2(n_64),
.Y(n_102)
);

MAJx2_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_43),
.C(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_89),
.C(n_65),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_52),
.B(n_41),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_71),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_37),
.Y(n_75)
);

NAND2x1_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_37),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_80),
.B(n_84),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_77),
.B1(n_89),
.B2(n_73),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_91),
.B1(n_64),
.B2(n_38),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_37),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_34),
.B1(n_39),
.B2(n_23),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_65),
.B(n_50),
.C(n_61),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_88),
.A2(n_59),
.B(n_62),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_18),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_25),
.B1(n_24),
.B2(n_34),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_38),
.B1(n_34),
.B2(n_24),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_53),
.B(n_51),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_95),
.B(n_107),
.Y(n_128)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_79),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_112),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_54),
.B1(n_60),
.B2(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_110),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_102),
.A2(n_105),
.B1(n_115),
.B2(n_119),
.Y(n_136)
);

MAJx2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_55),
.C(n_51),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_63),
.B1(n_60),
.B2(n_58),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_64),
.B1(n_46),
.B2(n_48),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_106),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_0),
.B(n_1),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_64),
.B1(n_46),
.B2(n_47),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_74),
.A2(n_48),
.B1(n_47),
.B2(n_34),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_79),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_119),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_71),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_50),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_61),
.B1(n_34),
.B2(n_2),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_87),
.B(n_76),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_119),
.A2(n_76),
.B1(n_81),
.B2(n_74),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_122),
.A2(n_136),
.B1(n_139),
.B2(n_142),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_72),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_125),
.B(n_147),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_99),
.A2(n_76),
.B1(n_87),
.B2(n_72),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_129),
.A2(n_138),
.B1(n_145),
.B2(n_50),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_130),
.A2(n_117),
.B1(n_97),
.B2(n_112),
.Y(n_152)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_76),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_103),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_76),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_138),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_87),
.B1(n_82),
.B2(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_101),
.B1(n_105),
.B2(n_113),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_140),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_130),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_114),
.B1(n_95),
.B2(n_109),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_149),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_94),
.A2(n_121),
.B1(n_117),
.B2(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_150),
.B1(n_122),
.B2(n_136),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_104),
.A2(n_87),
.B1(n_86),
.B2(n_93),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_85),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_148),
.B(n_110),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_118),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_94),
.A2(n_24),
.B1(n_29),
.B2(n_28),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_162),
.B1(n_150),
.B2(n_130),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_126),
.A2(n_116),
.B(n_103),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_153),
.A2(n_172),
.B(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_157),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_111),
.C(n_100),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_159),
.C(n_171),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_115),
.C(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_163),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_12),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_123),
.B1(n_137),
.B2(n_129),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_124),
.B(n_24),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_124),
.Y(n_187)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_166),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_169),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_61),
.B1(n_10),
.B2(n_11),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_145),
.B1(n_128),
.B2(n_146),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_135),
.B(n_28),
.C(n_29),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_128),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_127),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_29),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_176),
.Y(n_182)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_175),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_29),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_28),
.B(n_25),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_25),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_154),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_142),
.B(n_0),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_191),
.B1(n_208),
.B2(n_155),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_187),
.B(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_188),
.A2(n_189),
.B1(n_201),
.B2(n_206),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_123),
.B1(n_130),
.B2(n_137),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_192),
.A2(n_174),
.B(n_176),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_193),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_146),
.C(n_149),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_197),
.C(n_158),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_143),
.C(n_9),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_8),
.B(n_15),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_172),
.B(n_163),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_16),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_154),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_168),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_15),
.B1(n_13),
.B2(n_10),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_13),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_202),
.Y(n_218)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_180),
.A2(n_13),
.B1(n_10),
.B2(n_9),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_223),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_214),
.B1(n_201),
.B2(n_199),
.Y(n_246)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_187),
.B(n_157),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_215),
.B(n_216),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_220),
.Y(n_234)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_192),
.Y(n_221)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_221),
.Y(n_251)
);

XNOR2x2_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_160),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_222),
.A2(n_224),
.B1(n_232),
.B2(n_170),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g224 ( 
.A(n_183),
.B(n_161),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_184),
.B(n_166),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_229),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_188),
.A2(n_173),
.B1(n_164),
.B2(n_161),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_205),
.B1(n_182),
.B2(n_151),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_171),
.C(n_173),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_233),
.C(n_191),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_190),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_185),
.B(n_181),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_205),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_231),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_184),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_178),
.C(n_159),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_245),
.C(n_248),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_240),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_222),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_239),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_197),
.C(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_246),
.A2(n_210),
.B1(n_151),
.B2(n_167),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_200),
.C(n_189),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_227),
.A2(n_198),
.B1(n_156),
.B2(n_175),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_250),
.B1(n_253),
.B2(n_206),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_218),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_182),
.C(n_156),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_217),
.C(n_230),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_217),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_268),
.C(n_234),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_244),
.A2(n_232),
.B(n_231),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_256),
.A2(n_267),
.B(n_3),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_224),
.B(n_214),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_210),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_215),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_242),
.B(n_223),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_235),
.B(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_245),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_237),
.B(n_243),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_277),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_236),
.B(n_254),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_276),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_234),
.B(n_247),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_167),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_278),
.A2(n_265),
.B1(n_269),
.B2(n_6),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_1),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_282),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_2),
.B(n_3),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_285),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_287),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_296),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_261),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_273),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_261),
.C(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_293),
.C(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_259),
.C(n_255),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_258),
.B(n_5),
.Y(n_296)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_283),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_282),
.B1(n_5),
.B2(n_6),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_291),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_304),
.A2(n_288),
.B(n_286),
.C(n_293),
.Y(n_306)
);

AOI21x1_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_311),
.B(n_312),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_304),
.B(n_286),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_310),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_4),
.Y(n_310)
);

AOI21x1_ASAP7_75t_L g316 ( 
.A1(n_313),
.A2(n_314),
.B(n_306),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_303),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_307),
.B(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_297),
.C(n_4),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_4),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_6),
.Y(n_320)
);


endmodule