module fake_jpeg_31318_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_39),
.B1(n_3),
.B2(n_4),
.Y(n_49)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_15),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_42),
.Y(n_45)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_34),
.B1(n_5),
.B2(n_4),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_5),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_37),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_59),
.B(n_55),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_21),
.C(n_6),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_14),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_13),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_66),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_47),
.C(n_46),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_70),
.C(n_63),
.Y(n_74)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_67),
.B(n_68),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_52),
.B1(n_16),
.B2(n_17),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_19),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_62),
.B(n_23),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_76),
.B(n_77),
.C(n_73),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_75),
.C(n_72),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_74),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_24),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_82),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_83)
);


endmodule