module fake_jpeg_27852_n_218 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_218);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx8_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_11),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_17),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g41 ( 
.A(n_25),
.B(n_21),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_25),
.C(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_47),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_11),
.B(n_27),
.C(n_15),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_41),
.B(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_49),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_12),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_52),
.A2(n_53),
.B1(n_59),
.B2(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_19),
.B1(n_23),
.B2(n_17),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_54),
.B(n_25),
.C(n_26),
.Y(n_70)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_43),
.B(n_35),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_54),
.A2(n_41),
.B1(n_42),
.B2(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_50),
.B1(n_45),
.B2(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_29),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_26),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_44),
.A2(n_42),
.B1(n_35),
.B2(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_72),
.A2(n_73),
.B1(n_55),
.B2(n_29),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_42),
.B1(n_35),
.B2(n_34),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_14),
.B(n_22),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_81),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_91),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_84),
.A2(n_68),
.B1(n_24),
.B2(n_28),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_11),
.B(n_2),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_66),
.B(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_87),
.B(n_94),
.Y(n_123)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_89),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_37),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_67),
.B(n_32),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_92),
.B(n_93),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_62),
.B(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_16),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_32),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_18),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_24),
.B1(n_28),
.B2(n_68),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_75),
.A3(n_76),
.B1(n_79),
.B2(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_102),
.A2(n_57),
.B1(n_37),
.B2(n_32),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_110),
.B1(n_119),
.B2(n_124),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_117),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_95),
.A2(n_99),
.B1(n_84),
.B2(n_97),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_126),
.B(n_83),
.Y(n_128)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_113),
.A2(n_82),
.B1(n_98),
.B2(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_121),
.B1(n_21),
.B2(n_13),
.Y(n_143)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2x1_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_14),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_148),
.B(n_149),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_129),
.B(n_135),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_81),
.B1(n_80),
.B2(n_82),
.Y(n_130)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_131),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_93),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_141),
.C(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_21),
.B1(n_22),
.B2(n_14),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_139),
.B(n_140),
.Y(n_155)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_103),
.B(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_109),
.A2(n_1),
.B(n_3),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_13),
.C(n_22),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_111),
.A2(n_14),
.B(n_13),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_1),
.B(n_3),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_105),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_162),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_130),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_120),
.C(n_121),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_158),
.C(n_163),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_145),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_163),
.A2(n_146),
.B1(n_127),
.B2(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_176),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_148),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_170),
.B(n_173),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_165),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_164),
.C(n_144),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_133),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_146),
.B1(n_118),
.B2(n_125),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_154),
.B1(n_149),
.B2(n_126),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_151),
.B(n_104),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_104),
.C(n_134),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_152),
.C(n_156),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_184),
.C(n_113),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_160),
.B(n_164),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_183),
.A2(n_6),
.B(n_9),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_119),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_188),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_115),
.C(n_124),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_187),
.B(n_102),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_175),
.Y(n_188)
);

AOI221xp5_ASAP7_75t_SL g190 ( 
.A1(n_186),
.A2(n_173),
.B1(n_169),
.B2(n_171),
.C(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_194),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_193),
.A2(n_197),
.B(n_7),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_178),
.Y(n_194)
);

BUFx24_ASAP7_75t_SL g195 ( 
.A(n_180),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_6),
.Y(n_201)
);

AOI21x1_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_187),
.B(n_180),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_189),
.C(n_5),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_203),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_194),
.A2(n_6),
.B1(n_9),
.B2(n_4),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_204),
.B1(n_5),
.B2(n_8),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_4),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_205),
.B(n_206),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_207),
.A2(n_199),
.B(n_10),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_200),
.A2(n_9),
.B(n_10),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_208),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_210),
.B(n_209),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_213),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_1),
.B(n_3),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_1),
.C(n_3),
.Y(n_218)
);


endmodule