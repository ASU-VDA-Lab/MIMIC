module fake_jpeg_18153_n_298 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_298);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_298;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_260;
wire n_112;
wire n_199;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_45),
.Y(n_60)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_43),
.B(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_55),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_39),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_29),
.B(n_1),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_44),
.A2(n_26),
.B1(n_17),
.B2(n_30),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_42),
.B1(n_43),
.B2(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_39),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_64),
.B(n_72),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_59),
.A2(n_17),
.B1(n_26),
.B2(n_30),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_67),
.A2(n_84),
.B1(n_95),
.B2(n_97),
.Y(n_130)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_69),
.A2(n_71),
.B1(n_79),
.B2(n_82),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_37),
.B1(n_43),
.B2(n_38),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_29),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_29),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_78),
.Y(n_132)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_81),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_52),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_38),
.B1(n_33),
.B2(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_27),
.B1(n_22),
.B2(n_18),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_86),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_18),
.B1(n_35),
.B2(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_87),
.Y(n_106)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_57),
.A2(n_36),
.B(n_35),
.C(n_34),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_94),
.B(n_0),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_48),
.B(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_54),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_92),
.A2(n_56),
.B1(n_19),
.B2(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_29),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_101),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_28),
.B1(n_24),
.B2(n_31),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AO22x1_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_32),
.B1(n_31),
.B2(n_23),
.Y(n_97)
);

OR2x2_ASAP7_75t_SL g99 ( 
.A(n_48),
.B(n_32),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_32),
.CI(n_21),
.CON(n_107),
.SN(n_107)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_104),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_56),
.A2(n_31),
.B1(n_23),
.B2(n_21),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_56),
.A2(n_23),
.B1(n_21),
.B2(n_19),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_97),
.B1(n_81),
.B2(n_83),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_107),
.B(n_122),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_32),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_111),
.B(n_125),
.C(n_107),
.Y(n_143)
);

AO21x2_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_99),
.B(n_97),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_124),
.B1(n_68),
.B2(n_86),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_134),
.B(n_1),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_70),
.B(n_7),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_127),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_85),
.B(n_7),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_80),
.B(n_9),
.C(n_14),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_64),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_72),
.B1(n_75),
.B2(n_94),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_142),
.B1(n_149),
.B2(n_157),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_146),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_120),
.B1(n_113),
.B2(n_134),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_147),
.B(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_101),
.B1(n_67),
.B2(n_90),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_118),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_132),
.A2(n_103),
.B(n_87),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_133),
.B(n_129),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_132),
.A2(n_98),
.B(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_121),
.B(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_151),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_108),
.A2(n_96),
.B1(n_100),
.B2(n_10),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_121),
.B(n_128),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_2),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_116),
.B(n_10),
.C(n_14),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_106),
.C(n_115),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_156),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_108),
.A2(n_9),
.B1(n_13),
.B2(n_4),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_113),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_158),
.B(n_159),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_3),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_11),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_161),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_109),
.B(n_11),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_113),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_107),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_123),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_192),
.Y(n_197)
);

BUFx4f_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_123),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_173),
.B(n_178),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_141),
.C(n_154),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_179),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_143),
.B(n_120),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_117),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_115),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_181),
.B(n_169),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_140),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_156),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_106),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_191),
.B1(n_138),
.B2(n_163),
.Y(n_205)
);

XOR2x1_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_131),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g207 ( 
.A1(n_187),
.A2(n_153),
.B(n_138),
.C(n_157),
.D(n_162),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_105),
.Y(n_188)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_188),
.Y(n_200)
);

INVx13_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

OAI22x1_ASAP7_75t_SL g191 ( 
.A1(n_142),
.A2(n_114),
.B1(n_105),
.B2(n_126),
.Y(n_191)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_13),
.B(n_6),
.C(n_10),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_201),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_195),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_190),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_164),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_210),
.Y(n_226)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_207),
.B(n_215),
.C(n_192),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_173),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_185),
.C(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_181),
.C(n_186),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_217),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_162),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_182),
.A2(n_150),
.B1(n_161),
.B2(n_137),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_168),
.B1(n_177),
.B2(n_171),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_182),
.A2(n_150),
.B1(n_155),
.B2(n_126),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_216),
.B1(n_166),
.B2(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_165),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_137),
.B(n_3),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_168),
.A2(n_152),
.B1(n_114),
.B2(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_220),
.B1(n_197),
.B2(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_166),
.B1(n_191),
.B2(n_175),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_223),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_167),
.C(n_183),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_233),
.C(n_216),
.Y(n_255)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_206),
.B(n_189),
.CI(n_177),
.CON(n_225),
.SN(n_225)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_228),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_174),
.C(n_172),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_204),
.C(n_212),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_230),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_184),
.B1(n_12),
.B2(n_16),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_197),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_184),
.C(n_16),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_198),
.Y(n_234)
);

BUFx24_ASAP7_75t_SL g254 ( 
.A(n_234),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_16),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_202),
.B(n_3),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_237),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_201),
.B1(n_228),
.B2(n_207),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_244),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_223),
.B(n_204),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_245),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_246),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_248),
.A2(n_195),
.B1(n_218),
.B2(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_229),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_251),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_221),
.B(n_215),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_235),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_233),
.C(n_225),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_238),
.C(n_254),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_248),
.A2(n_228),
.B1(n_199),
.B2(n_237),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_228),
.B1(n_239),
.B2(n_241),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_264),
.B1(n_244),
.B2(n_247),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_251),
.B1(n_255),
.B2(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_276),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_263),
.B(n_267),
.Y(n_271)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_271),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_272),
.B(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_247),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_266),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_258),
.C(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_275),
.C(n_271),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_268),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_262),
.B1(n_260),
.B2(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_282),
.Y(n_286)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_287),
.C(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_280),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_289),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_283),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_279),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_293),
.A2(n_294),
.B(n_292),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_296),
.B(n_286),
.Y(n_297)
);

XNOR2x2_ASAP7_75t_SL g298 ( 
.A(n_297),
.B(n_278),
.Y(n_298)
);


endmodule