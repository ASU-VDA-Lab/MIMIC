module fake_jpeg_30386_n_161 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_161);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_161;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx4f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_29),
.B(n_27),
.C(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_23),
.B(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_0),
.C(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_45),
.A2(n_48),
.B1(n_28),
.B2(n_27),
.Y(n_65)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_47),
.Y(n_58)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_30),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_19),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_64),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_23),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_60),
.B(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_24),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_36),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_62),
.A2(n_63),
.B1(n_51),
.B2(n_65),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g66 ( 
.A1(n_39),
.A2(n_18),
.B(n_20),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_42),
.B(n_24),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_SL g68 ( 
.A(n_43),
.Y(n_68)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_28),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_22),
.B1(n_18),
.B2(n_20),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_72),
.A2(n_45),
.B1(n_38),
.B2(n_28),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_76),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_46),
.B1(n_34),
.B2(n_5),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_81),
.Y(n_99)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_4),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_85),
.B1(n_51),
.B2(n_57),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_4),
.B1(n_6),
.B2(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx13_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_54),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_52),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_57),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_66),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_88),
.B(n_52),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_94),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_98),
.C(n_100),
.Y(n_114)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_60),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_49),
.B(n_55),
.C(n_64),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_65),
.B1(n_72),
.B2(n_69),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_107),
.B(n_91),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_71),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_92),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_82),
.A2(n_71),
.B(n_57),
.C(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_108),
.A2(n_110),
.B1(n_90),
.B2(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_100),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_113),
.B(n_115),
.Y(n_133)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_84),
.Y(n_117)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_117),
.A2(n_122),
.B(n_123),
.C(n_107),
.D(n_110),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_76),
.B1(n_73),
.B2(n_80),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_109),
.Y(n_119)
);

AO221x1_ASAP7_75t_L g126 ( 
.A1(n_119),
.A2(n_121),
.B1(n_101),
.B2(n_103),
.C(n_95),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_92),
.C(n_74),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_92),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_94),
.B(n_77),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_115),
.B(n_97),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_135),
.Y(n_142)
);

NAND3xp33_ASAP7_75t_L g131 ( 
.A(n_124),
.B(n_103),
.C(n_96),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_134),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_110),
.B1(n_96),
.B2(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_123),
.Y(n_134)
);

NOR4xp25_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_96),
.C(n_87),
.D(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_122),
.C(n_112),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_143),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_112),
.C(n_117),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_141),
.A2(n_129),
.B1(n_133),
.B2(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_148),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_133),
.B(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_149),
.Y(n_153)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_138),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_119),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_147),
.A2(n_137),
.B1(n_121),
.B2(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_151),
.B1(n_86),
.B2(n_93),
.Y(n_156)
);

OAI321xp33_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_142),
.A3(n_130),
.B1(n_143),
.B2(n_139),
.C(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_154),
.B(n_155),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_144),
.B(n_86),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_156),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_158),
.C(n_93),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_93),
.Y(n_161)
);


endmodule