module fake_jpeg_9219_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_5),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_22),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_18),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_25),
.Y(n_37)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_13),
.B1(n_17),
.B2(n_10),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_10),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_38),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_22),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_22),
.A2(n_13),
.B1(n_15),
.B2(n_12),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_19),
.B1(n_11),
.B2(n_20),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_41),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_37),
.Y(n_41)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_0),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_12),
.B1(n_15),
.B2(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_48),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_34),
.B1(n_32),
.B2(n_30),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_44),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_34),
.B1(n_30),
.B2(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_65),
.B(n_66),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_39),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_40),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_40),
.Y(n_67)
);

A2O1A1O1Ixp25_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_53),
.B(n_24),
.C(n_43),
.D(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_27),
.C(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_58),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_60),
.C(n_61),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_52),
.B1(n_46),
.B2(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_73),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_75),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_36),
.B(n_51),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_45),
.B1(n_25),
.B2(n_36),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_16),
.B(n_43),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_66),
.C(n_65),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_78),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_27),
.C(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

AO221x1_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_0),
.B1(n_11),
.B2(n_26),
.C(n_19),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_73),
.B(n_72),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_85),
.B(n_11),
.Y(n_87)
);

NOR2xp67_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_71),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_76),
.C(n_79),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_88),
.B(n_4),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_84),
.A2(n_2),
.B(n_3),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_11),
.Y(n_89)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_4),
.B(n_7),
.Y(n_91)
);

A2O1A1O1Ixp25_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_8),
.B(n_9),
.C(n_89),
.D(n_44),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_8),
.Y(n_93)
);


endmodule