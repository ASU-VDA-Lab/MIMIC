module real_jpeg_21608_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_300;
wire n_215;
wire n_221;
wire n_288;
wire n_292;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_164;
wire n_48;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_306;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_297;
wire n_55;
wire n_125;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_209;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_244;
wire n_179;
wire n_167;
wire n_216;
wire n_133;
wire n_213;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_0),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_32),
.B1(n_58),
.B2(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_0),
.A2(n_32),
.B1(n_50),
.B2(n_51),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_53),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_57),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_57),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_58),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_3),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_66),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_66),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_4),
.A2(n_58),
.B1(n_59),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_4),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_91),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_91),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_91),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_5),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_5),
.B(n_64),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_5),
.A2(n_47),
.B(n_50),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_154),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_5),
.A2(n_79),
.B1(n_80),
.B2(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_42),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_30),
.B(n_241),
.Y(n_240)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_7),
.Y(n_80)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_8),
.A2(n_30),
.B1(n_31),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_8),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_10),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_150),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_150),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_150),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_11),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_11),
.A2(n_30),
.B1(n_31),
.B2(n_156),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_156),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_156),
.Y(n_210)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_13),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_127),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_127),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_127),
.Y(n_244)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_14),
.A2(n_30),
.A3(n_39),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_62),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx3_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_92),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_70),
.C(n_76),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_23),
.A2(n_24),
.B1(n_70),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_24)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_43),
.C(n_54),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_30),
.B(n_62),
.Y(n_168)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_35),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_31),
.A2(n_63),
.B1(n_153),
.B2(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_31),
.B(n_154),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_33),
.A2(n_40),
.B1(n_42),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_33),
.A2(n_42),
.B1(n_73),
.B2(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_33),
.A2(n_42),
.B1(n_179),
.B2(n_181),
.Y(n_178)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_34),
.A2(n_37),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_34),
.A2(n_37),
.B1(n_151),
.B2(n_164),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_34),
.A2(n_37),
.B1(n_180),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_34),
.A2(n_37),
.B1(n_123),
.B2(n_164),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_35),
.B(n_38),
.Y(n_236)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_39),
.A2(n_48),
.B(n_154),
.C(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_43),
.A2(n_44),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_49),
.B1(n_52),
.B2(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_49),
.B1(n_75),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_45),
.A2(n_49),
.B1(n_87),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_45),
.A2(n_49),
.B1(n_120),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_45),
.A2(n_49),
.B1(n_142),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_45),
.A2(n_49),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_45),
.A2(n_49),
.B1(n_206),
.B2(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_45),
.A2(n_49),
.B1(n_226),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_45),
.A2(n_49),
.B1(n_146),
.B2(n_244),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_49),
.B(n_154),
.Y(n_211)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_51),
.B(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_54),
.A2(n_69),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_65),
.B2(n_67),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_56),
.A2(n_61),
.B1(n_64),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_58),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_62),
.Y(n_63)
);

HAxp5_ASAP7_75t_SL g153 ( 
.A(n_58),
.B(n_154),
.CON(n_153),
.SN(n_153)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_65),
.B1(n_67),
.B2(n_97),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_60),
.A2(n_67),
.B1(n_90),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_60),
.A2(n_67),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_60),
.A2(n_67),
.B1(n_126),
.B2(n_162),
.Y(n_282)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_61),
.A2(n_64),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_71),
.B(n_74),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_76),
.A2(n_77),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_88),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_88),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_78),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_78),
.A2(n_86),
.B1(n_112),
.B2(n_297),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_84),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_83),
.B1(n_84),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_79),
.A2(n_80),
.B1(n_118),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_79),
.A2(n_83),
.B1(n_140),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_79),
.A2(n_83),
.B1(n_170),
.B2(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_79),
.A2(n_81),
.B1(n_196),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_79),
.A2(n_83),
.B1(n_198),
.B2(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_79),
.A2(n_81),
.B1(n_185),
.B2(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_80),
.B(n_154),
.Y(n_214)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_82),
.A2(n_194),
.B1(n_195),
.B2(n_197),
.Y(n_193)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_86),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_88),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.Y(n_92)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_98),
.B1(n_99),
.B2(n_103),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_132),
.B(n_306),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_128),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_108),
.B(n_128),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_114),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_109),
.B(n_113),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_114),
.A2(n_115),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_121),
.C(n_124),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_116),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_117),
.B(n_119),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_121),
.A2(n_124),
.B1(n_125),
.B2(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_300),
.B(n_305),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_287),
.B(n_299),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_186),
.B(n_269),
.C(n_286),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_171),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_136),
.B(n_171),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_157),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_138),
.B(n_143),
.C(n_157),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_139),
.B(n_141),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_147),
.C(n_152),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_152),
.B(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_166),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_165),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_159),
.B(n_165),
.C(n_166),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_163),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_169),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_176),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_183),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_182),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_268),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_263),
.B(n_267),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_249),
.B(n_262),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_230),
.B(n_248),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_218),
.B(n_229),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_207),
.B(n_217),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_199),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_212),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_211),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_211),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_220),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_227),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_225),
.C(n_227),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_232),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_238),
.B1(n_246),
.B2(n_247),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_233),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_235),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_259),
.C(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_259),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_264),
.B(n_265),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_271),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_285),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_278),
.C(n_285),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_281),
.C(n_284),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_288),
.B(n_289),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_298),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_295),
.B2(n_296),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_296),
.C(n_298),
.Y(n_301)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);


endmodule