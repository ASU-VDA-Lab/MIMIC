module fake_jpeg_349_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_54),
.Y(n_68)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

CKINVDCx6p67_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_61),
.Y(n_73)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_45),
.B1(n_48),
.B2(n_43),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_49),
.B1(n_40),
.B2(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_53),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_67),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_69),
.B(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_51),
.Y(n_70)
);

BUFx2_ASAP7_75t_SL g74 ( 
.A(n_72),
.Y(n_74)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_43),
.B1(n_55),
.B2(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_71),
.A2(n_50),
.B1(n_49),
.B2(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_78),
.B1(n_5),
.B2(n_6),
.Y(n_101)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_64),
.B(n_72),
.C(n_50),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_54),
.C(n_3),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_86),
.B(n_26),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_15),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_87),
.B(n_0),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_73),
.B(n_72),
.C(n_2),
.Y(n_88)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_6),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_1),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_101),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_17),
.B1(n_35),
.B2(n_32),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_97),
.B(n_103),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_99),
.B1(n_8),
.B2(n_10),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_84),
.B1(n_81),
.B2(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_38),
.C(n_28),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_119),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_108),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_114),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_23),
.B(n_24),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_10),
.B(n_11),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_96),
.B(n_12),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_99),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_19),
.C(n_25),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_120),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_96),
.B1(n_102),
.B2(n_13),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_125),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_27),
.B(n_12),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_104),
.A2(n_11),
.B(n_14),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_129),
.A2(n_115),
.B1(n_118),
.B2(n_106),
.C(n_110),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_126),
.B(n_124),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_124),
.C(n_105),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_136),
.B(n_123),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_112),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_132),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_140),
.A2(n_138),
.B(n_111),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_118),
.C(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_134),
.C(n_108),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_14),
.Y(n_145)
);


endmodule