module fake_aes_8485_n_835 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_835);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_835;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_807;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_786;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_721;
wire n_438;
wire n_656;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_198;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g182 ( .A(n_128), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_53), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_175), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_31), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_13), .Y(n_186) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_84), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_53), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_81), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_80), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_67), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_16), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_72), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_25), .Y(n_195) );
INVxp67_ASAP7_75t_SL g196 ( .A(n_159), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_174), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_32), .Y(n_198) );
INVxp33_ASAP7_75t_L g199 ( .A(n_42), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_50), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_47), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_61), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_29), .Y(n_203) );
INVx1_ASAP7_75t_SL g204 ( .A(n_34), .Y(n_204) );
INVxp67_ASAP7_75t_SL g205 ( .A(n_177), .Y(n_205) );
NOR2xp67_ASAP7_75t_L g206 ( .A(n_152), .B(n_90), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_7), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_44), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_2), .Y(n_209) );
INVxp33_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
INVxp33_ASAP7_75t_SL g211 ( .A(n_12), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_149), .Y(n_212) );
CKINVDCx5p33_ASAP7_75t_R g213 ( .A(n_143), .Y(n_213) );
NOR2xp67_ASAP7_75t_L g214 ( .A(n_170), .B(n_167), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_145), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_82), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_19), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_157), .Y(n_218) );
CKINVDCx14_ASAP7_75t_R g219 ( .A(n_78), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_30), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_39), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_16), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_104), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_71), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_69), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_14), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_38), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_94), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_54), .Y(n_230) );
CKINVDCx14_ASAP7_75t_R g231 ( .A(n_8), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g232 ( .A(n_135), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_49), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_110), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_29), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_86), .Y(n_236) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_27), .Y(n_237) );
BUFx8_ASAP7_75t_SL g238 ( .A(n_9), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_178), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_85), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_98), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
INVxp33_ASAP7_75t_SL g243 ( .A(n_107), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_148), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_142), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_150), .Y(n_246) );
INVxp33_ASAP7_75t_L g247 ( .A(n_140), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_100), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_63), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_114), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_124), .Y(n_251) );
INVxp33_ASAP7_75t_SL g252 ( .A(n_31), .Y(n_252) );
BUFx5_ASAP7_75t_L g253 ( .A(n_127), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_180), .B(n_154), .Y(n_254) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_56), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_46), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_138), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_51), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_47), .Y(n_259) );
INVx2_ASAP7_75t_L g260 ( .A(n_64), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_77), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_36), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_144), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_164), .Y(n_264) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_65), .Y(n_265) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_48), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_66), .Y(n_267) );
INVxp67_ASAP7_75t_SL g268 ( .A(n_48), .Y(n_268) );
INVxp67_ASAP7_75t_SL g269 ( .A(n_173), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_21), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_83), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_131), .Y(n_272) );
INVx1_ASAP7_75t_SL g273 ( .A(n_27), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_253), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_231), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_186), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_255), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g279 ( .A1(n_211), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_279) );
OAI22xp33_ASAP7_75t_SL g280 ( .A1(n_211), .A2(n_0), .B1(n_3), .B2(n_4), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_253), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_187), .Y(n_283) );
INVx6_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_187), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_186), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_187), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_198), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_198), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_199), .B(n_4), .Y(n_290) );
AND2x2_ASAP7_75t_SL g291 ( .A(n_271), .B(n_181), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_221), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_187), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_227), .B(n_5), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_242), .Y(n_296) );
INVx5_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_256), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_224), .B(n_6), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_256), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_265), .B(n_6), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_262), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_262), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_182), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_278), .B(n_210), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_284), .Y(n_306) );
AND2x2_ASAP7_75t_SL g307 ( .A(n_291), .B(n_189), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_295), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_276), .B(n_247), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_274), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_276), .B(n_266), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_295), .A2(n_185), .B1(n_188), .B2(n_183), .Y(n_313) );
AND2x4_ASAP7_75t_L g314 ( .A(n_295), .B(n_200), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_290), .B(n_201), .Y(n_315) );
NAND2xp5_ASAP7_75t_SL g316 ( .A(n_304), .B(n_247), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_283), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_304), .B(n_202), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_219), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_274), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_301), .Y(n_322) );
INVxp67_ASAP7_75t_SL g323 ( .A(n_301), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_284), .B(n_192), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_284), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_279), .A2(n_252), .B1(n_243), .B2(n_233), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_275), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_297), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_292), .B(n_203), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_275), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_286), .B(n_191), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_283), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_275), .B(n_237), .C(n_233), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_286), .B(n_207), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_292), .B(n_237), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_292), .B(n_259), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
BUFx4f_ASAP7_75t_L g339 ( .A(n_289), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_281), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_289), .B(n_259), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_281), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_305), .B(n_243), .Y(n_343) );
AND2x4_ASAP7_75t_L g344 ( .A(n_320), .B(n_315), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_309), .B(n_213), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_335), .Y(n_347) );
INVx2_ASAP7_75t_SL g348 ( .A(n_320), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_327), .Y(n_350) );
NAND2xp5_ASAP7_75t_SL g351 ( .A(n_322), .B(n_213), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_315), .A2(n_280), .B1(n_282), .B2(n_281), .Y(n_352) );
AO21x1_ASAP7_75t_L g353 ( .A1(n_308), .A2(n_282), .B(n_314), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_311), .B(n_216), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_316), .B(n_216), .Y(n_355) );
INVx4_ASAP7_75t_L g356 ( .A(n_306), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_314), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_319), .B(n_282), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_326), .A2(n_268), .B1(n_273), .B2(n_235), .C(n_204), .Y(n_360) );
AND3x1_ASAP7_75t_L g361 ( .A(n_313), .B(n_238), .C(n_220), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_331), .B(n_236), .Y(n_362) );
AND2x6_ASAP7_75t_SL g363 ( .A(n_329), .B(n_217), .Y(n_363) );
OR2x6_ASAP7_75t_L g364 ( .A(n_336), .B(n_223), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_337), .B(n_293), .Y(n_366) );
INVx5_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_339), .B(n_239), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_333), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_325), .B(n_239), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_330), .B(n_240), .Y(n_372) );
INVx3_ASAP7_75t_L g373 ( .A(n_327), .Y(n_373) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_306), .Y(n_374) );
INVx5_ASAP7_75t_L g375 ( .A(n_328), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_340), .B(n_241), .Y(n_376) );
AND2x4_ASAP7_75t_L g377 ( .A(n_306), .B(n_293), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_340), .B(n_241), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_342), .Y(n_379) );
INVx5_ASAP7_75t_L g380 ( .A(n_328), .Y(n_380) );
BUFx6f_ASAP7_75t_SL g381 ( .A(n_317), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_312), .B(n_249), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_310), .B(n_249), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_321), .B(n_257), .Y(n_384) );
NOR3xp33_ASAP7_75t_SL g385 ( .A(n_321), .B(n_209), .C(n_257), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_317), .B(n_184), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_317), .B(n_196), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_317), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_332), .B(n_195), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_332), .B(n_205), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_332), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_332), .B(n_298), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_332), .Y(n_393) );
AND2x4_ASAP7_75t_L g394 ( .A(n_323), .B(n_300), .Y(n_394) );
INVx3_ASAP7_75t_L g395 ( .A(n_334), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_341), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_323), .Y(n_397) );
BUFx2_ASAP7_75t_SL g398 ( .A(n_323), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_323), .B(n_269), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_318), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_318), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_323), .B(n_232), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_398), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_396), .B(n_208), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_397), .B(n_228), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_402), .A2(n_193), .B(n_190), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_374), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_348), .B(n_230), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_395), .B(n_302), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_358), .A2(n_197), .B(n_194), .Y(n_410) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_SL g412 ( .A1(n_343), .A2(n_254), .B(n_303), .C(n_302), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_352), .A2(n_270), .B1(n_258), .B2(n_303), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_394), .Y(n_415) );
INVx3_ASAP7_75t_L g416 ( .A(n_356), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_396), .B(n_212), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
AND2x4_ASAP7_75t_L g419 ( .A(n_364), .B(n_222), .Y(n_419) );
BUFx4f_ASAP7_75t_SL g420 ( .A(n_389), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_377), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_369), .A2(n_244), .B(n_234), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_353), .A2(n_246), .B(n_245), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_379), .Y(n_424) );
A2O1A1Ixp33_ASAP7_75t_L g425 ( .A1(n_349), .A2(n_250), .B(n_251), .C(n_248), .Y(n_425) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_367), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_357), .B(n_359), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_354), .Y(n_428) );
BUFx3_ASAP7_75t_L g429 ( .A(n_367), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_399), .B(n_261), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_366), .B(n_264), .Y(n_431) );
INVx1_ASAP7_75t_SL g432 ( .A(n_377), .Y(n_432) );
AOI221x1_ASAP7_75t_L g433 ( .A1(n_387), .A2(n_260), .B1(n_226), .B2(n_229), .C(n_225), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_346), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_347), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
OAI21x1_ASAP7_75t_L g437 ( .A1(n_390), .A2(n_226), .B(n_215), .Y(n_437) );
INVx1_ASAP7_75t_SL g438 ( .A(n_372), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_350), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_390), .A2(n_214), .B(n_206), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_366), .A2(n_272), .B1(n_218), .B2(n_260), .Y(n_442) );
OR2x6_ASAP7_75t_L g443 ( .A(n_351), .B(n_229), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_375), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_345), .B(n_8), .Y(n_445) );
INVx5_ASAP7_75t_L g446 ( .A(n_375), .Y(n_446) );
INVx4_ASAP7_75t_L g447 ( .A(n_375), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_376), .B(n_263), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_376), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_378), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_375), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_365), .B(n_9), .Y(n_452) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_383), .A2(n_267), .B(n_263), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_370), .B(n_267), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_392), .A2(n_383), .B(n_384), .C(n_355), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_380), .Y(n_456) );
AND3x1_ASAP7_75t_SL g457 ( .A(n_360), .B(n_10), .C(n_11), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_380), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_361), .B(n_10), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_371), .B(n_253), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_382), .Y(n_461) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_388), .Y(n_462) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_362), .A2(n_242), .B1(n_297), .B2(n_294), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_385), .B(n_297), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_368), .A2(n_297), .B(n_285), .Y(n_465) );
BUFx3_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_391), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_381), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_363), .A2(n_296), .B(n_294), .C(n_287), .Y(n_469) );
BUFx3_ASAP7_75t_L g470 ( .A(n_381), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_398), .A2(n_297), .B1(n_296), .B2(n_294), .Y(n_471) );
NOR2xp33_ASAP7_75t_SL g472 ( .A(n_398), .B(n_283), .Y(n_472) );
O2A1O1Ixp5_ASAP7_75t_SL g473 ( .A1(n_386), .A2(n_296), .B(n_294), .C(n_287), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_374), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_367), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_352), .A2(n_296), .B1(n_294), .B2(n_287), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_402), .A2(n_285), .B(n_283), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_398), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_398), .A2(n_296), .B1(n_287), .B2(n_285), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_428), .A2(n_287), .B1(n_285), .B2(n_17), .C(n_18), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_404), .B(n_15), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_470), .Y(n_482) );
NAND2x1p5_ASAP7_75t_L g483 ( .A(n_403), .B(n_285), .Y(n_483) );
OAI21x1_ASAP7_75t_L g484 ( .A1(n_437), .A2(n_287), .B(n_285), .Y(n_484) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_478), .B(n_17), .Y(n_485) );
OAI21x1_ASAP7_75t_L g486 ( .A1(n_473), .A2(n_68), .B(n_62), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
AO32x2_ASAP7_75t_L g488 ( .A1(n_476), .A2(n_18), .A3(n_19), .B1(n_20), .B2(n_21), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
OAI21x1_ASAP7_75t_L g490 ( .A1(n_477), .A2(n_73), .B(n_70), .Y(n_490) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_423), .A2(n_75), .B(n_74), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_436), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_439), .Y(n_493) );
AO21x2_ASAP7_75t_L g494 ( .A1(n_423), .A2(n_79), .B(n_76), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_434), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_415), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_405), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_414), .B(n_22), .Y(n_498) );
OAI21x1_ASAP7_75t_L g499 ( .A1(n_465), .A2(n_88), .B(n_87), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_438), .B(n_23), .Y(n_500) );
OAI21x1_ASAP7_75t_L g501 ( .A1(n_453), .A2(n_91), .B(n_89), .Y(n_501) );
AO31x2_ASAP7_75t_L g502 ( .A1(n_433), .A2(n_24), .A3(n_25), .B(n_26), .Y(n_502) );
OA21x2_ASAP7_75t_L g503 ( .A1(n_455), .A2(n_93), .B(n_92), .Y(n_503) );
AOI21x1_ASAP7_75t_L g504 ( .A1(n_460), .A2(n_96), .B(n_95), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_440), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_406), .A2(n_121), .B(n_179), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_420), .B(n_28), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_449), .A2(n_30), .B(n_32), .C(n_33), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_447), .Y(n_510) );
AOI21x1_ASAP7_75t_L g511 ( .A1(n_448), .A2(n_122), .B(n_176), .Y(n_511) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_409), .A2(n_123), .B(n_172), .Y(n_512) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_469), .A2(n_120), .B(n_169), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_450), .B(n_35), .Y(n_514) );
AND2x4_ASAP7_75t_L g515 ( .A(n_446), .B(n_37), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_408), .Y(n_516) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_409), .A2(n_119), .B(n_168), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g518 ( .A(n_446), .B(n_37), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_417), .B(n_38), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_426), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_464), .A2(n_125), .B(n_166), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_438), .B(n_40), .Y(n_522) );
AO31x2_ASAP7_75t_L g523 ( .A1(n_413), .A2(n_40), .A3(n_41), .B(n_42), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_411), .Y(n_524) );
INVx2_ASAP7_75t_SL g525 ( .A(n_446), .Y(n_525) );
OAI21x1_ASAP7_75t_L g526 ( .A1(n_479), .A2(n_126), .B(n_165), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_417), .B(n_43), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_411), .Y(n_528) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_421), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_427), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_475), .B(n_44), .Y(n_531) );
BUFx3_ASAP7_75t_L g532 ( .A(n_426), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_412), .A2(n_129), .B(n_163), .C(n_162), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_427), .Y(n_534) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_410), .A2(n_117), .B(n_161), .Y(n_535) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_472), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_462), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_431), .B(n_45), .Y(n_538) );
OAI21x1_ASAP7_75t_L g539 ( .A1(n_471), .A2(n_118), .B(n_160), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_411), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_422), .A2(n_130), .B(n_156), .Y(n_541) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_407), .A2(n_116), .B(n_153), .Y(n_542) );
INVx2_ASAP7_75t_SL g543 ( .A(n_462), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_462), .Y(n_544) );
OR2x6_ASAP7_75t_L g545 ( .A(n_475), .B(n_50), .Y(n_545) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_418), .A2(n_115), .B(n_151), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_474), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_452), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_474), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_452), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_432), .B(n_52), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_454), .Y(n_552) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_426), .B(n_55), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_451), .Y(n_554) );
OR2x6_ASAP7_75t_L g555 ( .A(n_468), .B(n_57), .Y(n_555) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_441), .A2(n_133), .B(n_147), .Y(n_556) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_425), .A2(n_132), .B(n_146), .Y(n_557) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_451), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_430), .A2(n_58), .B(n_59), .C(n_60), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_419), .B(n_58), .Y(n_560) );
INVx2_ASAP7_75t_SL g561 ( .A(n_451), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g562 ( .A(n_472), .B(n_134), .Y(n_562) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_416), .A2(n_97), .B(n_99), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_430), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_564) );
OAI21x1_ASAP7_75t_L g565 ( .A1(n_416), .A2(n_105), .B(n_106), .Y(n_565) );
OAI21x1_ASAP7_75t_L g566 ( .A1(n_463), .A2(n_108), .B(n_109), .Y(n_566) );
OAI21x1_ASAP7_75t_L g567 ( .A1(n_442), .A2(n_111), .B(n_112), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_474), .Y(n_568) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_429), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_461), .B(n_113), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_497), .B(n_419), .Y(n_571) );
INVx4_ASAP7_75t_L g572 ( .A(n_545), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_492), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_493), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_514), .A2(n_457), .B1(n_459), .B2(n_445), .Y(n_575) );
AOI21xp5_ASAP7_75t_SL g576 ( .A1(n_536), .A2(n_466), .B(n_443), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_545), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_545), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_481), .B(n_458), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_533), .A2(n_441), .B(n_467), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_552), .A2(n_444), .B(n_456), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_485), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_544), .Y(n_583) );
INVx3_ASAP7_75t_L g584 ( .A(n_532), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_489), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_544), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g587 ( .A1(n_508), .A2(n_137), .B(n_139), .C(n_141), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_496), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_530), .B(n_534), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_489), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_519), .A2(n_560), .B1(n_555), .B2(n_529), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_503), .A2(n_562), .B(n_541), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_537), .B(n_543), .Y(n_594) );
INVx3_ASAP7_75t_L g595 ( .A(n_532), .Y(n_595) );
AOI21xp33_ASAP7_75t_L g596 ( .A1(n_538), .A2(n_527), .B(n_516), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_531), .A2(n_548), .B1(n_550), .B2(n_498), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_518), .B(n_515), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_531), .A2(n_529), .B1(n_500), .B2(n_522), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_480), .B(n_509), .C(n_559), .Y(n_600) );
AO31x2_ASAP7_75t_L g601 ( .A1(n_509), .A2(n_559), .A3(n_564), .B(n_507), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_506), .Y(n_602) );
BUFx3_ASAP7_75t_L g603 ( .A(n_482), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_505), .B(n_510), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_531), .A2(n_570), .B1(n_515), .B2(n_551), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_553), .Y(n_606) );
INVx4_ASAP7_75t_L g607 ( .A(n_515), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_505), .B(n_510), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_525), .B(n_554), .Y(n_609) );
OR2x6_ASAP7_75t_L g610 ( .A(n_520), .B(n_558), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_561), .B(n_520), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g612 ( .A1(n_483), .A2(n_554), .B1(n_569), .B2(n_558), .Y(n_612) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_483), .A2(n_569), .B1(n_520), .B2(n_558), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_569), .A2(n_494), .B1(n_491), .B2(n_557), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_523), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_523), .B(n_488), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_524), .A2(n_540), .B1(n_568), .B2(n_528), .Y(n_617) );
INVx5_ASAP7_75t_L g618 ( .A(n_528), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_523), .B(n_540), .Y(n_619) );
OA21x2_ASAP7_75t_L g620 ( .A1(n_566), .A2(n_535), .B(n_567), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_547), .A2(n_549), .B1(n_556), .B2(n_513), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
INVx3_ASAP7_75t_L g623 ( .A(n_547), .Y(n_623) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_502), .Y(n_624) );
OAI22xp33_ASAP7_75t_SL g625 ( .A1(n_488), .A2(n_504), .B1(n_502), .B2(n_511), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_488), .A2(n_512), .B1(n_517), .B2(n_563), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_521), .B(n_539), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_488), .B(n_565), .Y(n_628) );
AND2x4_ASAP7_75t_L g629 ( .A(n_521), .B(n_526), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g630 ( .A1(n_501), .A2(n_490), .B1(n_499), .B2(n_542), .C(n_546), .Y(n_630) );
AND2x4_ASAP7_75t_L g631 ( .A(n_497), .B(n_403), .Y(n_631) );
AND2x2_ASAP7_75t_SL g632 ( .A(n_514), .B(n_307), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_487), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_497), .B(n_396), .Y(n_634) );
AND2x4_ASAP7_75t_L g635 ( .A(n_497), .B(n_403), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_487), .Y(n_636) );
OA21x2_ASAP7_75t_L g637 ( .A1(n_484), .A2(n_486), .B(n_566), .Y(n_637) );
AO31x2_ASAP7_75t_L g638 ( .A1(n_509), .A2(n_433), .A3(n_476), .B(n_455), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_591), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_634), .B(n_590), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_585), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_598), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_615), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_632), .B(n_602), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_573), .B(n_574), .Y(n_645) );
AND2x4_ASAP7_75t_SL g646 ( .A(n_607), .B(n_598), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_622), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_592), .B(n_572), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_572), .B(n_586), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_633), .B(n_636), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_586), .B(n_609), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_588), .B(n_631), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_623), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_607), .B(n_576), .Y(n_655) );
BUFx3_ASAP7_75t_L g656 ( .A(n_610), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_620), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_635), .B(n_589), .Y(n_658) );
NAND2x1p5_ASAP7_75t_L g659 ( .A(n_618), .B(n_582), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_616), .Y(n_660) );
AND2x4_ASAP7_75t_L g661 ( .A(n_610), .B(n_611), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_624), .Y(n_662) );
BUFx3_ASAP7_75t_L g663 ( .A(n_603), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_628), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_577), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_606), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_583), .Y(n_667) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_594), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_571), .B(n_578), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_575), .B(n_605), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_581), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_637), .Y(n_672) );
NOR2x1p5_ASAP7_75t_L g673 ( .A(n_600), .B(n_584), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_581), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_626), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_627), .Y(n_676) );
AND2x4_ASAP7_75t_L g677 ( .A(n_611), .B(n_584), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_627), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_625), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_604), .B(n_608), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_625), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_604), .B(n_608), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_579), .B(n_597), .Y(n_683) );
OR2x6_ASAP7_75t_L g684 ( .A(n_613), .B(n_612), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_618), .B(n_595), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_629), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_629), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_638), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_638), .Y(n_689) );
AND2x2_ASAP7_75t_L g690 ( .A(n_596), .B(n_599), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_638), .Y(n_691) );
OR2x2_ASAP7_75t_L g692 ( .A(n_601), .B(n_617), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_601), .B(n_587), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_640), .B(n_621), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_660), .B(n_614), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_643), .Y(n_696) );
HB1xp67_ASAP7_75t_L g697 ( .A(n_668), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_660), .B(n_580), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_647), .Y(n_699) );
INVx2_ASAP7_75t_SL g700 ( .A(n_646), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_647), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_648), .Y(n_702) );
INVx4_ASAP7_75t_L g703 ( .A(n_655), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_664), .B(n_593), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_664), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_669), .B(n_630), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_679), .B(n_681), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_684), .Y(n_708) );
NAND2x1p5_ASAP7_75t_SL g709 ( .A(n_693), .B(n_690), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_662), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_657), .Y(n_711) );
OR2x2_ASAP7_75t_L g712 ( .A(n_669), .B(n_665), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_665), .B(n_649), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_670), .B(n_645), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_651), .B(n_693), .Y(n_715) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_653), .Y(n_716) );
INVx1_ASAP7_75t_SL g717 ( .A(n_663), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_639), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_639), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_690), .B(n_641), .Y(n_720) );
INVx5_ASAP7_75t_L g721 ( .A(n_655), .Y(n_721) );
OR2x2_ASAP7_75t_L g722 ( .A(n_683), .B(n_652), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_676), .B(n_678), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_676), .B(n_678), .Y(n_724) );
BUFx3_ASAP7_75t_L g725 ( .A(n_646), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_683), .B(n_652), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_675), .B(n_692), .Y(n_727) );
AND2x2_ASAP7_75t_L g728 ( .A(n_692), .B(n_658), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_650), .B(n_667), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_658), .B(n_689), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_715), .B(n_687), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_696), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_696), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_718), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_714), .B(n_650), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_715), .B(n_686), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_711), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_728), .B(n_686), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_728), .B(n_686), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_730), .B(n_687), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_722), .B(n_691), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g742 ( .A(n_725), .B(n_642), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_718), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_719), .Y(n_744) );
INVx2_ASAP7_75t_SL g745 ( .A(n_717), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_699), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_730), .B(n_688), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_719), .Y(n_748) );
OR2x2_ASAP7_75t_L g749 ( .A(n_726), .B(n_688), .Y(n_749) );
BUFx2_ASAP7_75t_L g750 ( .A(n_703), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_707), .B(n_674), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_697), .Y(n_752) );
INVx2_ASAP7_75t_SL g753 ( .A(n_725), .Y(n_753) );
BUFx3_ASAP7_75t_L g754 ( .A(n_725), .Y(n_754) );
INVxp67_ASAP7_75t_L g755 ( .A(n_729), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_701), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_701), .Y(n_757) );
AOI21xp5_ASAP7_75t_SL g758 ( .A1(n_700), .A2(n_655), .B(n_673), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_716), .B(n_666), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_710), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_727), .B(n_671), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_720), .B(n_644), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_710), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_705), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_720), .B(n_644), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_727), .B(n_671), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_709), .B(n_672), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_732), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_733), .Y(n_769) );
OR2x6_ASAP7_75t_L g770 ( .A(n_758), .B(n_703), .Y(n_770) );
INVx2_ASAP7_75t_SL g771 ( .A(n_745), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_737), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_752), .B(n_702), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_735), .B(n_712), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_762), .B(n_712), .Y(n_775) );
AND2x4_ASAP7_75t_L g776 ( .A(n_750), .B(n_708), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_765), .B(n_713), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_731), .B(n_736), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_751), .B(n_694), .Y(n_779) );
INVx2_ASAP7_75t_SL g780 ( .A(n_745), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_737), .Y(n_781) );
INVx3_ASAP7_75t_SL g782 ( .A(n_753), .Y(n_782) );
AND2x2_ASAP7_75t_L g783 ( .A(n_738), .B(n_695), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_738), .B(n_704), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g785 ( .A(n_755), .B(n_706), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_746), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_754), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_773), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_768), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g790 ( .A1(n_785), .A2(n_766), .B(n_761), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g791 ( .A(n_782), .B(n_721), .Y(n_791) );
OAI332xp33_ASAP7_75t_L g792 ( .A1(n_785), .A2(n_749), .A3(n_741), .B1(n_759), .B2(n_767), .B3(n_760), .C1(n_763), .C2(n_764), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_769), .Y(n_793) );
AOI21xp5_ASAP7_75t_L g794 ( .A1(n_770), .A2(n_721), .B(n_742), .Y(n_794) );
INVx2_ASAP7_75t_L g795 ( .A(n_772), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_778), .B(n_739), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_776), .A2(n_747), .B1(n_740), .B2(n_723), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g798 ( .A1(n_779), .A2(n_709), .B1(n_756), .B2(n_757), .C(n_744), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_795), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_792), .B(n_783), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g801 ( .A1(n_790), .A2(n_776), .B1(n_780), .B2(n_771), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_791), .A2(n_780), .B(n_787), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_797), .A2(n_782), .B1(n_777), .B2(n_774), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_789), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_793), .Y(n_805) );
HB1xp67_ASAP7_75t_L g806 ( .A(n_796), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_788), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_791), .B(n_772), .Y(n_808) );
INVx2_ASAP7_75t_SL g809 ( .A(n_795), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_798), .B(n_784), .Y(n_810) );
NAND2xp5_ASAP7_75t_SL g811 ( .A(n_794), .B(n_781), .Y(n_811) );
INVx2_ASAP7_75t_L g812 ( .A(n_809), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_806), .Y(n_813) );
HB1xp67_ASAP7_75t_L g814 ( .A(n_809), .Y(n_814) );
OAI222xp33_ASAP7_75t_L g815 ( .A1(n_800), .A2(n_801), .B1(n_803), .B2(n_810), .C1(n_811), .C2(n_802), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_804), .Y(n_816) );
XOR2xp5_ASAP7_75t_L g817 ( .A(n_807), .B(n_775), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_815), .A2(n_805), .B1(n_799), .B2(n_808), .C(n_786), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_814), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_813), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_816), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g822 ( .A(n_820), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_819), .Y(n_823) );
NAND4xp75_ASAP7_75t_L g824 ( .A(n_818), .B(n_812), .C(n_685), .D(n_682), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_821), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_823), .Y(n_826) );
AOI311xp33_ASAP7_75t_L g827 ( .A1(n_825), .A2(n_817), .A3(n_734), .B(n_748), .C(n_743), .Y(n_827) );
BUFx2_ASAP7_75t_L g828 ( .A(n_822), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_828), .A2(n_822), .B1(n_824), .B2(n_680), .Y(n_829) );
NAND4xp25_ASAP7_75t_L g830 ( .A(n_826), .B(n_682), .C(n_680), .D(n_685), .Y(n_830) );
AND2x2_ASAP7_75t_SL g831 ( .A(n_829), .B(n_827), .Y(n_831) );
OAI22xp5_ASAP7_75t_SL g832 ( .A1(n_831), .A2(n_830), .B1(n_659), .B2(n_656), .Y(n_832) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_832), .A2(n_677), .B1(n_656), .B2(n_661), .C1(n_698), .C2(n_654), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_833), .A2(n_656), .B1(n_661), .B2(n_724), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_834), .A2(n_661), .B1(n_724), .B2(n_723), .Y(n_835) );
endmodule