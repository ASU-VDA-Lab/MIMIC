module real_aes_1705_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_546;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g100 ( .A1(n_0), .A2(n_57), .B1(n_88), .B2(n_101), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_1), .A2(n_49), .B1(n_150), .B2(n_152), .Y(n_149) );
INVx1_ASAP7_75t_L g164 ( .A(n_2), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_3), .B(n_191), .Y(n_214) );
INVx1_ASAP7_75t_L g236 ( .A(n_4), .Y(n_236) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_5), .A2(n_17), .B1(n_88), .B2(n_98), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_6), .Y(n_252) );
INVx2_ASAP7_75t_L g190 ( .A(n_7), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g550 ( .A1(n_8), .A2(n_62), .B1(n_551), .B2(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g552 ( .A(n_8), .Y(n_552) );
INVx1_ASAP7_75t_L g224 ( .A(n_9), .Y(n_224) );
INVx1_ASAP7_75t_L g221 ( .A(n_10), .Y(n_221) );
INVx1_ASAP7_75t_SL g296 ( .A(n_11), .Y(n_296) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_12), .B(n_201), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g109 ( .A1(n_13), .A2(n_51), .B1(n_110), .B2(n_114), .Y(n_109) );
AOI33xp33_ASAP7_75t_L g273 ( .A1(n_14), .A2(n_38), .A3(n_181), .B1(n_196), .B2(n_274), .B3(n_275), .Y(n_273) );
INVx1_ASAP7_75t_L g245 ( .A(n_15), .Y(n_245) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_16), .A2(n_18), .B1(n_125), .B2(n_128), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_17), .A2(n_57), .B1(n_60), .B2(n_556), .C(n_558), .Y(n_555) );
OA21x2_ASAP7_75t_L g189 ( .A1(n_19), .A2(n_70), .B(n_190), .Y(n_189) );
OR2x2_ASAP7_75t_L g192 ( .A(n_19), .B(n_70), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_20), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_20), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_21), .B(n_234), .Y(n_293) );
AOI22xp33_ASAP7_75t_L g142 ( .A1(n_22), .A2(n_43), .B1(n_143), .B2(n_145), .Y(n_142) );
INVx3_ASAP7_75t_L g88 ( .A(n_23), .Y(n_88) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_24), .A2(n_37), .B1(n_119), .B2(n_121), .Y(n_118) );
INVx1_ASAP7_75t_SL g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g166 ( .A(n_26), .Y(n_166) );
AND2x2_ASAP7_75t_L g185 ( .A(n_26), .B(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_L g210 ( .A(n_26), .B(n_164), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_27), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_28), .B(n_234), .Y(n_260) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_29), .A2(n_178), .B1(n_188), .B2(n_191), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_30), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_31), .B(n_201), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_32), .A2(n_80), .B1(n_159), .B2(n_160), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_32), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_33), .B(n_212), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_34), .B(n_201), .Y(n_237) );
AO22x2_ASAP7_75t_L g87 ( .A1(n_35), .A2(n_60), .B1(n_88), .B2(n_89), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_36), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_39), .B(n_201), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_40), .A2(n_53), .B1(n_84), .B2(n_102), .Y(n_83) );
INVx1_ASAP7_75t_L g182 ( .A(n_41), .Y(n_182) );
INVx1_ASAP7_75t_L g203 ( .A(n_41), .Y(n_203) );
AND2x2_ASAP7_75t_L g265 ( .A(n_42), .B(n_266), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g233 ( .A1(n_44), .A2(n_63), .B1(n_194), .B2(n_234), .C(n_235), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_45), .B(n_234), .Y(n_288) );
INVx1_ASAP7_75t_L g94 ( .A(n_46), .Y(n_94) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_47), .B(n_188), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_47), .A2(n_541), .B1(n_554), .B2(n_562), .Y(n_540) );
INVx1_ASAP7_75t_L g568 ( .A(n_47), .Y(n_568) );
AOI21xp5_ASAP7_75t_SL g284 ( .A1(n_48), .A2(n_194), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g217 ( .A(n_50), .Y(n_217) );
INVx1_ASAP7_75t_L g263 ( .A(n_52), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_54), .A2(n_61), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_54), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_55), .A2(n_194), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_56), .B(n_156), .Y(n_155) );
INVxp33_ASAP7_75t_L g560 ( .A(n_57), .Y(n_560) );
INVx1_ASAP7_75t_L g186 ( .A(n_58), .Y(n_186) );
INVx1_ASAP7_75t_L g205 ( .A(n_58), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_59), .A2(n_76), .B1(n_134), .B2(n_137), .Y(n_133) );
INVxp67_ASAP7_75t_L g559 ( .A(n_60), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_61), .B(n_234), .Y(n_276) );
INVx1_ASAP7_75t_L g545 ( .A(n_61), .Y(n_545) );
INVx1_ASAP7_75t_L g551 ( .A(n_62), .Y(n_551) );
AND2x2_ASAP7_75t_L g298 ( .A(n_64), .B(n_241), .Y(n_298) );
INVx1_ASAP7_75t_L g218 ( .A(n_65), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_66), .A2(n_194), .B(n_295), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g193 ( .A1(n_67), .A2(n_194), .B(n_199), .C(n_211), .Y(n_193) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_68), .B(n_241), .Y(n_282) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_69), .A2(n_194), .B1(n_271), .B2(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g286 ( .A(n_71), .Y(n_286) );
AND2x2_ASAP7_75t_L g277 ( .A(n_72), .B(n_241), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_73), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
BUFx2_ASAP7_75t_SL g557 ( .A(n_74), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_75), .B(n_201), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_161), .B1(n_167), .B2(n_538), .C(n_539), .Y(n_77) );
INVxp67_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_80), .Y(n_160) );
OAI222xp33_ASAP7_75t_L g539 ( .A1(n_80), .A2(n_160), .B1(n_252), .B2(n_540), .C1(n_567), .C2(n_570), .Y(n_539) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2xp67_ASAP7_75t_L g81 ( .A(n_82), .B(n_132), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_109), .C(n_118), .D(n_124), .Y(n_82) );
BUFx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
AND2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_95), .Y(n_85) );
AND2x2_ASAP7_75t_L g120 ( .A(n_86), .B(n_107), .Y(n_120) );
AND2x4_ASAP7_75t_L g144 ( .A(n_86), .B(n_131), .Y(n_144) );
AND2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
INVx2_ASAP7_75t_L g106 ( .A(n_87), .Y(n_106) );
BUFx2_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
AND2x2_ASAP7_75t_L g139 ( .A(n_87), .B(n_91), .Y(n_139) );
INVx1_ASAP7_75t_L g89 ( .A(n_88), .Y(n_89) );
OAI22x1_ASAP7_75t_L g91 ( .A1(n_88), .A2(n_92), .B1(n_93), .B2(n_94), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_88), .Y(n_92) );
INVx2_ASAP7_75t_L g98 ( .A(n_88), .Y(n_98) );
INVx1_ASAP7_75t_L g101 ( .A(n_88), .Y(n_101) );
AND2x4_ASAP7_75t_L g105 ( .A(n_90), .B(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
AND2x2_ASAP7_75t_L g113 ( .A(n_91), .B(n_106), .Y(n_113) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_91), .Y(n_154) );
AND2x4_ASAP7_75t_L g112 ( .A(n_95), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g127 ( .A(n_95), .B(n_105), .Y(n_127) );
AND2x2_ASAP7_75t_L g158 ( .A(n_95), .B(n_139), .Y(n_158) );
AND2x4_ASAP7_75t_L g95 ( .A(n_96), .B(n_99), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
INVx1_ASAP7_75t_L g108 ( .A(n_97), .Y(n_108) );
AND2x2_ASAP7_75t_L g117 ( .A(n_97), .B(n_100), .Y(n_117) );
AND2x4_ASAP7_75t_L g131 ( .A(n_97), .B(n_99), .Y(n_131) );
INVxp67_ASAP7_75t_L g148 ( .A(n_99), .Y(n_148) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x2_ASAP7_75t_L g107 ( .A(n_100), .B(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx8_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_107), .Y(n_104) );
AND2x4_ASAP7_75t_L g116 ( .A(n_105), .B(n_117), .Y(n_116) );
AND2x4_ASAP7_75t_L g130 ( .A(n_105), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g136 ( .A(n_107), .B(n_113), .Y(n_136) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_108), .Y(n_141) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx6_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g151 ( .A(n_113), .B(n_131), .Y(n_151) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
AND2x4_ASAP7_75t_L g122 ( .A(n_117), .B(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g153 ( .A(n_117), .B(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
INVx8_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NAND4xp25_ASAP7_75t_L g132 ( .A(n_133), .B(n_142), .C(n_149), .D(n_155), .Y(n_132) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx4f_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
AND2x4_ASAP7_75t_L g147 ( .A(n_139), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx3_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx12f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx6_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OR2x2_ASAP7_75t_SL g162 ( .A(n_163), .B(n_165), .Y(n_162) );
AND2x2_ASAP7_75t_L g180 ( .A(n_163), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g561 ( .A(n_163), .Y(n_561) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AND2x2_ASAP7_75t_L g198 ( .A(n_164), .B(n_182), .Y(n_198) );
AND3x1_ASAP7_75t_SL g554 ( .A(n_165), .B(n_555), .C(n_561), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_165), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NOR2x1p5_ASAP7_75t_L g195 ( .A(n_166), .B(n_196), .Y(n_195) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_170), .B(n_472), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_171), .B(n_395), .Y(n_170) );
NAND3xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_342), .C(n_375), .Y(n_171) );
AOI211xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_299), .B(n_308), .C(n_332), .Y(n_172) );
OAI21xp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_228), .B(n_278), .Y(n_173) );
OR2x2_ASAP7_75t_L g352 ( .A(n_174), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g507 ( .A(n_174), .B(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_175), .A2(n_398), .B1(n_402), .B2(n_404), .Y(n_397) );
AND2x2_ASAP7_75t_L g434 ( .A(n_175), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_213), .Y(n_175) );
INVx1_ASAP7_75t_L g331 ( .A(n_176), .Y(n_331) );
AND2x4_ASAP7_75t_L g348 ( .A(n_176), .B(n_329), .Y(n_348) );
INVx2_ASAP7_75t_L g370 ( .A(n_176), .Y(n_370) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_176), .Y(n_453) );
AND2x2_ASAP7_75t_L g524 ( .A(n_176), .B(n_281), .Y(n_524) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_193), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_183), .C(n_187), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g571 ( .A1(n_179), .A2(n_561), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x4_ASAP7_75t_L g234 ( .A(n_180), .B(n_184), .Y(n_234) );
OR2x6_ASAP7_75t_L g208 ( .A(n_181), .B(n_197), .Y(n_208) );
INVxp33_ASAP7_75t_L g274 ( .A(n_181), .Y(n_274) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x4_ASAP7_75t_L g226 ( .A(n_182), .B(n_204), .Y(n_226) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g197 ( .A(n_186), .Y(n_197) );
AND2x6_ASAP7_75t_L g223 ( .A(n_186), .B(n_202), .Y(n_223) );
INVx4_ASAP7_75t_L g241 ( .A(n_188), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_188), .B(n_251), .Y(n_250) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_189), .Y(n_212) );
AND2x4_ASAP7_75t_L g191 ( .A(n_190), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_190), .B(n_192), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_191), .B(n_209), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_191), .A2(n_284), .B(n_288), .Y(n_283) );
INVxp67_ASAP7_75t_L g253 ( .A(n_194), .Y(n_253) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_194), .Y(n_538) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_198), .Y(n_194) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_195), .Y(n_572) );
INVx1_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
INVx3_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_200), .A2(n_206), .B(n_209), .Y(n_199) );
INVx1_ASAP7_75t_L g219 ( .A(n_201), .Y(n_219) );
AND2x4_ASAP7_75t_L g201 ( .A(n_202), .B(n_204), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_208), .A2(n_217), .B1(n_218), .B2(n_219), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_208), .A2(n_209), .B(n_236), .C(n_237), .Y(n_235) );
INVxp67_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_208), .A2(n_209), .B(n_263), .C(n_264), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g285 ( .A1(n_208), .A2(n_209), .B(n_286), .C(n_287), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_SL g295 ( .A1(n_208), .A2(n_209), .B(n_296), .C(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g271 ( .A(n_209), .Y(n_271) );
INVx5_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_210), .Y(n_246) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_211), .A2(n_269), .B(n_277), .Y(n_268) );
AO21x2_ASAP7_75t_L g313 ( .A1(n_211), .A2(n_269), .B(n_277), .Y(n_313) );
INVx2_ASAP7_75t_SL g211 ( .A(n_212), .Y(n_211) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_212), .A2(n_233), .B(n_238), .Y(n_232) );
AND2x2_ASAP7_75t_L g289 ( .A(n_213), .B(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g318 ( .A(n_213), .Y(n_318) );
INVx3_ASAP7_75t_L g329 ( .A(n_213), .Y(n_329) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_220), .B(n_227), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_219), .B(n_245), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B1(n_224), .B2(n_225), .Y(n_220) );
INVxp67_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVxp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_228), .A2(n_519), .B1(n_521), .B2(n_523), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_228), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_SL g228 ( .A(n_229), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_256), .Y(n_229) );
INVx3_ASAP7_75t_L g302 ( .A(n_230), .Y(n_302) );
AND2x2_ASAP7_75t_L g310 ( .A(n_230), .B(n_311), .Y(n_310) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_230), .Y(n_340) );
NAND2x1_ASAP7_75t_SL g534 ( .A(n_230), .B(n_301), .Y(n_534) );
AND2x4_ASAP7_75t_L g230 ( .A(n_231), .B(n_239), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g307 ( .A(n_232), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_232), .B(n_313), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_232), .B(n_239), .Y(n_338) );
AND2x4_ASAP7_75t_L g345 ( .A(n_232), .B(n_346), .Y(n_345) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_232), .Y(n_394) );
INVxp67_ASAP7_75t_L g401 ( .A(n_232), .Y(n_401) );
INVx1_ASAP7_75t_L g406 ( .A(n_232), .Y(n_406) );
INVx1_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
INVx1_ASAP7_75t_L g305 ( .A(n_239), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_239), .B(n_315), .Y(n_324) );
INVx2_ASAP7_75t_L g392 ( .A(n_239), .Y(n_392) );
INVx1_ASAP7_75t_L g431 ( .A(n_239), .Y(n_431) );
OR2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_249), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B1(n_247), .B2(n_248), .Y(n_240) );
INVx3_ASAP7_75t_L g248 ( .A(n_241), .Y(n_248) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_248), .A2(n_259), .B(n_265), .Y(n_258) );
AO21x2_ASAP7_75t_L g315 ( .A1(n_248), .A2(n_259), .B(n_265), .Y(n_315) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_253), .B1(n_254), .B2(n_255), .Y(n_249) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g361 ( .A(n_256), .B(n_338), .Y(n_361) );
AND2x2_ASAP7_75t_L g429 ( .A(n_256), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g443 ( .A(n_256), .B(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_256), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_268), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2x1_ASAP7_75t_L g306 ( .A(n_258), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g399 ( .A(n_258), .B(n_392), .Y(n_399) );
AND2x2_ASAP7_75t_L g490 ( .A(n_258), .B(n_312), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_266), .Y(n_291) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g301 ( .A(n_268), .Y(n_301) );
INVx2_ASAP7_75t_L g346 ( .A(n_268), .Y(n_346) );
AND2x2_ASAP7_75t_L g391 ( .A(n_268), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_270), .B(n_276), .Y(n_269) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_289), .Y(n_279) );
AND2x2_ASAP7_75t_L g433 ( .A(n_280), .B(n_434), .Y(n_433) );
OR2x6_ASAP7_75t_L g492 ( .A(n_280), .B(n_493), .Y(n_492) );
BUFx6f_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx4_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
AND2x4_ASAP7_75t_L g330 ( .A(n_281), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g365 ( .A(n_281), .B(n_290), .Y(n_365) );
INVx2_ASAP7_75t_L g414 ( .A(n_281), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_281), .B(n_388), .Y(n_463) );
AND2x2_ASAP7_75t_L g500 ( .A(n_281), .B(n_318), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_281), .B(n_383), .Y(n_508) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g341 ( .A(n_289), .B(n_330), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_289), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_289), .B(n_368), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_289), .B(n_381), .Y(n_502) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_290), .Y(n_320) );
AND2x2_ASAP7_75t_L g328 ( .A(n_290), .B(n_329), .Y(n_328) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_290), .Y(n_351) );
INVx2_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
INVx1_ASAP7_75t_L g387 ( .A(n_290), .Y(n_387) );
INVx1_ASAP7_75t_L g435 ( .A(n_290), .Y(n_435) );
AO21x2_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_298), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
NAND2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
OR2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_301), .B(n_304), .Y(n_377) );
OR2x2_ASAP7_75t_L g449 ( .A(n_301), .B(n_450), .Y(n_449) );
AND4x1_ASAP7_75t_SL g495 ( .A(n_301), .B(n_477), .C(n_496), .D(n_497), .Y(n_495) );
OR2x2_ASAP7_75t_L g519 ( .A(n_302), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
AND2x2_ASAP7_75t_L g356 ( .A(n_305), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_305), .B(n_314), .Y(n_506) );
AND2x2_ASAP7_75t_L g531 ( .A(n_306), .B(n_391), .Y(n_531) );
OAI32xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_316), .A3(n_321), .B1(n_323), .B2(n_326), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g404 ( .A(n_311), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g504 ( .A(n_311), .B(n_458), .Y(n_504) );
AND2x4_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
AND2x2_ASAP7_75t_L g400 ( .A(n_312), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g486 ( .A(n_312), .Y(n_486) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_313), .B(n_315), .Y(n_520) );
INVx3_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g515 ( .A(n_314), .B(n_442), .Y(n_515) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_315), .Y(n_374) );
AND2x2_ASAP7_75t_L g393 ( .A(n_315), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g527 ( .A(n_317), .Y(n_527) );
NAND2x1_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g367 ( .A(n_318), .Y(n_367) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_318), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_321), .B(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_327), .Y(n_359) );
AND2x4_ASAP7_75t_L g381 ( .A(n_322), .B(n_331), .Y(n_381) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_322), .B(n_453), .Y(n_452) );
NOR2x1_ASAP7_75t_L g478 ( .A(n_322), .B(n_403), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g445 ( .A1(n_323), .A2(n_446), .B1(n_449), .B2(n_451), .Y(n_445) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_SL g465 ( .A(n_324), .Y(n_465) );
INVx2_ASAP7_75t_L g357 ( .A(n_325), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_330), .Y(n_326) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_328), .B(n_334), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g466 ( .A1(n_328), .A2(n_464), .B1(n_467), .B2(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
AND2x2_ASAP7_75t_L g411 ( .A(n_329), .B(n_370), .Y(n_411) );
INVx2_ASAP7_75t_L g334 ( .A(n_330), .Y(n_334) );
OAI21xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_335), .B(n_339), .Y(n_332) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_336), .A2(n_408), .B1(n_412), .B2(n_413), .Y(n_407) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_337), .B(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_337), .B(n_405), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_337), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NOR3xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_358), .C(n_362), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_347), .B1(n_352), .B2(n_355), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g372 ( .A(n_345), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_399), .Y(n_412) );
AND2x2_ASAP7_75t_L g464 ( .A(n_345), .B(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g481 ( .A(n_345), .B(n_431), .Y(n_481) );
AND2x2_ASAP7_75t_L g536 ( .A(n_345), .B(n_430), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx4_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
AND2x2_ASAP7_75t_L g413 ( .A(n_348), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g418 ( .A(n_351), .Y(n_418) );
AND2x2_ASAP7_75t_L g427 ( .A(n_351), .B(n_411), .Y(n_427) );
INVx1_ASAP7_75t_L g462 ( .A(n_353), .Y(n_462) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g383 ( .A(n_354), .Y(n_383) );
INVxp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_356), .B(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_357), .B(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_366), .B(n_371), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_364), .B(n_403), .Y(n_512) );
INVx2_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_367), .A2(n_376), .B(n_378), .Y(n_375) );
AND2x2_ASAP7_75t_L g522 ( .A(n_367), .B(n_381), .Y(n_522) );
AND2x4_ASAP7_75t_L g385 ( .A(n_368), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g419 ( .A(n_368), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_368), .B(n_435), .Y(n_501) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_384), .B(n_389), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_381), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_381), .B(n_386), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_382), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g444 ( .A(n_382), .Y(n_444) );
INVx1_ASAP7_75t_L g448 ( .A(n_382), .Y(n_448) );
AND2x2_ASAP7_75t_L g532 ( .A(n_382), .B(n_500), .Y(n_532) );
AND2x2_ASAP7_75t_L g535 ( .A(n_382), .B(n_452), .Y(n_535) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x4_ASAP7_75t_SL g386 ( .A(n_387), .B(n_388), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_387), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g514 ( .A(n_391), .Y(n_514) );
AND2x2_ASAP7_75t_L g405 ( .A(n_392), .B(n_406), .Y(n_405) );
NAND4xp75_ASAP7_75t_L g395 ( .A(n_396), .B(n_415), .C(n_436), .D(n_454), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_407), .Y(n_396) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_399), .B(n_486), .Y(n_485) );
NAND2x1p5_ASAP7_75t_L g471 ( .A(n_400), .B(n_465), .Y(n_471) );
NAND2xp5_ASAP7_75t_R g487 ( .A(n_403), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g537 ( .A(n_403), .Y(n_537) );
INVx2_ASAP7_75t_L g450 ( .A(n_405), .Y(n_450) );
BUFx3_ASAP7_75t_L g442 ( .A(n_406), .Y(n_442) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g493 ( .A(n_411), .Y(n_493) );
AND2x2_ASAP7_75t_L g447 ( .A(n_413), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g469 ( .A(n_414), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_420), .B(n_422), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_418), .B(n_452), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_419), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_421), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_426), .B1(n_428), .B2(n_432), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_430), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g489 ( .A(n_431), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g497 ( .A(n_431), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_432), .B(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g467 ( .A(n_435), .B(n_468), .Y(n_467) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_443), .B(n_445), .Y(n_436) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g484 ( .A(n_441), .B(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_448), .Y(n_496) );
INVx2_ASAP7_75t_SL g488 ( .A(n_452), .Y(n_488) );
AND2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_459), .B1(n_461), .B2(n_464), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_509), .Y(n_472) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_482), .C(n_494), .Y(n_473) );
NOR2x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_479), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g482 ( .A1(n_483), .A2(n_487), .B1(n_489), .B2(n_491), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .C(n_505), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_502), .B(n_503), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_528), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_518), .C(n_525), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B1(n_516), .B2(n_517), .Y(n_511) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_515), .Y(n_513) );
NOR3xp33_ASAP7_75t_L g525 ( .A(n_519), .B(n_524), .C(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI222xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_532), .B1(n_533), .B2(n_535), .C1(n_536), .C2(n_537), .Y(n_528) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
INVx2_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_542), .A2(n_554), .B1(n_568), .B2(n_569), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_544), .B1(n_547), .B2(n_553), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_544), .Y(n_543) );
CKINVDCx16_ASAP7_75t_R g553 ( .A(n_547), .Y(n_553) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVxp67_ASAP7_75t_L g566 ( .A(n_555), .Y(n_566) );
CKINVDCx8_ASAP7_75t_R g556 ( .A(n_557), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
CKINVDCx16_ASAP7_75t_R g564 ( .A(n_561), .Y(n_564) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_563), .Y(n_569) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_571), .Y(n_570) );
endmodule