module fake_jpeg_8475_n_65 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_65);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_65;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_31),
.B(n_1),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_2),
.Y(n_38)
);

NOR2xp67_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_4),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_29),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_2),
.B(n_3),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_50),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_29),
.B1(n_32),
.B2(n_30),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_55)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_15),
.B1(n_22),
.B2(n_21),
.Y(n_49)
);

AND2x6_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_36),
.A2(n_13),
.B1(n_20),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_5),
.C(n_7),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_56),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_46),
.Y(n_56)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_55),
.C(n_54),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_57),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_41),
.Y(n_63)
);

AOI322xp5_ASAP7_75t_L g64 ( 
.A1(n_63),
.A2(n_56),
.A3(n_58),
.B1(n_46),
.B2(n_43),
.C1(n_23),
.C2(n_16),
.Y(n_64)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);


endmodule