module fake_netlist_6_4156_n_1598 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1598);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1598;

wire n_992;
wire n_801;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_250;
wire n_544;
wire n_1140;
wire n_1444;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1069;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_1412;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1388;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_1207;
wire n_683;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1224;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1437;
wire n_385;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_1429;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1024;
wire n_248;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_785;
wire n_746;
wire n_609;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_1350;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_1346;
wire n_711;
wire n_579;
wire n_1352;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_1121;
wire n_330;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_482;
wire n_934;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_1574;
wire n_240;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1240;

BUFx3_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_6),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_217),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_21),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_214),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_102),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_135),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_150),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_162),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_67),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_2),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_79),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_33),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_204),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_107),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_171),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_105),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_114),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_215),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_72),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_77),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_86),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_137),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_180),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_108),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_218),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_167),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_126),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_85),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_193),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_223),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_196),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_194),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_181),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_178),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_186),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_177),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_173),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_168),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_87),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_205),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_35),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_161),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_64),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_138),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_170),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_198),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_157),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_212),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_11),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_151),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_148),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_113),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_48),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_145),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_52),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_8),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_100),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_190),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_91),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_82),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_140),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_60),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_120),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_143),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_43),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_26),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_110),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_58),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_160),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_65),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_128),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_192),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_30),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_78),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_15),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_15),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_34),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_208),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_83),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_207),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_5),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_154),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_189),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_197),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_201),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_40),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_30),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_134),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_175),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_191),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_89),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_21),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_93),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_13),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_37),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_56),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_27),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_75),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_60),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_125),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_50),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_132),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_159),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_57),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_56),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_129),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_59),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_147),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_206),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_58),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_44),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_210),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_31),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_22),
.Y(n_361)
);

BUFx8_ASAP7_75t_SL g362 ( 
.A(n_139),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_84),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_133),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_8),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_225),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_41),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_32),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_19),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_142),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_24),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_16),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_315),
.B(n_0),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_226),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_221),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_253),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_226),
.B(n_327),
.Y(n_377)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_253),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_253),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_228),
.Y(n_380)
);

AND2x6_ASAP7_75t_L g381 ( 
.A(n_253),
.B(n_74),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_234),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_328),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_0),
.Y(n_385)
);

BUFx12f_ASAP7_75t_L g386 ( 
.A(n_227),
.Y(n_386)
);

BUFx12f_ASAP7_75t_L g387 ( 
.A(n_227),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_1),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_294),
.B(n_1),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_253),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_294),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_240),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_242),
.B(n_2),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_239),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_328),
.Y(n_395)
);

BUFx8_ASAP7_75t_SL g396 ( 
.A(n_362),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_242),
.B(n_3),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_285),
.B(n_3),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_285),
.B(n_4),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_300),
.B(n_4),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_332),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_286),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_300),
.B(n_5),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

BUFx12f_ASAP7_75t_L g405 ( 
.A(n_230),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_302),
.B(n_6),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_302),
.B(n_76),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_314),
.B(n_220),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_286),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_314),
.B(n_7),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_349),
.B(n_80),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_248),
.Y(n_412)
);

AND2x4_ASAP7_75t_L g413 ( 
.A(n_251),
.B(n_88),
.Y(n_413)
);

BUFx12f_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx5_ASAP7_75t_L g415 ( 
.A(n_286),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_332),
.B(n_7),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_286),
.Y(n_417)
);

BUFx12f_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_243),
.Y(n_421)
);

BUFx12f_ASAP7_75t_L g422 ( 
.A(n_230),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_255),
.B(n_9),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_281),
.Y(n_424)
);

AND2x4_ASAP7_75t_L g425 ( 
.A(n_257),
.B(n_259),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_328),
.B(n_9),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_328),
.B(n_10),
.Y(n_428)
);

BUFx12f_ASAP7_75t_L g429 ( 
.A(n_232),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_328),
.B(n_10),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_263),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_264),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_328),
.B(n_267),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_273),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_232),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_328),
.B(n_11),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_299),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_308),
.B(n_12),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_275),
.B(n_12),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_277),
.B(n_219),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_371),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_309),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_287),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_319),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_288),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_307),
.B(n_13),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_323),
.B(n_14),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_316),
.B(n_14),
.Y(n_449)
);

AND2x6_ASAP7_75t_L g450 ( 
.A(n_325),
.B(n_90),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_229),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_334),
.B(n_337),
.Y(n_452)
);

BUFx12f_ASAP7_75t_L g453 ( 
.A(n_241),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_324),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_333),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_338),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_340),
.Y(n_457)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_289),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_353),
.B(n_17),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_339),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_377),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_376),
.Y(n_462)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_385),
.A2(n_365),
.B1(n_369),
.B2(n_368),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_231),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_342),
.B1(n_369),
.B2(n_368),
.Y(n_465)
);

AND2x2_ASAP7_75t_SL g466 ( 
.A(n_375),
.B(n_370),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_376),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_412),
.B(n_229),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_447),
.A2(n_449),
.B1(n_459),
.B2(n_373),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

AO22x2_ASAP7_75t_L g471 ( 
.A1(n_375),
.A2(n_367),
.B1(n_341),
.B2(n_351),
.Y(n_471)
);

OA22x2_ASAP7_75t_L g472 ( 
.A1(n_377),
.A2(n_360),
.B1(n_365),
.B2(n_241),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_376),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_393),
.A2(n_358),
.B1(n_256),
.B2(n_357),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_374),
.B(n_383),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_399),
.A2(n_358),
.B1(n_256),
.B2(n_357),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_403),
.A2(n_354),
.B1(n_361),
.B2(n_345),
.Y(n_477)
);

OAI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_397),
.A2(n_354),
.B1(n_361),
.B2(n_284),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_R g480 ( 
.A1(n_424),
.A2(n_278),
.B1(n_290),
.B2(n_292),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_423),
.A2(n_238),
.B1(n_260),
.B2(n_280),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_423),
.A2(n_301),
.B1(n_298),
.B2(n_296),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_233),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_451),
.B(n_233),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g485 ( 
.A1(n_398),
.A2(n_406),
.B1(n_410),
.B2(n_400),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_451),
.B(n_374),
.Y(n_486)
);

AO22x2_ASAP7_75t_L g487 ( 
.A1(n_375),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_376),
.Y(n_488)
);

OAI22xp33_ASAP7_75t_SL g489 ( 
.A1(n_426),
.A2(n_305),
.B1(n_311),
.B2(n_313),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_375),
.B(n_235),
.Y(n_490)
);

AO22x2_ASAP7_75t_L g491 ( 
.A1(n_407),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_491)
);

OAI22xp33_ASAP7_75t_L g492 ( 
.A1(n_439),
.A2(n_343),
.B1(n_317),
.B2(n_320),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_386),
.A2(n_344),
.B1(n_346),
.B2(n_322),
.Y(n_493)
);

OAI22xp33_ASAP7_75t_L g494 ( 
.A1(n_446),
.A2(n_348),
.B1(n_352),
.B2(n_366),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_383),
.B(n_235),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_428),
.A2(n_366),
.B1(n_364),
.B2(n_363),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_386),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

AO22x2_ASAP7_75t_L g499 ( 
.A1(n_407),
.A2(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_R g500 ( 
.A1(n_424),
.A2(n_23),
.B1(n_26),
.B2(n_27),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_430),
.A2(n_364),
.B1(n_363),
.B2(n_359),
.Y(n_501)
);

AO22x2_ASAP7_75t_L g502 ( 
.A1(n_407),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_379),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_407),
.A2(n_28),
.B1(n_29),
.B2(n_32),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_431),
.Y(n_505)
);

OA22x2_ASAP7_75t_L g506 ( 
.A1(n_392),
.A2(n_455),
.B1(n_421),
.B2(n_460),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_389),
.A2(n_359),
.B1(n_356),
.B2(n_355),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_379),
.Y(n_508)
);

OAI22xp33_ASAP7_75t_R g509 ( 
.A1(n_441),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_379),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_431),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_408),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_413),
.B(n_236),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_431),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_413),
.B(n_236),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_438),
.A2(n_356),
.B1(n_355),
.B2(n_244),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_436),
.A2(n_237),
.B1(n_244),
.B2(n_245),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_408),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_519)
);

OAI22xp33_ASAP7_75t_L g520 ( 
.A1(n_387),
.A2(n_237),
.B1(n_245),
.B2(n_246),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_396),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_380),
.B(n_246),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_380),
.B(n_247),
.Y(n_523)
);

NAND3x1_ASAP7_75t_L g524 ( 
.A(n_389),
.B(n_42),
.C(n_43),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_433),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_408),
.B(n_249),
.Y(n_526)
);

OA22x2_ASAP7_75t_L g527 ( 
.A1(n_460),
.A2(n_250),
.B1(n_252),
.B2(n_254),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_431),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_387),
.Y(n_529)
);

AO22x2_ASAP7_75t_L g530 ( 
.A1(n_408),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_382),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_470),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_505),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_461),
.B(n_413),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_511),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_469),
.B(n_405),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g537 ( 
.A(n_481),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_475),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_462),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_481),
.B(n_45),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_528),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_464),
.B(n_482),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_469),
.B(n_483),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_514),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_514),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_467),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_473),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_479),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_486),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_510),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_466),
.B(n_458),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_531),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_482),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_531),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_513),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_523),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_491),
.B(n_499),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_468),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_493),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_468),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_521),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_506),
.Y(n_568)
);

INVxp67_ASAP7_75t_SL g569 ( 
.A(n_516),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_506),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_495),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_507),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_471),
.Y(n_573)
);

XNOR2x2_ASAP7_75t_L g574 ( 
.A(n_491),
.B(n_416),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_471),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_513),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_493),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_521),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_484),
.B(n_405),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_497),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_526),
.B(n_425),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_490),
.B(n_425),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_472),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_499),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_477),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g587 ( 
.A(n_529),
.B(n_414),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_527),
.B(n_425),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_502),
.B(n_411),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_485),
.B(n_414),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_517),
.A2(n_411),
.B(n_440),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_524),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_527),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_517),
.B(n_411),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_558),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_578),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_561),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_540),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_591),
.B(n_525),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_411),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_593),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_548),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_582),
.B(n_416),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_566),
.B(n_504),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_548),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_573),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_583),
.B(n_425),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_549),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_583),
.B(n_452),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_L g615 ( 
.A1(n_545),
.A2(n_525),
.B(n_518),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_588),
.B(n_504),
.Y(n_616)
);

AND2x4_ASAP7_75t_SL g617 ( 
.A(n_561),
.B(n_452),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_588),
.B(n_582),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_569),
.B(n_452),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_549),
.Y(n_620)
);

INVx3_ASAP7_75t_SL g621 ( 
.A(n_589),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_551),
.B(n_512),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_575),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_561),
.B(n_518),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_452),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_551),
.B(n_512),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

INVx3_ASAP7_75t_SL g628 ( 
.A(n_589),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_539),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_580),
.B(n_519),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_550),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_580),
.B(n_519),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_568),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_552),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_570),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

INVxp67_ASAP7_75t_SL g637 ( 
.A(n_561),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_R g638 ( 
.A(n_578),
.B(n_418),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_534),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_553),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_584),
.B(n_530),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_576),
.B(n_440),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_595),
.B(n_440),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_584),
.B(n_530),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_594),
.B(n_487),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_539),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_594),
.B(n_487),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_553),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_534),
.B(n_474),
.Y(n_649)
);

AND2x2_ASAP7_75t_SL g650 ( 
.A(n_536),
.B(n_438),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_567),
.Y(n_651)
);

BUFx4f_ASAP7_75t_SL g652 ( 
.A(n_567),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_534),
.B(n_476),
.Y(n_654)
);

AND2x6_ASAP7_75t_L g655 ( 
.A(n_585),
.B(n_412),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_589),
.B(n_440),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_557),
.B(n_489),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_589),
.B(n_440),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_571),
.B(n_476),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_562),
.B(n_412),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_542),
.B(n_477),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_542),
.B(n_592),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_574),
.B(n_440),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_532),
.B(n_440),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_547),
.A2(n_395),
.B(n_384),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_532),
.B(n_450),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_554),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_572),
.B(n_382),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_574),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_555),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_579),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_555),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_590),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_535),
.B(n_489),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_556),
.Y(n_675)
);

INVx3_ASAP7_75t_L g676 ( 
.A(n_556),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_535),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_596),
.B(n_394),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_533),
.B(n_496),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_563),
.B(n_394),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_547),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_563),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_538),
.B(n_450),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_618),
.B(n_537),
.Y(n_684)
);

NOR2xp67_ASAP7_75t_L g685 ( 
.A(n_671),
.B(n_581),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_662),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_619),
.B(n_543),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_618),
.Y(n_688)
);

INVx6_ASAP7_75t_L g689 ( 
.A(n_599),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_681),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_601),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_601),
.Y(n_693)
);

AND2x2_ASAP7_75t_SL g694 ( 
.A(n_650),
.B(n_587),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_618),
.Y(n_695)
);

NOR2xp67_ASAP7_75t_SL g696 ( 
.A(n_607),
.B(n_402),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_606),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_619),
.B(n_546),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_662),
.B(n_437),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_668),
.B(n_581),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_650),
.B(n_507),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_650),
.B(n_501),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_599),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_598),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_662),
.B(n_437),
.Y(n_705)
);

BUFx6f_ASAP7_75t_L g706 ( 
.A(n_599),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_677),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_662),
.B(n_637),
.Y(n_708)
);

AOI21x1_ASAP7_75t_L g709 ( 
.A1(n_664),
.A2(n_395),
.B(n_384),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_599),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_662),
.B(n_444),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_629),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_650),
.B(n_520),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_604),
.B(n_492),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_601),
.Y(n_715)
);

NOR2x1_ASAP7_75t_L g716 ( 
.A(n_639),
.B(n_541),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_637),
.B(n_444),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_604),
.B(n_494),
.Y(n_718)
);

INVx4_ASAP7_75t_L g719 ( 
.A(n_607),
.Y(n_719)
);

OR2x2_ASAP7_75t_L g720 ( 
.A(n_605),
.B(n_544),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_668),
.B(n_465),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_681),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_610),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_651),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_668),
.B(n_465),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_610),
.Y(n_726)
);

NAND2x1p5_ASAP7_75t_L g727 ( 
.A(n_607),
.B(n_427),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_678),
.B(n_434),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_633),
.B(n_441),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_633),
.B(n_442),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_SL g731 ( 
.A(n_598),
.B(n_567),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_629),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_677),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_677),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_671),
.B(n_646),
.Y(n_735)
);

INVx4_ASAP7_75t_L g736 ( 
.A(n_607),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_478),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_606),
.Y(n_738)
);

OR2x6_ASAP7_75t_L g739 ( 
.A(n_639),
.B(n_418),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_606),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_605),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_607),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_678),
.B(n_434),
.Y(n_743)
);

BUFx6f_ASAP7_75t_SL g744 ( 
.A(n_663),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_677),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_603),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_612),
.B(n_478),
.Y(n_747)
);

CKINVDCx11_ASAP7_75t_R g748 ( 
.A(n_646),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_613),
.Y(n_749)
);

BUFx2_ASAP7_75t_L g750 ( 
.A(n_605),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_658),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_678),
.B(n_635),
.Y(n_752)
);

AND2x2_ASAP7_75t_SL g753 ( 
.A(n_663),
.B(n_541),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_635),
.B(n_586),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_614),
.B(n_458),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_614),
.B(n_458),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_658),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_660),
.B(n_586),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_597),
.B(n_559),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_603),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_658),
.B(n_422),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_597),
.B(n_458),
.Y(n_762)
);

BUFx8_ASAP7_75t_L g763 ( 
.A(n_649),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_615),
.B(n_458),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_606),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_603),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_615),
.B(n_458),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_660),
.B(n_559),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_677),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_669),
.B(n_544),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_655),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_679),
.B(n_463),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_631),
.Y(n_773)
);

NAND2x1p5_ASAP7_75t_L g774 ( 
.A(n_658),
.B(n_427),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_613),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_676),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_679),
.B(n_608),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_603),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_638),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_638),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_651),
.Y(n_781)
);

BUFx2_ASAP7_75t_L g782 ( 
.A(n_741),
.Y(n_782)
);

BUFx2_ASAP7_75t_SL g783 ( 
.A(n_703),
.Y(n_783)
);

INVx5_ASAP7_75t_L g784 ( 
.A(n_751),
.Y(n_784)
);

BUFx4_ASAP7_75t_SL g785 ( 
.A(n_704),
.Y(n_785)
);

BUFx3_ASAP7_75t_L g786 ( 
.A(n_741),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_769),
.Y(n_787)
);

BUFx4f_ASAP7_75t_SL g788 ( 
.A(n_724),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_728),
.B(n_600),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_748),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_697),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_750),
.Y(n_792)
);

BUFx12f_ASAP7_75t_L g793 ( 
.A(n_748),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_732),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_697),
.Y(n_795)
);

BUFx2_ASAP7_75t_L g796 ( 
.A(n_750),
.Y(n_796)
);

INVx6_ASAP7_75t_L g797 ( 
.A(n_751),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_688),
.B(n_649),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_688),
.B(n_649),
.Y(n_799)
);

INVx3_ASAP7_75t_SL g800 ( 
.A(n_779),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_751),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_751),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_690),
.Y(n_803)
);

BUFx12f_ASAP7_75t_L g804 ( 
.A(n_724),
.Y(n_804)
);

CKINVDCx11_ASAP7_75t_R g805 ( 
.A(n_781),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_732),
.Y(n_806)
);

CKINVDCx16_ASAP7_75t_R g807 ( 
.A(n_704),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_722),
.Y(n_808)
);

BUFx2_ASAP7_75t_SL g809 ( 
.A(n_703),
.Y(n_809)
);

INVx1_ASAP7_75t_SL g810 ( 
.A(n_712),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_738),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_738),
.Y(n_812)
);

BUFx2_ASAP7_75t_SL g813 ( 
.A(n_703),
.Y(n_813)
);

INVx4_ASAP7_75t_L g814 ( 
.A(n_689),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_751),
.Y(n_815)
);

HB1xp67_ASAP7_75t_L g816 ( 
.A(n_752),
.Y(n_816)
);

BUFx12f_ASAP7_75t_L g817 ( 
.A(n_781),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_691),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_740),
.Y(n_819)
);

BUFx3_ASAP7_75t_L g820 ( 
.A(n_757),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_769),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_769),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_701),
.A2(n_669),
.B1(n_673),
.B2(n_600),
.Y(n_823)
);

BUFx4f_ASAP7_75t_L g824 ( 
.A(n_757),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_740),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_765),
.Y(n_826)
);

INVx2_ASAP7_75t_SL g827 ( 
.A(n_689),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_765),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_744),
.A2(n_673),
.B1(n_654),
.B2(n_608),
.Y(n_829)
);

NAND2x1p5_ASAP7_75t_L g830 ( 
.A(n_719),
.B(n_676),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_708),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_773),
.Y(n_832)
);

INVx4_ASAP7_75t_L g833 ( 
.A(n_689),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_728),
.B(n_654),
.Y(n_834)
);

INVx4_ASAP7_75t_L g835 ( 
.A(n_689),
.Y(n_835)
);

NOR2x1_ASAP7_75t_SL g836 ( 
.A(n_773),
.B(n_643),
.Y(n_836)
);

NAND2x1p5_ASAP7_75t_L g837 ( 
.A(n_719),
.B(n_676),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_691),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_723),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_757),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_708),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_757),
.Y(n_842)
);

BUFx3_ASAP7_75t_L g843 ( 
.A(n_757),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_763),
.Y(n_844)
);

INVx6_ASAP7_75t_L g845 ( 
.A(n_703),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_719),
.B(n_676),
.Y(n_846)
);

INVx1_ASAP7_75t_SL g847 ( 
.A(n_754),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_763),
.Y(n_848)
);

BUFx5_ASAP7_75t_L g849 ( 
.A(n_771),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_703),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_706),
.Y(n_851)
);

BUFx4f_ASAP7_75t_SL g852 ( 
.A(n_763),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_706),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_726),
.Y(n_854)
);

BUFx6f_ASAP7_75t_SL g855 ( 
.A(n_761),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_749),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_686),
.Y(n_857)
);

INVx8_ASAP7_75t_L g858 ( 
.A(n_744),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_736),
.B(n_676),
.Y(n_859)
);

INVx8_ASAP7_75t_L g860 ( 
.A(n_744),
.Y(n_860)
);

INVxp67_ASAP7_75t_SL g861 ( 
.A(n_706),
.Y(n_861)
);

INVx3_ASAP7_75t_SL g862 ( 
.A(n_779),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_775),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_692),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_713),
.A2(n_602),
.B1(n_663),
.B2(n_657),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_708),
.Y(n_867)
);

INVx2_ASAP7_75t_SL g868 ( 
.A(n_706),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_695),
.B(n_654),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_702),
.A2(n_602),
.B1(n_663),
.B2(n_657),
.Y(n_870)
);

BUFx12f_ASAP7_75t_L g871 ( 
.A(n_780),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_686),
.Y(n_872)
);

INVx4_ASAP7_75t_L g873 ( 
.A(n_710),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_752),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_692),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_780),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_866),
.A2(n_694),
.B1(n_777),
.B2(n_753),
.Y(n_877)
);

INVx6_ASAP7_75t_L g878 ( 
.A(n_784),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_870),
.A2(n_694),
.B1(n_753),
.B2(n_772),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_814),
.Y(n_880)
);

BUFx12f_ASAP7_75t_L g881 ( 
.A(n_805),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_803),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_808),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_834),
.A2(n_747),
.B1(n_737),
.B2(n_721),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_SL g885 ( 
.A1(n_852),
.A2(n_577),
.B1(n_565),
.B2(n_768),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_876),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_839),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_854),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_856),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_863),
.Y(n_890)
);

INVx1_ASAP7_75t_SL g891 ( 
.A(n_810),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

BUFx8_ASAP7_75t_L g893 ( 
.A(n_804),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_798),
.A2(n_721),
.B1(n_725),
.B2(n_718),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_791),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_831),
.A2(n_735),
.B1(n_695),
.B2(n_685),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_818),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_798),
.A2(n_725),
.B1(n_714),
.B2(n_500),
.Y(n_899)
);

CKINVDCx11_ASAP7_75t_R g900 ( 
.A(n_805),
.Y(n_900)
);

CKINVDCx11_ASAP7_75t_R g901 ( 
.A(n_793),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_814),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_791),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_799),
.A2(n_509),
.B1(n_674),
.B2(n_743),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_847),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_831),
.A2(n_776),
.B1(n_700),
.B2(n_771),
.Y(n_906)
);

INVx3_ASAP7_75t_SL g907 ( 
.A(n_800),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_844),
.A2(n_577),
.B1(n_565),
.B2(n_768),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_795),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_841),
.A2(n_867),
.B1(n_829),
.B2(n_824),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_799),
.A2(n_674),
.B1(n_743),
.B2(n_624),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_786),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_795),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_785),
.Y(n_914)
);

OAI22xp33_ASAP7_75t_L g915 ( 
.A1(n_789),
.A2(n_720),
.B1(n_770),
.B2(n_731),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_811),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_786),
.Y(n_917)
);

OR2x2_ASAP7_75t_L g918 ( 
.A(n_874),
.B(n_770),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_876),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_800),
.Y(n_920)
);

CKINVDCx11_ASAP7_75t_R g921 ( 
.A(n_793),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_838),
.Y(n_922)
);

OAI21xp33_ASAP7_75t_L g923 ( 
.A1(n_874),
.A2(n_700),
.B(n_759),
.Y(n_923)
);

OAI22xp33_ASAP7_75t_L g924 ( 
.A1(n_807),
.A2(n_720),
.B1(n_758),
.B2(n_716),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_869),
.B(n_684),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_792),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_811),
.Y(n_927)
);

INVx6_ASAP7_75t_L g928 ( 
.A(n_784),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_814),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_812),
.Y(n_930)
);

AOI22xp33_ASAP7_75t_L g931 ( 
.A1(n_869),
.A2(n_624),
.B1(n_684),
.B2(n_659),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_812),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_833),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_823),
.A2(n_659),
.B1(n_758),
.B2(n_687),
.Y(n_934)
);

OAI22xp33_ASAP7_75t_L g935 ( 
.A1(n_844),
.A2(n_754),
.B1(n_739),
.B2(n_652),
.Y(n_935)
);

OAI22xp33_ASAP7_75t_L g936 ( 
.A1(n_848),
.A2(n_739),
.B1(n_652),
.B2(n_761),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_858),
.A2(n_659),
.B1(n_608),
.B2(n_661),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_832),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_850),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_784),
.Y(n_940)
);

BUFx2_ASAP7_75t_L g941 ( 
.A(n_792),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_832),
.Y(n_942)
);

BUFx12f_ASAP7_75t_L g943 ( 
.A(n_804),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_858),
.A2(n_608),
.B1(n_661),
.B2(n_717),
.Y(n_944)
);

AOI22xp33_ASAP7_75t_L g945 ( 
.A1(n_858),
.A2(n_608),
.B1(n_661),
.B2(n_717),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_858),
.A2(n_608),
.B1(n_860),
.B2(n_717),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_838),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_860),
.A2(n_608),
.B1(n_730),
.B2(n_729),
.Y(n_948)
);

NAND2x1p5_ASAP7_75t_L g949 ( 
.A(n_784),
.B(n_710),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_SL g950 ( 
.A1(n_848),
.A2(n_680),
.B1(n_608),
.B2(n_656),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_SL g951 ( 
.A1(n_860),
.A2(n_680),
.B1(n_608),
.B2(n_656),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_819),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_782),
.B(n_680),
.Y(n_953)
);

BUFx8_ASAP7_75t_L g954 ( 
.A(n_855),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_841),
.A2(n_625),
.B1(n_733),
.B2(n_707),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_875),
.Y(n_956)
);

OAI22xp5_ASAP7_75t_SL g957 ( 
.A1(n_790),
.A2(n_682),
.B1(n_739),
.B2(n_761),
.Y(n_957)
);

INVx4_ASAP7_75t_L g958 ( 
.A(n_784),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_825),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_867),
.A2(n_824),
.B1(n_860),
.B2(n_835),
.Y(n_960)
);

CKINVDCx11_ASAP7_75t_R g961 ( 
.A(n_817),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_855),
.A2(n_608),
.B1(n_739),
.B2(n_480),
.Y(n_962)
);

CKINVDCx6p67_ASAP7_75t_R g963 ( 
.A(n_862),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_855),
.A2(n_729),
.B1(n_730),
.B2(n_660),
.Y(n_964)
);

BUFx12f_ASAP7_75t_L g965 ( 
.A(n_817),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_SL g966 ( 
.A1(n_788),
.A2(n_429),
.B1(n_453),
.B2(n_422),
.Y(n_966)
);

BUFx2_ASAP7_75t_SL g967 ( 
.A(n_794),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_824),
.A2(n_625),
.B1(n_733),
.B2(n_707),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_833),
.A2(n_835),
.B1(n_821),
.B2(n_822),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_782),
.B(n_699),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_796),
.Y(n_971)
);

OAI22xp5_ASAP7_75t_L g972 ( 
.A1(n_833),
.A2(n_733),
.B1(n_734),
.B2(n_707),
.Y(n_972)
);

BUFx8_ASAP7_75t_SL g973 ( 
.A(n_871),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_871),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_794),
.B(n_729),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_826),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_875),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_796),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_862),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_SL g980 ( 
.A1(n_806),
.A2(n_453),
.B1(n_429),
.B2(n_609),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_828),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_864),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_835),
.A2(n_734),
.B1(n_745),
.B2(n_710),
.Y(n_983)
);

BUFx4_ASAP7_75t_SL g984 ( 
.A(n_857),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_865),
.Y(n_985)
);

CKINVDCx20_ASAP7_75t_R g986 ( 
.A(n_857),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_934),
.A2(n_872),
.B1(n_761),
.B2(n_821),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_940),
.Y(n_989)
);

OAI21xp33_ASAP7_75t_L g990 ( 
.A1(n_934),
.A2(n_705),
.B(n_699),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_939),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_925),
.B(n_730),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_931),
.A2(n_872),
.B1(n_787),
.B2(n_822),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_900),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_931),
.A2(n_787),
.B1(n_822),
.B2(n_821),
.Y(n_995)
);

OAI21xp5_ASAP7_75t_SL g996 ( 
.A1(n_962),
.A2(n_682),
.B(n_609),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_964),
.A2(n_895),
.B1(n_884),
.B2(n_879),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_956),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_882),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_956),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_877),
.A2(n_705),
.B1(n_711),
.B2(n_699),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_915),
.A2(n_711),
.B1(n_705),
.B2(n_764),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_900),
.Y(n_1003)
);

OAI21xp5_ASAP7_75t_SL g1004 ( 
.A1(n_899),
.A2(n_609),
.B(n_622),
.Y(n_1004)
);

AOI22xp33_ASAP7_75t_SL g1005 ( 
.A1(n_957),
.A2(n_643),
.B1(n_626),
.B2(n_622),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_891),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_940),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_918),
.B(n_616),
.Y(n_1008)
);

NOR2x1p5_ASAP7_75t_L g1009 ( 
.A(n_963),
.B(n_820),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_923),
.A2(n_711),
.B1(n_767),
.B2(n_655),
.Y(n_1010)
);

AOI22xp33_ASAP7_75t_L g1011 ( 
.A1(n_924),
.A2(n_655),
.B1(n_840),
.B2(n_820),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_SL g1012 ( 
.A(n_943),
.Y(n_1012)
);

CKINVDCx20_ASAP7_75t_R g1013 ( 
.A(n_886),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_884),
.A2(n_655),
.B1(n_842),
.B2(n_840),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_895),
.A2(n_698),
.B(n_762),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_899),
.B(n_905),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_971),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_950),
.A2(n_655),
.B1(n_843),
.B2(n_842),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_SL g1019 ( 
.A1(n_954),
.A2(n_626),
.B1(n_622),
.B2(n_783),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_937),
.A2(n_655),
.B1(n_843),
.B2(n_450),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_937),
.A2(n_964),
.B1(n_908),
.B2(n_951),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_SL g1022 ( 
.A1(n_885),
.A2(n_626),
.B(n_616),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_897),
.B(n_787),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_SL g1024 ( 
.A1(n_954),
.A2(n_809),
.B1(n_813),
.B2(n_783),
.Y(n_1024)
);

AOI22xp33_ASAP7_75t_L g1025 ( 
.A1(n_953),
.A2(n_655),
.B1(n_450),
.B2(n_797),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_904),
.B(n_616),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_919),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_904),
.A2(n_837),
.B1(n_846),
.B2(n_830),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_896),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_970),
.B(n_630),
.Y(n_1030)
);

AOI222xp33_ASAP7_75t_L g1031 ( 
.A1(n_892),
.A2(n_454),
.B1(n_448),
.B2(n_442),
.C1(n_647),
.C2(n_645),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_935),
.A2(n_628),
.B1(n_621),
.B2(n_655),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_944),
.A2(n_837),
.B1(n_846),
.B2(n_830),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_939),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_911),
.A2(n_655),
.B1(n_450),
.B2(n_797),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_883),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_911),
.A2(n_655),
.B1(n_450),
.B2(n_797),
.Y(n_1037)
);

OAI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_920),
.A2(n_628),
.B1(n_621),
.B2(n_801),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_SL g1039 ( 
.A1(n_954),
.A2(n_809),
.B1(n_813),
.B2(n_849),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_944),
.A2(n_830),
.B1(n_846),
.B2(n_837),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_945),
.A2(n_859),
.B1(n_861),
.B2(n_710),
.Y(n_1041)
);

OAI21xp5_ASAP7_75t_SL g1042 ( 
.A1(n_966),
.A2(n_658),
.B(n_632),
.Y(n_1042)
);

NAND3xp33_ASAP7_75t_L g1043 ( 
.A(n_980),
.B(n_948),
.C(n_975),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_910),
.A2(n_450),
.B1(n_815),
.B2(n_797),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_960),
.B(n_850),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_887),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_SL g1047 ( 
.A1(n_920),
.A2(n_849),
.B1(n_836),
.B2(n_802),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_L g1048 ( 
.A1(n_948),
.A2(n_815),
.B1(n_617),
.B2(n_667),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_888),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_986),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_971),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_889),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_945),
.A2(n_815),
.B1(n_617),
.B2(n_667),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_890),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_978),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_952),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_SL g1057 ( 
.A1(n_967),
.A2(n_849),
.B1(n_836),
.B2(n_802),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_973),
.Y(n_1058)
);

OAI21xp5_ASAP7_75t_SL g1059 ( 
.A1(n_936),
.A2(n_632),
.B(n_630),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_958),
.Y(n_1060)
);

BUFx4f_ASAP7_75t_SL g1061 ( 
.A(n_943),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_906),
.A2(n_978),
.B1(n_917),
.B2(n_941),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_955),
.A2(n_756),
.B(n_755),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_973),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_977),
.B(n_853),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_959),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_907),
.A2(n_815),
.B1(n_617),
.B2(n_648),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_977),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_976),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_894),
.B(n_853),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_981),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_SL g1072 ( 
.A1(n_903),
.A2(n_742),
.B(n_736),
.Y(n_1072)
);

OAI21xp33_ASAP7_75t_L g1073 ( 
.A1(n_912),
.A2(n_632),
.B(n_630),
.Y(n_1073)
);

AOI22xp33_ASAP7_75t_L g1074 ( 
.A1(n_907),
.A2(n_617),
.B1(n_672),
.B2(n_648),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_909),
.Y(n_1075)
);

BUFx12f_ASAP7_75t_L g1076 ( 
.A(n_961),
.Y(n_1076)
);

OAI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_979),
.A2(n_621),
.B1(n_628),
.B2(n_801),
.Y(n_1077)
);

BUFx4f_ASAP7_75t_SL g1078 ( 
.A(n_965),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_894),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_946),
.A2(n_859),
.B1(n_710),
.B2(n_745),
.Y(n_1080)
);

AOI22xp33_ASAP7_75t_L g1081 ( 
.A1(n_997),
.A2(n_974),
.B1(n_881),
.B2(n_921),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_1043),
.A2(n_974),
.B1(n_881),
.B2(n_921),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_1051),
.Y(n_1083)
);

AOI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_996),
.A2(n_965),
.B1(n_987),
.B2(n_946),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1021),
.A2(n_990),
.B1(n_1005),
.B2(n_1016),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1026),
.A2(n_901),
.B1(n_987),
.B2(n_926),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_1008),
.A2(n_901),
.B1(n_926),
.B2(n_912),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_SL g1088 ( 
.A1(n_1028),
.A2(n_893),
.B1(n_928),
.B2(n_878),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_SL g1089 ( 
.A1(n_988),
.A2(n_893),
.B1(n_928),
.B2(n_878),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1006),
.B(n_982),
.Y(n_1090)
);

OAI222xp33_ASAP7_75t_L g1091 ( 
.A1(n_1019),
.A2(n_252),
.B1(n_254),
.B2(n_258),
.C1(n_930),
.C2(n_942),
.Y(n_1091)
);

OAI221xp5_ASAP7_75t_L g1092 ( 
.A1(n_1042),
.A2(n_454),
.B1(n_448),
.B2(n_628),
.C(n_621),
.Y(n_1092)
);

AOI221xp5_ASAP7_75t_L g1093 ( 
.A1(n_1004),
.A2(n_647),
.B1(n_645),
.B2(n_644),
.C(n_641),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_998),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1011),
.A2(n_961),
.B1(n_627),
.B2(n_636),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_992),
.B(n_913),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1002),
.A2(n_627),
.B1(n_636),
.B2(n_620),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1029),
.B(n_916),
.Y(n_1098)
);

OAI22x1_ASAP7_75t_L g1099 ( 
.A1(n_1051),
.A2(n_932),
.B1(n_938),
.B2(n_927),
.Y(n_1099)
);

OAI221xp5_ASAP7_75t_SL g1100 ( 
.A1(n_1022),
.A2(n_644),
.B1(n_641),
.B2(n_647),
.C(n_645),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_SL g1101 ( 
.A1(n_1041),
.A2(n_949),
.B(n_958),
.Y(n_1101)
);

AOI222xp33_ASAP7_75t_L g1102 ( 
.A1(n_1059),
.A2(n_391),
.B1(n_401),
.B2(n_420),
.C1(n_644),
.C2(n_641),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1030),
.B(n_898),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1029),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_SL g1105 ( 
.A1(n_1076),
.A2(n_928),
.B1(n_878),
.B2(n_914),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1001),
.A2(n_672),
.B1(n_620),
.B2(n_802),
.Y(n_1106)
);

OAI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1032),
.A2(n_880),
.B1(n_902),
.B2(n_929),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1050),
.A2(n_1074),
.B1(n_1010),
.B2(n_1014),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1050),
.A2(n_801),
.B1(n_802),
.B2(n_381),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_L g1110 ( 
.A1(n_1018),
.A2(n_801),
.B1(n_802),
.B2(n_381),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1073),
.A2(n_801),
.B1(n_381),
.B2(n_968),
.Y(n_1111)
);

OAI21xp5_ASAP7_75t_SL g1112 ( 
.A1(n_1044),
.A2(n_642),
.B(n_401),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_998),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1076),
.A2(n_381),
.B1(n_849),
.B2(n_827),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1000),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1031),
.A2(n_258),
.B1(n_274),
.B2(n_318),
.Y(n_1116)
);

AOI22xp33_ASAP7_75t_L g1117 ( 
.A1(n_1062),
.A2(n_381),
.B1(n_849),
.B2(n_827),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1067),
.A2(n_1048),
.B1(n_1053),
.B2(n_1017),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1000),
.Y(n_1119)
);

OAI222xp33_ASAP7_75t_L g1120 ( 
.A1(n_1077),
.A2(n_898),
.B1(n_922),
.B2(n_947),
.C1(n_304),
.C2(n_272),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1038),
.B(n_880),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_L g1122 ( 
.A(n_1015),
.B(n_420),
.C(n_391),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1055),
.A2(n_381),
.B1(n_849),
.B2(n_845),
.Y(n_1123)
);

HB1xp67_ASAP7_75t_L g1124 ( 
.A(n_1065),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_1023),
.A2(n_1061),
.B1(n_1078),
.B2(n_1012),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1023),
.A2(n_1027),
.B1(n_1013),
.B2(n_1045),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_SL g1127 ( 
.A1(n_1013),
.A2(n_969),
.B1(n_929),
.B2(n_902),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1027),
.A2(n_933),
.B1(n_859),
.B2(n_985),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1045),
.A2(n_381),
.B1(n_849),
.B2(n_845),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1068),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1045),
.A2(n_849),
.B1(n_845),
.B2(n_933),
.Y(n_1131)
);

AOI222xp33_ASAP7_75t_L g1132 ( 
.A1(n_999),
.A2(n_419),
.B1(n_623),
.B2(n_611),
.C1(n_262),
.C2(n_347),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1045),
.A2(n_845),
.B1(n_865),
.B2(n_873),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1033),
.A2(n_1040),
.B1(n_993),
.B2(n_1009),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1063),
.A2(n_665),
.B(n_709),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1039),
.A2(n_985),
.B1(n_949),
.B2(n_734),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1036),
.B(n_922),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1046),
.A2(n_865),
.B1(n_873),
.B2(n_868),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1049),
.A2(n_873),
.B1(n_868),
.B2(n_851),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1052),
.A2(n_947),
.B1(n_611),
.B2(n_623),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1054),
.A2(n_1020),
.B1(n_1056),
.B2(n_1066),
.Y(n_1141)
);

OA21x2_ASAP7_75t_L g1142 ( 
.A1(n_1075),
.A2(n_665),
.B(n_709),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_994),
.A2(n_972),
.B1(n_939),
.B2(n_850),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1069),
.B(n_939),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_1071),
.A2(n_850),
.B1(n_851),
.B2(n_634),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_SL g1146 ( 
.A1(n_994),
.A2(n_850),
.B1(n_851),
.B2(n_983),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1084),
.B(n_1125),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1124),
.B(n_1068),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1092),
.A2(n_1118),
.B1(n_1122),
.B2(n_1128),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1104),
.B(n_1065),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1090),
.B(n_1070),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1082),
.B(n_1003),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1104),
.B(n_1070),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1096),
.B(n_1079),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1098),
.B(n_1079),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_SL g1156 ( 
.A1(n_1081),
.A2(n_1024),
.B(n_1047),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1132),
.B(n_1037),
.C(n_1035),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1087),
.B(n_1003),
.Y(n_1158)
);

AOI22xp33_ASAP7_75t_L g1159 ( 
.A1(n_1085),
.A2(n_1057),
.B1(n_1025),
.B2(n_419),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1126),
.A2(n_419),
.B1(n_1058),
.B2(n_1064),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1098),
.B(n_991),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1083),
.B(n_991),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1083),
.B(n_991),
.Y(n_1163)
);

NAND2xp33_ASAP7_75t_L g1164 ( 
.A(n_1084),
.B(n_851),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1091),
.A2(n_1007),
.B(n_989),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_1088),
.B(n_989),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_1116),
.A2(n_261),
.B1(n_265),
.B2(n_312),
.C(n_266),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1103),
.B(n_991),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1113),
.B(n_991),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1137),
.B(n_1034),
.Y(n_1170)
);

OAI221xp5_ASAP7_75t_L g1171 ( 
.A1(n_1086),
.A2(n_1058),
.B1(n_1064),
.B2(n_283),
.C(n_291),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1144),
.B(n_1034),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_L g1173 ( 
.A(n_1132),
.B(n_269),
.C(n_268),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1102),
.A2(n_995),
.B1(n_1080),
.B2(n_1072),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1113),
.B(n_1034),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1115),
.B(n_1034),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_L g1177 ( 
.A(n_1116),
.B(n_271),
.C(n_270),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_L g1178 ( 
.A(n_1102),
.B(n_279),
.C(n_276),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1089),
.A2(n_1060),
.B1(n_1007),
.B2(n_989),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_1134),
.A2(n_1060),
.B(n_1007),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_1141),
.B(n_293),
.C(n_282),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1115),
.B(n_1034),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1122),
.B(n_295),
.C(n_297),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1130),
.B(n_1060),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1130),
.B(n_46),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1120),
.B(n_984),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1094),
.B(n_303),
.Y(n_1187)
);

OA21x2_ASAP7_75t_L g1188 ( 
.A1(n_1094),
.A2(n_665),
.B(n_631),
.Y(n_1188)
);

AND2x2_ASAP7_75t_SL g1189 ( 
.A(n_1131),
.B(n_1129),
.Y(n_1189)
);

NAND2xp33_ASAP7_75t_SL g1190 ( 
.A(n_1121),
.B(n_851),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1119),
.B(n_46),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1119),
.B(n_306),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1099),
.B(n_47),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1099),
.B(n_310),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_L g1195 ( 
.A(n_1108),
.B(n_326),
.C(n_329),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1146),
.B(n_47),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1127),
.B(n_49),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1107),
.B(n_330),
.Y(n_1198)
);

NAND3xp33_ASAP7_75t_L g1199 ( 
.A(n_1173),
.B(n_1177),
.C(n_1181),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1150),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_L g1201 ( 
.A(n_1173),
.B(n_1105),
.C(n_1100),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1150),
.B(n_1143),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_SL g1203 ( 
.A1(n_1186),
.A2(n_1136),
.B1(n_1140),
.B2(n_1101),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1153),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1177),
.B(n_1112),
.C(n_1140),
.Y(n_1205)
);

OA211x2_ASAP7_75t_L g1206 ( 
.A1(n_1147),
.A2(n_1139),
.B(n_1117),
.C(n_1111),
.Y(n_1206)
);

NAND4xp75_ASAP7_75t_L g1207 ( 
.A(n_1197),
.B(n_1093),
.C(n_51),
.D(n_52),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1169),
.B(n_1135),
.Y(n_1208)
);

OR2x2_ASAP7_75t_L g1209 ( 
.A(n_1161),
.B(n_1135),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_SL g1210 ( 
.A(n_1149),
.B(n_1194),
.Y(n_1210)
);

XNOR2xp5_ASAP7_75t_L g1211 ( 
.A(n_1197),
.B(n_49),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1152),
.B(n_51),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1153),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1151),
.B(n_1135),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1148),
.Y(n_1215)
);

NOR3xp33_ASAP7_75t_L g1216 ( 
.A(n_1195),
.B(n_1112),
.C(n_331),
.Y(n_1216)
);

AOI211xp5_ASAP7_75t_L g1217 ( 
.A1(n_1165),
.A2(n_1101),
.B(n_335),
.C(n_443),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1169),
.B(n_1135),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_1158),
.B(n_53),
.Y(n_1219)
);

CKINVDCx20_ASAP7_75t_R g1220 ( 
.A(n_1172),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1155),
.B(n_1142),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1175),
.B(n_1133),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1175),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1184),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1184),
.B(n_1138),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1193),
.B(n_1145),
.Y(n_1226)
);

AO21x2_ASAP7_75t_L g1227 ( 
.A1(n_1181),
.A2(n_631),
.B(n_634),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1178),
.A2(n_1095),
.B1(n_1106),
.B2(n_1097),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_1176),
.Y(n_1229)
);

NAND4xp75_ASAP7_75t_L g1230 ( 
.A(n_1196),
.B(n_53),
.C(n_54),
.D(n_55),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1180),
.B(n_1142),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1193),
.B(n_1142),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_SL g1233 ( 
.A(n_1166),
.B(n_1114),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1195),
.B(n_1109),
.C(n_1123),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1178),
.A2(n_1110),
.B1(n_670),
.B2(n_640),
.Y(n_1235)
);

AOI221xp5_ASAP7_75t_L g1236 ( 
.A1(n_1196),
.A2(n_457),
.B1(n_456),
.B2(n_445),
.C(n_443),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1162),
.B(n_1142),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1182),
.Y(n_1238)
);

NAND3xp33_ASAP7_75t_L g1239 ( 
.A(n_1167),
.B(n_457),
.C(n_456),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1164),
.A2(n_670),
.B(n_634),
.Y(n_1240)
);

AO21x2_ASAP7_75t_L g1241 ( 
.A1(n_1164),
.A2(n_670),
.B(n_634),
.Y(n_1241)
);

NAND3xp33_ASAP7_75t_L g1242 ( 
.A(n_1198),
.B(n_457),
.C(n_432),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1157),
.B(n_457),
.C(n_432),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

NAND4xp75_ASAP7_75t_L g1245 ( 
.A(n_1189),
.B(n_54),
.C(n_57),
.D(n_59),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1168),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1163),
.B(n_61),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1185),
.B(n_1191),
.Y(n_1248)
);

NOR3xp33_ASAP7_75t_L g1249 ( 
.A(n_1171),
.B(n_675),
.C(n_631),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1185),
.B(n_61),
.Y(n_1250)
);

NAND4xp75_ASAP7_75t_L g1251 ( 
.A(n_1189),
.B(n_62),
.C(n_63),
.D(n_64),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1154),
.Y(n_1252)
);

INVx2_ASAP7_75t_SL g1253 ( 
.A(n_1191),
.Y(n_1253)
);

NAND2x1_ASAP7_75t_L g1254 ( 
.A(n_1174),
.B(n_736),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1252),
.B(n_1174),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1215),
.B(n_1189),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1246),
.B(n_1244),
.Y(n_1257)
);

INVx3_ASAP7_75t_L g1258 ( 
.A(n_1224),
.Y(n_1258)
);

NAND4xp75_ASAP7_75t_L g1259 ( 
.A(n_1210),
.B(n_1192),
.C(n_1187),
.D(n_1157),
.Y(n_1259)
);

HB1xp67_ASAP7_75t_L g1260 ( 
.A(n_1229),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1200),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1208),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1200),
.Y(n_1263)
);

NOR3xp33_ASAP7_75t_L g1264 ( 
.A(n_1199),
.B(n_1156),
.C(n_1183),
.Y(n_1264)
);

INVx2_ASAP7_75t_SL g1265 ( 
.A(n_1224),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1223),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1204),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1213),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1253),
.B(n_1179),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1223),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1237),
.B(n_1190),
.Y(n_1271)
);

NAND4xp75_ASAP7_75t_SL g1272 ( 
.A(n_1212),
.B(n_1188),
.C(n_696),
.D(n_1160),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1232),
.B(n_1188),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1208),
.Y(n_1274)
);

NOR4xp75_ASAP7_75t_L g1275 ( 
.A(n_1245),
.B(n_62),
.C(n_63),
.D(n_65),
.Y(n_1275)
);

INVx1_ASAP7_75t_SL g1276 ( 
.A(n_1220),
.Y(n_1276)
);

NAND4xp75_ASAP7_75t_SL g1277 ( 
.A(n_1219),
.B(n_1232),
.C(n_1217),
.D(n_1247),
.Y(n_1277)
);

NAND4xp75_ASAP7_75t_SL g1278 ( 
.A(n_1247),
.B(n_1188),
.C(n_696),
.D(n_1159),
.Y(n_1278)
);

XOR2x2_ASAP7_75t_L g1279 ( 
.A(n_1211),
.B(n_1183),
.Y(n_1279)
);

NOR4xp25_ASAP7_75t_L g1280 ( 
.A(n_1243),
.B(n_66),
.C(n_67),
.D(n_68),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1253),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1218),
.B(n_1188),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_SL g1283 ( 
.A(n_1205),
.B(n_1201),
.C(n_1203),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1237),
.B(n_66),
.Y(n_1284)
);

NAND4xp25_ASAP7_75t_L g1285 ( 
.A(n_1228),
.B(n_68),
.C(n_69),
.D(n_70),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1218),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1221),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1258),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1261),
.Y(n_1289)
);

XOR2x2_ASAP7_75t_L g1290 ( 
.A(n_1279),
.B(n_1283),
.Y(n_1290)
);

XNOR2xp5_ASAP7_75t_L g1291 ( 
.A(n_1279),
.B(n_1211),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1256),
.B(n_1284),
.Y(n_1292)
);

XNOR2xp5_ASAP7_75t_L g1293 ( 
.A(n_1279),
.B(n_1245),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1261),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_1276),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1256),
.B(n_1238),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1263),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1263),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1284),
.Y(n_1299)
);

INVxp67_ASAP7_75t_SL g1300 ( 
.A(n_1260),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1267),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1269),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1267),
.Y(n_1303)
);

AND2x4_ASAP7_75t_L g1304 ( 
.A(n_1262),
.B(n_1274),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_R g1305 ( 
.A(n_1277),
.B(n_1233),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1268),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1257),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1258),
.Y(n_1308)
);

XNOR2xp5_ASAP7_75t_L g1309 ( 
.A(n_1285),
.B(n_1251),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1287),
.B(n_1214),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1276),
.Y(n_1311)
);

XOR2x2_ASAP7_75t_L g1312 ( 
.A(n_1259),
.B(n_1251),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1281),
.Y(n_1313)
);

OAI22x1_ASAP7_75t_L g1314 ( 
.A1(n_1270),
.A2(n_1250),
.B1(n_1248),
.B2(n_1238),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1258),
.Y(n_1315)
);

XNOR2x2_ASAP7_75t_L g1316 ( 
.A(n_1275),
.B(n_1230),
.Y(n_1316)
);

XOR2x2_ASAP7_75t_L g1317 ( 
.A(n_1259),
.B(n_1230),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1271),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1255),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1293),
.A2(n_1309),
.B1(n_1291),
.B2(n_1319),
.Y(n_1320)
);

INVx3_ASAP7_75t_L g1321 ( 
.A(n_1304),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1301),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1313),
.Y(n_1323)
);

XOR2x2_ASAP7_75t_L g1324 ( 
.A(n_1290),
.B(n_1264),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1303),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1304),
.Y(n_1326)
);

AO22x1_ASAP7_75t_L g1327 ( 
.A1(n_1300),
.A2(n_1250),
.B1(n_1275),
.B2(n_1271),
.Y(n_1327)
);

OAI22x1_ASAP7_75t_SL g1328 ( 
.A1(n_1290),
.A2(n_1220),
.B1(n_1285),
.B2(n_1287),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1313),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1306),
.Y(n_1330)
);

AOI22x1_ASAP7_75t_SL g1331 ( 
.A1(n_1295),
.A2(n_1286),
.B1(n_1262),
.B2(n_1274),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1293),
.A2(n_1255),
.B1(n_1207),
.B2(n_1231),
.Y(n_1332)
);

XNOR2x1_ASAP7_75t_L g1333 ( 
.A(n_1291),
.B(n_1207),
.Y(n_1333)
);

AOI22x1_ASAP7_75t_L g1334 ( 
.A1(n_1309),
.A2(n_1248),
.B1(n_1226),
.B2(n_1202),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1304),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1295),
.A2(n_1280),
.B1(n_1254),
.B2(n_1231),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1319),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1307),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1289),
.Y(n_1339)
);

OA22x2_ASAP7_75t_L g1340 ( 
.A1(n_1311),
.A2(n_1270),
.B1(n_1231),
.B2(n_1265),
.Y(n_1340)
);

XNOR2x2_ASAP7_75t_L g1341 ( 
.A(n_1317),
.B(n_1239),
.Y(n_1341)
);

XNOR2x1_ASAP7_75t_L g1342 ( 
.A(n_1317),
.B(n_1272),
.Y(n_1342)
);

AO22x1_ASAP7_75t_L g1343 ( 
.A1(n_1312),
.A2(n_1216),
.B1(n_1202),
.B2(n_1249),
.Y(n_1343)
);

XOR2x2_ASAP7_75t_L g1344 ( 
.A(n_1312),
.B(n_1278),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1288),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1294),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1302),
.A2(n_1231),
.B1(n_1254),
.B2(n_1226),
.Y(n_1347)
);

INVx1_ASAP7_75t_SL g1348 ( 
.A(n_1307),
.Y(n_1348)
);

AOI22x1_ASAP7_75t_SL g1349 ( 
.A1(n_1318),
.A2(n_1305),
.B1(n_1316),
.B2(n_1297),
.Y(n_1349)
);

INVx2_ASAP7_75t_SL g1350 ( 
.A(n_1314),
.Y(n_1350)
);

AOI22x1_ASAP7_75t_L g1351 ( 
.A1(n_1314),
.A2(n_1273),
.B1(n_1262),
.B2(n_1274),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1299),
.A2(n_1234),
.B1(n_1242),
.B2(n_1214),
.Y(n_1352)
);

XNOR2x1_ASAP7_75t_L g1353 ( 
.A(n_1316),
.B(n_1206),
.Y(n_1353)
);

INVx5_ASAP7_75t_SL g1354 ( 
.A(n_1341),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1346),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1337),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1346),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1322),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1321),
.Y(n_1359)
);

OA22x2_ASAP7_75t_L g1360 ( 
.A1(n_1320),
.A2(n_1292),
.B1(n_1296),
.B2(n_1298),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1338),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1339),
.Y(n_1362)
);

XOR2x2_ASAP7_75t_L g1363 ( 
.A(n_1324),
.B(n_1236),
.Y(n_1363)
);

INVx2_ASAP7_75t_SL g1364 ( 
.A(n_1323),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1325),
.Y(n_1365)
);

INVx2_ASAP7_75t_SL g1366 ( 
.A(n_1323),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1330),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1329),
.Y(n_1368)
);

INVxp67_ASAP7_75t_SL g1369 ( 
.A(n_1328),
.Y(n_1369)
);

OAI322xp33_ASAP7_75t_L g1370 ( 
.A1(n_1333),
.A2(n_1310),
.A3(n_1209),
.B1(n_1268),
.B2(n_1286),
.C1(n_1221),
.C2(n_1315),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1329),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1348),
.Y(n_1372)
);

INVxp67_ASAP7_75t_L g1373 ( 
.A(n_1349),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1326),
.Y(n_1374)
);

NOR2x1_ASAP7_75t_SL g1375 ( 
.A(n_1350),
.B(n_1240),
.Y(n_1375)
);

BUFx2_ASAP7_75t_L g1376 ( 
.A(n_1350),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1324),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1326),
.Y(n_1378)
);

INVx1_ASAP7_75t_SL g1379 ( 
.A(n_1333),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1321),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1335),
.Y(n_1381)
);

INVxp67_ASAP7_75t_SL g1382 ( 
.A(n_1334),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1321),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1335),
.Y(n_1384)
);

AOI322xp5_ASAP7_75t_L g1385 ( 
.A1(n_1341),
.A2(n_1273),
.A3(n_1286),
.B1(n_1282),
.B2(n_1265),
.C1(n_1266),
.C2(n_1222),
.Y(n_1385)
);

AOI22x1_ASAP7_75t_L g1386 ( 
.A1(n_1377),
.A2(n_1353),
.B1(n_1344),
.B2(n_1342),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1361),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1361),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1369),
.A2(n_1336),
.B1(n_1344),
.B2(n_1342),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1362),
.Y(n_1390)
);

AOI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1354),
.A2(n_1332),
.B1(n_1353),
.B2(n_1343),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1354),
.A2(n_1327),
.B1(n_1347),
.B2(n_1352),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1354),
.A2(n_1331),
.B1(n_1340),
.B2(n_1280),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1362),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1365),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1365),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1377),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1355),
.Y(n_1398)
);

INVxp67_ASAP7_75t_SL g1399 ( 
.A(n_1356),
.Y(n_1399)
);

BUFx4_ASAP7_75t_R g1400 ( 
.A(n_1354),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1373),
.A2(n_1340),
.B1(n_1345),
.B2(n_1351),
.Y(n_1401)
);

OA22x2_ASAP7_75t_L g1402 ( 
.A1(n_1379),
.A2(n_1382),
.B1(n_1372),
.B2(n_1376),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1357),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1376),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1358),
.Y(n_1405)
);

INVx1_ASAP7_75t_SL g1406 ( 
.A(n_1364),
.Y(n_1406)
);

AOI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1363),
.A2(n_1225),
.B1(n_1222),
.B2(n_1345),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1367),
.Y(n_1408)
);

OA22x2_ASAP7_75t_L g1409 ( 
.A1(n_1368),
.A2(n_1315),
.B1(n_1308),
.B2(n_1288),
.Y(n_1409)
);

OAI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1360),
.A2(n_1310),
.B1(n_1209),
.B2(n_1308),
.Y(n_1410)
);

NAND4xp25_ASAP7_75t_L g1411 ( 
.A(n_1385),
.B(n_1235),
.C(n_1225),
.D(n_71),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1378),
.Y(n_1412)
);

AOI22x1_ASAP7_75t_L g1413 ( 
.A1(n_1364),
.A2(n_1282),
.B1(n_1258),
.B2(n_71),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1366),
.Y(n_1414)
);

AOI22x1_ASAP7_75t_L g1415 ( 
.A1(n_1366),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_1415)
);

NAND4xp25_ASAP7_75t_L g1416 ( 
.A(n_1363),
.B(n_73),
.C(n_378),
.D(n_1227),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1397),
.A2(n_1370),
.B(n_1371),
.C(n_1360),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1391),
.A2(n_1360),
.B1(n_1381),
.B2(n_1374),
.Y(n_1418)
);

AO22x2_ASAP7_75t_L g1419 ( 
.A1(n_1404),
.A2(n_1383),
.B1(n_1380),
.B2(n_1359),
.Y(n_1419)
);

OAI31xp33_ASAP7_75t_L g1420 ( 
.A1(n_1411),
.A2(n_1384),
.A3(n_1378),
.B(n_1380),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1387),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1388),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1399),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_SL g1424 ( 
.A1(n_1389),
.A2(n_1383),
.B(n_1359),
.C(n_1384),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1392),
.A2(n_1375),
.B1(n_73),
.B2(n_1241),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1400),
.Y(n_1426)
);

AND4x1_ASAP7_75t_L g1427 ( 
.A(n_1393),
.B(n_1375),
.C(n_94),
.D(n_95),
.Y(n_1427)
);

OAI211xp5_ASAP7_75t_L g1428 ( 
.A1(n_1386),
.A2(n_443),
.B(n_432),
.C(n_445),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1412),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1406),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1411),
.A2(n_1241),
.B1(n_1240),
.B2(n_1227),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1402),
.A2(n_1241),
.B1(n_1240),
.B2(n_1227),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1406),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1414),
.Y(n_1434)
);

AO22x2_ASAP7_75t_L g1435 ( 
.A1(n_1398),
.A2(n_378),
.B1(n_640),
.B2(n_653),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1415),
.Y(n_1436)
);

INVxp67_ASAP7_75t_L g1437 ( 
.A(n_1413),
.Y(n_1437)
);

OA22x2_ASAP7_75t_L g1438 ( 
.A1(n_1407),
.A2(n_378),
.B1(n_640),
.B2(n_653),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_SL g1439 ( 
.A(n_1416),
.B(n_742),
.Y(n_1439)
);

OAI211xp5_ASAP7_75t_L g1440 ( 
.A1(n_1416),
.A2(n_432),
.B(n_443),
.C(n_457),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1401),
.A2(n_445),
.B1(n_456),
.B2(n_443),
.Y(n_1441)
);

INVxp33_ASAP7_75t_SL g1442 ( 
.A(n_1403),
.Y(n_1442)
);

AND4x1_ASAP7_75t_L g1443 ( 
.A(n_1390),
.B(n_92),
.C(n_96),
.D(n_97),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1405),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1394),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1410),
.A2(n_432),
.B1(n_445),
.B2(n_456),
.Y(n_1446)
);

AOI22x1_ASAP7_75t_L g1447 ( 
.A1(n_1408),
.A2(n_390),
.B1(n_404),
.B2(n_417),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1409),
.A2(n_445),
.B1(n_456),
.B2(n_675),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_L g1449 ( 
.A1(n_1395),
.A2(n_390),
.B1(n_404),
.B2(n_417),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1396),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1391),
.A2(n_390),
.B1(n_404),
.B2(n_417),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1391),
.A2(n_640),
.B1(n_653),
.B2(n_670),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1391),
.A2(n_390),
.B1(n_404),
.B2(n_417),
.Y(n_1453)
);

OAI211xp5_ASAP7_75t_L g1454 ( 
.A1(n_1391),
.A2(n_390),
.B(n_404),
.C(n_417),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1436),
.B(n_98),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1419),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1419),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1423),
.Y(n_1458)
);

OA22x2_ASAP7_75t_L g1459 ( 
.A1(n_1431),
.A2(n_653),
.B1(n_675),
.B2(n_642),
.Y(n_1459)
);

NOR4xp25_ASAP7_75t_L g1460 ( 
.A(n_1418),
.B(n_675),
.C(n_664),
.D(n_666),
.Y(n_1460)
);

NOR4xp25_ASAP7_75t_L g1461 ( 
.A(n_1417),
.B(n_666),
.C(n_766),
.D(n_760),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1421),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1426),
.Y(n_1463)
);

INVxp67_ASAP7_75t_SL g1464 ( 
.A(n_1437),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1425),
.A2(n_642),
.B1(n_693),
.B2(n_766),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1430),
.B(n_1433),
.Y(n_1466)
);

AO22x2_ASAP7_75t_L g1467 ( 
.A1(n_1422),
.A2(n_99),
.B1(n_101),
.B2(n_103),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1420),
.B(n_104),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1441),
.A2(n_745),
.B1(n_715),
.B2(n_760),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1429),
.Y(n_1470)
);

AO22x2_ASAP7_75t_L g1471 ( 
.A1(n_1445),
.A2(n_106),
.B1(n_112),
.B2(n_115),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1434),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1439),
.A2(n_642),
.B1(n_693),
.B2(n_746),
.Y(n_1473)
);

AOI221xp5_ASAP7_75t_L g1474 ( 
.A1(n_1424),
.A2(n_642),
.B1(n_683),
.B2(n_118),
.C(n_119),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1442),
.A2(n_683),
.B1(n_117),
.B2(n_122),
.C(n_123),
.Y(n_1475)
);

NOR2x1_ASAP7_75t_L g1476 ( 
.A(n_1428),
.B(n_742),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1450),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1444),
.B(n_1452),
.Y(n_1478)
);

AOI221xp5_ASAP7_75t_L g1479 ( 
.A1(n_1451),
.A2(n_683),
.B1(n_124),
.B2(n_127),
.C(n_130),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1435),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1453),
.A2(n_683),
.B1(n_131),
.B2(n_136),
.C(n_141),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1435),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1438),
.Y(n_1483)
);

AOI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1440),
.A2(n_778),
.B1(n_715),
.B2(n_746),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1446),
.A2(n_778),
.B1(n_774),
.B2(n_683),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1449),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1427),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1454),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1448),
.Y(n_1489)
);

NOR2x1_ASAP7_75t_L g1490 ( 
.A(n_1427),
.B(n_116),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1490),
.A2(n_1432),
.B1(n_1443),
.B2(n_1447),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1466),
.Y(n_1492)
);

AOI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1487),
.A2(n_1443),
.B1(n_774),
.B2(n_415),
.Y(n_1493)
);

AOI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1474),
.A2(n_774),
.B1(n_727),
.B2(n_415),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1472),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1464),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1463),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1456),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1457),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1462),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1467),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1461),
.A2(n_1468),
.B1(n_1458),
.B2(n_1465),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1482),
.Y(n_1503)
);

NOR2xp67_ASAP7_75t_L g1504 ( 
.A(n_1470),
.B(n_1477),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1467),
.Y(n_1505)
);

NOR2xp67_ASAP7_75t_L g1506 ( 
.A(n_1480),
.B(n_144),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1471),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1482),
.Y(n_1508)
);

AOI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1455),
.A2(n_415),
.B1(n_409),
.B2(n_402),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1483),
.A2(n_727),
.B1(n_415),
.B2(n_409),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1486),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1478),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1488),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1476),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1489),
.A2(n_727),
.B1(n_415),
.B2(n_409),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1459),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1460),
.B(n_1473),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1471),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1469),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1485),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1484),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1479),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1481),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1496),
.Y(n_1524)
);

NOR2xp67_ASAP7_75t_L g1525 ( 
.A(n_1497),
.B(n_146),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1498),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1499),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1495),
.Y(n_1528)
);

INVx1_ASAP7_75t_SL g1529 ( 
.A(n_1501),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1522),
.A2(n_1475),
.B1(n_415),
.B2(n_409),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1503),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1504),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1492),
.B(n_149),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1505),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1493),
.A2(n_1491),
.B1(n_1518),
.B2(n_1512),
.Y(n_1536)
);

AO211x2_ASAP7_75t_L g1537 ( 
.A1(n_1523),
.A2(n_153),
.B(n_155),
.C(n_156),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_158),
.Y(n_1538)
);

AND4x1_ASAP7_75t_L g1539 ( 
.A(n_1511),
.B(n_163),
.C(n_164),
.D(n_165),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1514),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1513),
.A2(n_409),
.B1(n_402),
.B2(n_172),
.Y(n_1541)
);

AOI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1493),
.A2(n_409),
.B1(n_402),
.B2(n_174),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1500),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1521),
.Y(n_1545)
);

AND4x1_ASAP7_75t_L g1546 ( 
.A(n_1491),
.B(n_166),
.C(n_169),
.D(n_176),
.Y(n_1546)
);

INVxp33_ASAP7_75t_L g1547 ( 
.A(n_1525),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1529),
.A2(n_1502),
.B1(n_1506),
.B2(n_1520),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1533),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1536),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1540),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1535),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1535),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1526),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1526),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1528),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1540),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1528),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1538),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1538),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1531),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1532),
.Y(n_1562)
);

INVxp33_ASAP7_75t_SL g1563 ( 
.A(n_1544),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1527),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1534),
.Y(n_1565)
);

OA22x2_ASAP7_75t_L g1566 ( 
.A1(n_1544),
.A2(n_1519),
.B1(n_1517),
.B2(n_1509),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1524),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1545),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1557),
.Y(n_1569)
);

AO22x1_ASAP7_75t_L g1570 ( 
.A1(n_1551),
.A2(n_1545),
.B1(n_1543),
.B2(n_1537),
.Y(n_1570)
);

OAI22x1_ASAP7_75t_L g1571 ( 
.A1(n_1551),
.A2(n_1546),
.B1(n_1559),
.B2(n_1560),
.Y(n_1571)
);

OAI22x1_ASAP7_75t_L g1572 ( 
.A1(n_1557),
.A2(n_1539),
.B1(n_1530),
.B2(n_1542),
.Y(n_1572)
);

AOI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1550),
.A2(n_1537),
.B1(n_1541),
.B2(n_1494),
.Y(n_1573)
);

AOI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1563),
.A2(n_1515),
.B1(n_1509),
.B2(n_1510),
.Y(n_1574)
);

AOI22xp5_ASAP7_75t_L g1575 ( 
.A1(n_1548),
.A2(n_402),
.B1(n_183),
.B2(n_184),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1552),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1565),
.A2(n_402),
.B1(n_185),
.B2(n_187),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1547),
.A2(n_179),
.B1(n_188),
.B2(n_199),
.Y(n_1578)
);

OAI22x1_ASAP7_75t_L g1579 ( 
.A1(n_1549),
.A2(n_200),
.B1(n_203),
.B2(n_209),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1569),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1571),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1576),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1570),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1572),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1584),
.A2(n_1553),
.B1(n_1549),
.B2(n_1568),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1583),
.A2(n_1575),
.B1(n_1547),
.B2(n_1573),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1581),
.A2(n_1556),
.B1(n_1566),
.B2(n_1554),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1581),
.A2(n_1566),
.B1(n_1558),
.B2(n_1555),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1588),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1587),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1585),
.Y(n_1591)
);

AOI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1590),
.A2(n_1586),
.B1(n_1580),
.B2(n_1567),
.Y(n_1592)
);

AOI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1591),
.A2(n_1558),
.B1(n_1564),
.B2(n_1582),
.Y(n_1593)
);

OAI22x1_ASAP7_75t_L g1594 ( 
.A1(n_1589),
.A2(n_1562),
.B1(n_1561),
.B2(n_1574),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1593),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1592),
.Y(n_1596)
);

AOI221xp5_ASAP7_75t_L g1597 ( 
.A1(n_1596),
.A2(n_1589),
.B1(n_1594),
.B2(n_1579),
.C(n_1578),
.Y(n_1597)
);

AOI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1597),
.A2(n_1595),
.B(n_1589),
.C(n_1577),
.Y(n_1598)
);


endmodule