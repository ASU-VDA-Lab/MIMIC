module fake_jpeg_1552_n_515 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_17),
.B(n_14),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_53),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_55),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_58),
.Y(n_120)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_64),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_17),
.B(n_13),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_66),
.Y(n_159)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_68),
.B(n_73),
.Y(n_151)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx11_ASAP7_75t_L g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_74),
.Y(n_164)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_75),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_79),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_80),
.B(n_84),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g144 ( 
.A(n_81),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_83),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx11_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_16),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_92),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_93),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_44),
.B(n_13),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_94),
.B(n_102),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_2),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_100),
.Y(n_155)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_25),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

BUFx16f_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx4_ASAP7_75t_SL g169 ( 
.A(n_112),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_118),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_103),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_67),
.B(n_45),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_125),
.B(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_89),
.A2(n_47),
.B1(n_48),
.B2(n_35),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_134),
.A2(n_41),
.B1(n_46),
.B2(n_38),
.Y(n_174)
);

CKINVDCx12_ASAP7_75t_R g136 ( 
.A(n_58),
.Y(n_136)
);

INVx4_ASAP7_75t_SL g183 ( 
.A(n_136),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_90),
.A2(n_47),
.B(n_39),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_137),
.B(n_19),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_100),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_78),
.B(n_41),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_34),
.B1(n_25),
.B2(n_32),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_145),
.A2(n_86),
.B1(n_34),
.B2(n_62),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_77),
.B(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_147),
.B(n_148),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_21),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_92),
.C(n_98),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_149),
.B(n_121),
.C(n_97),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_125),
.B1(n_137),
.B2(n_129),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_167),
.A2(n_168),
.B1(n_193),
.B2(n_208),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_152),
.B1(n_130),
.B2(n_159),
.Y(n_168)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_171),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_174),
.A2(n_175),
.B1(n_202),
.B2(n_215),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_112),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_180),
.Y(n_216)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_177),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_151),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_120),
.Y(n_182)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_185),
.Y(n_219)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_191),
.B(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_38),
.B1(n_46),
.B2(n_35),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_151),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_110),
.B(n_31),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_106),
.Y(n_197)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_123),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_201),
.Y(n_230)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_157),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_128),
.A2(n_54),
.B1(n_60),
.B2(n_82),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_131),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_204),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_110),
.B(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_146),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_111),
.B(n_31),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_209),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_207),
.B(n_20),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_116),
.A2(n_70),
.B1(n_81),
.B2(n_79),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_140),
.B(n_30),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_126),
.B(n_30),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_210),
.Y(n_236)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_132),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_211),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_108),
.A2(n_56),
.B1(n_76),
.B2(n_74),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_145),
.B1(n_165),
.B2(n_153),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_161),
.B(n_122),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_162),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_229),
.A2(n_249),
.B1(n_252),
.B2(n_182),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_172),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_167),
.A2(n_28),
.B(n_32),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_179),
.B(n_20),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_168),
.B(n_39),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_28),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_174),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_154),
.B1(n_34),
.B2(n_142),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_207),
.A2(n_122),
.B1(n_109),
.B2(n_107),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_221),
.B(n_170),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_266),
.Y(n_288)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_255),
.Y(n_286)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_257),
.Y(n_307)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_258),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_217),
.B1(n_223),
.B2(n_229),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_260),
.A2(n_274),
.B1(n_280),
.B2(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_198),
.C(n_178),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_261),
.B(n_265),
.C(n_183),
.Y(n_314)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_264),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_187),
.C(n_169),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_203),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_267),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_271),
.Y(n_285)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_190),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_236),
.B(n_169),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_242),
.A2(n_165),
.B1(n_115),
.B2(n_133),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_230),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_275),
.B(n_276),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_211),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_277),
.B(n_282),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_251),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_278),
.Y(n_309)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_231),
.A2(n_177),
.A3(n_186),
.B1(n_189),
.B2(n_173),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_218),
.B(n_246),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_217),
.A2(n_124),
.B1(n_133),
.B2(n_135),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_235),
.A2(n_202),
.B1(n_241),
.B2(n_226),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_281),
.A2(n_244),
.B1(n_225),
.B2(n_237),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_183),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_218),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_244),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_239),
.A2(n_124),
.B1(n_135),
.B2(n_164),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_290),
.A2(n_315),
.B1(n_274),
.B2(n_257),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_301),
.C(n_219),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_295),
.A2(n_300),
.B(n_306),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_225),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_303),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_259),
.A2(n_246),
.B(n_250),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_219),
.Y(n_301)
);

OA22x2_ASAP7_75t_L g303 ( 
.A1(n_281),
.A2(n_247),
.B1(n_239),
.B2(n_227),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_254),
.B(n_247),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_304),
.B(n_266),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_260),
.A2(n_250),
.B(n_228),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_228),
.B(n_222),
.Y(n_308)
);

AOI21xp33_ASAP7_75t_SL g335 ( 
.A1(n_308),
.A2(n_279),
.B(n_264),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_273),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_275),
.Y(n_317)
);

XNOR2x1_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_224),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_314),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_269),
.A2(n_188),
.B1(n_200),
.B2(n_238),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_317),
.B(n_328),
.Y(n_368)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_311),
.Y(n_319)
);

INVxp33_ASAP7_75t_L g372 ( 
.A(n_319),
.Y(n_372)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_320),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_310),
.Y(n_323)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_254),
.Y(n_325)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_325),
.Y(n_353)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_268),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_288),
.B(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_329),
.B(n_339),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_340),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_305),
.A2(n_280),
.B1(n_283),
.B2(n_271),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_332),
.A2(n_346),
.B1(n_295),
.B2(n_290),
.Y(n_352)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_292),
.Y(n_333)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_258),
.Y(n_334)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_334),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_335),
.A2(n_285),
.B(n_303),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_277),
.B1(n_284),
.B2(n_263),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_343),
.B1(n_309),
.B2(n_297),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_292),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_341),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_288),
.B(n_256),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_307),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_294),
.B(n_309),
.Y(n_342)
);

NOR3xp33_ASAP7_75t_SL g371 ( 
.A(n_342),
.B(n_303),
.C(n_286),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_314),
.C(n_293),
.Y(n_361)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_307),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_345),
.B(n_315),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_306),
.A2(n_238),
.B1(n_270),
.B2(n_255),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_350),
.A2(n_262),
.B1(n_248),
.B2(n_197),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_352),
.A2(n_356),
.B1(n_358),
.B2(n_339),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_316),
.A2(n_291),
.B1(n_289),
.B2(n_301),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_326),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_357),
.B(n_362),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_289),
.B1(n_301),
.B2(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_359),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_222),
.C(n_319),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_293),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_318),
.A2(n_335),
.B(n_328),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_366),
.B(n_369),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_314),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_371),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_318),
.A2(n_308),
.B(n_296),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_367),
.A2(n_375),
.B(n_319),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_296),
.B(n_285),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_334),
.A2(n_321),
.B(n_320),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_344),
.B(n_303),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_361),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_321),
.A2(n_303),
.B1(n_286),
.B2(n_287),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_332),
.B1(n_336),
.B2(n_343),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_379),
.A2(n_385),
.B1(n_387),
.B2(n_389),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_380),
.B(n_383),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_381),
.B(n_392),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_347),
.A2(n_346),
.B1(n_325),
.B2(n_330),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_382),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_330),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_384),
.B(n_396),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_352),
.A2(n_345),
.B1(n_340),
.B2(n_337),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_386),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_374),
.A2(n_358),
.B1(n_363),
.B2(n_353),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_377),
.A2(n_333),
.B1(n_323),
.B2(n_327),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_390),
.Y(n_411)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_355),
.Y(n_391)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_391),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_302),
.Y(n_393)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_393),
.Y(n_421)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_355),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_394),
.A2(n_395),
.B1(n_400),
.B2(n_403),
.Y(n_415)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_375),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_376),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_364),
.C(n_360),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_399),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_347),
.B(n_181),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_374),
.A2(n_215),
.B1(n_153),
.B2(n_164),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_354),
.B(n_224),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_404),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_353),
.A2(n_184),
.B1(n_156),
.B2(n_71),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_368),
.B(n_185),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_407),
.B(n_408),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_366),
.C(n_372),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_428),
.C(n_400),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_364),
.C(n_367),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_416),
.B(n_418),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_384),
.B(n_360),
.C(n_373),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_368),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_422),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_382),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_348),
.C(n_373),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_423),
.B(n_348),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_387),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_424),
.B(n_156),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_402),
.B(n_359),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_426),
.B(n_412),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_401),
.B(n_399),
.C(n_404),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_430),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_425),
.Y(n_431)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_405),
.B1(n_378),
.B2(n_379),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_432),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_389),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

XOR2x2_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_371),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_434),
.B(n_435),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_411),
.Y(n_436)
);

INVx11_ASAP7_75t_L g461 ( 
.A(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_440),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_439),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_426),
.A2(n_87),
.B(n_55),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_418),
.B(n_199),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_441),
.B(n_447),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_419),
.A2(n_199),
.B(n_109),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_444),
.B(n_448),
.C(n_412),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_413),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_446),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_409),
.A2(n_72),
.B1(n_163),
.B2(n_107),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_415),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_445),
.B(n_406),
.C(n_427),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_452),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_406),
.C(n_417),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_448),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_428),
.C(n_417),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_460),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_163),
.C(n_127),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_438),
.B(n_163),
.C(n_127),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_465),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_117),
.C(n_93),
.Y(n_465)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_453),
.Y(n_467)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_467),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_452),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_468),
.B(n_472),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_431),
.C(n_433),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_469),
.B(n_473),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_461),
.A2(n_429),
.B1(n_434),
.B2(n_436),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_471),
.A2(n_476),
.B1(n_465),
.B2(n_3),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_463),
.C(n_451),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_454),
.B(n_440),
.Y(n_474)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_446),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_457),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_478),
.B(n_479),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_459),
.B(n_117),
.Y(n_479)
);

MAJx2_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_93),
.C(n_3),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_480),
.B(n_481),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_51),
.C(n_22),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_466),
.C(n_464),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_487),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_475),
.Y(n_487)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_488),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_22),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_489),
.B(n_491),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_2),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_490),
.B(n_3),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_477),
.B(n_51),
.C(n_4),
.Y(n_491)
);

NAND3xp33_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_480),
.C(n_481),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_SL g502 ( 
.A(n_494),
.B(n_497),
.C(n_499),
.Y(n_502)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_493),
.A2(n_5),
.B(n_6),
.Y(n_497)
);

NOR3xp33_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_6),
.C(n_7),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_498),
.A2(n_483),
.B(n_489),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_485),
.A2(n_7),
.B(n_8),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_504),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_500),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_506),
.A2(n_485),
.B1(n_482),
.B2(n_486),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_502),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_508),
.B(n_509),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_507),
.A2(n_505),
.B(n_491),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_8),
.B(n_9),
.Y(n_512)
);

NOR5xp2_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_8),
.C(n_9),
.D(n_10),
.E(n_11),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_510),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_514),
.B(n_11),
.Y(n_515)
);


endmodule