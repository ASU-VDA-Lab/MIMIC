module fake_jpeg_4823_n_72 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_72);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_72;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_5),
.B(n_9),
.Y(n_13)
);

CKINVDCx5p33_ASAP7_75t_R g14 ( 
.A(n_8),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx24_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_27),
.Y(n_32)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_1),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_14),
.B(n_1),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_17),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_28),
.A2(n_17),
.B1(n_20),
.B2(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_18),
.C(n_21),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_41),
.C(n_48),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_22),
.C(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_15),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_55),
.C(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_47),
.B(n_37),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_46),
.B1(n_40),
.B2(n_42),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_29),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_39),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_62),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_56),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_50),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_12),
.B(n_10),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_63),
.B(n_65),
.C(n_54),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.C(n_64),
.Y(n_70)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_61),
.A3(n_59),
.B1(n_58),
.B2(n_8),
.C1(n_4),
.C2(n_3),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_67),
.Y(n_69)
);

BUFx24_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_65),
.B1(n_70),
.B2(n_61),
.Y(n_72)
);


endmodule