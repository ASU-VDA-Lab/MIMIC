module real_jpeg_23784_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_11;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_3),
.A2(n_20),
.B1(n_21),
.B2(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_27),
.B1(n_41),
.B2(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_4),
.A2(n_20),
.B1(n_21),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_7),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_7),
.A2(n_18),
.B(n_28),
.C(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_7),
.B(n_16),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_7),
.A2(n_20),
.B1(n_21),
.B2(n_34),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_7),
.B(n_40),
.C(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_7),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_7),
.B(n_38),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_8),
.B(n_72),
.Y(n_93)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_8),
.Y(n_101)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_8),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_75),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_73),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_58),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_12),
.B(n_58),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_48),
.Y(n_12)
);

XNOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_35),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_29),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_24),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_17)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_18),
.A2(n_23),
.B1(n_25),
.B2(n_28),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_20),
.A2(n_21),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_20),
.A2(n_23),
.B(n_34),
.Y(n_56)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_21),
.B(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_43),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_41),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_44),
.B(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B(n_54),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_71),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_51),
.B(n_54),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.C(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_65),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_70),
.B(n_108),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_88),
.B(n_112),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_84),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_77),
.B(n_84),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_81),
.B1(n_82),
.B2(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_96),
.B(n_111),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_94),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_109),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_105),
.B(n_110),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);


endmodule