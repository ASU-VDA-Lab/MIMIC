module fake_jpeg_24301_n_110 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_110);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_110;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_30;
wire n_106;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_10),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_26),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_0),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_32),
.B(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

AND2x4_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_25),
.Y(n_62)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_46),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

AND2x6_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_18),
.B1(n_13),
.B2(n_12),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_23),
.B1(n_20),
.B2(n_14),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_59),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_60),
.Y(n_69)
);

OR2x2_ASAP7_75t_SL g72 ( 
.A(n_62),
.B(n_41),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_29),
.C(n_33),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_59),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_73),
.B(n_62),
.C(n_52),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_79),
.C(n_80),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_67),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_71),
.B(n_62),
.C(n_61),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_65),
.C(n_68),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_43),
.C(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_54),
.C(n_37),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_50),
.C(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_64),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_72),
.C(n_74),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_2),
.C(n_3),
.Y(n_96)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_89),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_92),
.B1(n_67),
.B2(n_42),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_42),
.B1(n_90),
.B2(n_48),
.Y(n_99)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_1),
.B(n_2),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_97),
.B(n_88),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_96),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_96),
.B(n_9),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_101),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_48),
.C(n_24),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_7),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_22),
.B1(n_17),
.B2(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_100),
.B1(n_99),
.B2(n_101),
.Y(n_105)
);

AOI321xp33_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_106),
.A3(n_104),
.B1(n_10),
.B2(n_17),
.C(n_5),
.Y(n_107)
);

AO22x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_105),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_2),
.C(n_4),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_22),
.Y(n_110)
);


endmodule