module fake_jpeg_1173_n_95 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_95);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_95;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_41),
.B(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_28),
.B(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_29),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_45),
.Y(n_52)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_29),
.Y(n_46)
);

AO21x1_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_37),
.B(n_30),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_53),
.Y(n_60)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_55),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_35),
.B(n_33),
.C(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.Y(n_62)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_31),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_52),
.A2(n_54),
.B1(n_42),
.B2(n_56),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_59),
.A2(n_65),
.B1(n_6),
.B2(n_7),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_40),
.B1(n_38),
.B2(n_49),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_57),
.B1(n_51),
.B2(n_4),
.Y(n_72)
);

OAI32xp33_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_26),
.A3(n_49),
.B1(n_43),
.B2(n_3),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_68),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_49),
.B1(n_1),
.B2(n_2),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_66),
.A2(n_67),
.B(n_6),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_12),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_71),
.B(n_73),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_72),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_59),
.B(n_61),
.C(n_65),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_7),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_79),
.B(n_82),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_74),
.B1(n_25),
.B2(n_72),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_70),
.B(n_13),
.C(n_22),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_70),
.A2(n_17),
.B(n_19),
.Y(n_84)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_85),
.B(n_83),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_87),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_80),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_81),
.B(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_86),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_10),
.Y(n_95)
);


endmodule