module fake_jpeg_1668_n_314 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_23),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_49),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_47),
.Y(n_113)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

CKINVDCx9p33_ASAP7_75t_R g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_2),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_3),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_56),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_54),
.B(n_62),
.Y(n_134)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_3),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_31),
.Y(n_64)
);

INVx5_ASAP7_75t_SL g121 ( 
.A(n_64),
.Y(n_121)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_24),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_33),
.B1(n_36),
.B2(n_44),
.Y(n_101)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

AND2x4_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_89),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_24),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_71),
.B(n_84),
.Y(n_118)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_72),
.Y(n_106)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_17),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_77),
.Y(n_107)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_35),
.B(n_12),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_SL g80 ( 
.A1(n_28),
.A2(n_12),
.B(n_7),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_29),
.C(n_40),
.Y(n_117)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_83),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_6),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_86),
.B(n_87),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_34),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_27),
.B(n_34),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_27),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_56),
.A2(n_34),
.B1(n_25),
.B2(n_32),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_94),
.A2(n_97),
.B1(n_131),
.B2(n_39),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_44),
.B1(n_43),
.B2(n_40),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_61),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_109),
.B(n_66),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_25),
.B1(n_36),
.B2(n_33),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_112),
.A2(n_120),
.B1(n_93),
.B2(n_99),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_123),
.Y(n_145)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_79),
.C(n_57),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_48),
.A2(n_25),
.B1(n_43),
.B2(n_30),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_77),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_53),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_124),
.B(n_135),
.Y(n_162)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_127),
.Y(n_160)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_58),
.A2(n_38),
.B1(n_37),
.B2(n_30),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_64),
.B(n_38),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_67),
.B(n_37),
.C(n_39),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_79),
.C(n_76),
.Y(n_149)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_128),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_153),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_146),
.A2(n_152),
.B(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_91),
.B(n_65),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_154),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_149),
.B(n_151),
.Y(n_201)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_98),
.Y(n_150)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_150),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_60),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_133),
.B(n_78),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_74),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_69),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_168),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_97),
.B(n_66),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_92),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_159),
.B(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_7),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_166),
.B(n_106),
.Y(n_208)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_102),
.B(n_7),
.Y(n_168)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

BUFx24_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVx2_ASAP7_75t_R g172 ( 
.A(n_110),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_176),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_134),
.B(n_8),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_178),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_135),
.A2(n_57),
.B1(n_85),
.B2(n_39),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_110),
.B(n_8),
.Y(n_176)
);

AOI32xp33_ASAP7_75t_L g178 ( 
.A1(n_132),
.A2(n_9),
.A3(n_12),
.B1(n_115),
.B2(n_103),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_112),
.B(n_120),
.C(n_121),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_179),
.A2(n_180),
.B(n_149),
.C(n_151),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_109),
.A2(n_121),
.B(n_113),
.C(n_129),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_95),
.B(n_104),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_95),
.B(n_108),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_183),
.Y(n_200)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_138),
.B(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_125),
.B(n_108),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_190),
.A2(n_204),
.B(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_177),
.A2(n_126),
.B1(n_130),
.B2(n_141),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_199),
.B1(n_204),
.B2(n_212),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_144),
.A2(n_130),
.B1(n_139),
.B2(n_104),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_193),
.A2(n_160),
.B1(n_150),
.B2(n_143),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_157),
.A2(n_139),
.B1(n_100),
.B2(n_127),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_106),
.B1(n_129),
.B2(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_193),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_160),
.B(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_153),
.A2(n_179),
.B1(n_166),
.B2(n_162),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_216),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_169),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_151),
.B(n_173),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_171),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_170),
.C(n_164),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_190),
.C(n_217),
.Y(n_233)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_188),
.B(n_201),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_220),
.B(n_221),
.C(n_222),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_188),
.B(n_173),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_224),
.A2(n_237),
.B(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_225),
.A2(n_198),
.B1(n_214),
.B2(n_203),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_171),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_226),
.B(n_228),
.C(n_198),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_240),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_165),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_231),
.B(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_205),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_241),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_210),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_202),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_197),
.B(n_200),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_209),
.B(n_208),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_210),
.A2(n_207),
.B(n_205),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_238),
.A2(n_192),
.B(n_199),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_189),
.Y(n_239)
);

NOR2x1_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_218),
.Y(n_241)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_211),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_206),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_253),
.C(n_233),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_260),
.C(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_252),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_217),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_220),
.B(n_207),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_229),
.B(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_203),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_226),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_228),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_262),
.B(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_268),
.C(n_273),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_232),
.B1(n_243),
.B2(n_238),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_265),
.A2(n_272),
.B1(n_271),
.B2(n_247),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_258),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

BUFx12_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_252),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_240),
.B1(n_237),
.B2(n_230),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_222),
.C(n_221),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_274),
.B1(n_283),
.B2(n_271),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_253),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_257),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_284),
.C(n_261),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_285),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_257),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_274),
.A2(n_249),
.B1(n_250),
.B2(n_256),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_275),
.B(n_258),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_272),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_287),
.B(n_248),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_291),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_276),
.A2(n_275),
.B1(n_265),
.B2(n_245),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_284),
.C(n_280),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_275),
.B1(n_279),
.B2(n_278),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_293),
.A2(n_277),
.B1(n_248),
.B2(n_279),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_294),
.A2(n_286),
.B(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_300),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_292),
.C(n_280),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_293),
.C(n_288),
.Y(n_303)
);

OAI221xp5_ASAP7_75t_L g307 ( 
.A1(n_301),
.A2(n_290),
.B1(n_288),
.B2(n_294),
.C(n_298),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_307),
.B(n_308),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_296),
.B(n_279),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_304),
.C(n_291),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_304),
.C(n_282),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_311),
.B(n_312),
.C(n_227),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_242),
.A3(n_227),
.B1(n_259),
.B2(n_219),
.C1(n_225),
.C2(n_211),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_211),
.Y(n_314)
);


endmodule