module fake_jpeg_13427_n_177 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_48),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_16),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_0),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_58),
.B(n_2),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_3),
.Y(n_90)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_81),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_69),
.B(n_2),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_57),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_76),
.B1(n_70),
.B2(n_52),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_87),
.A2(n_67),
.B1(n_68),
.B2(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_88),
.B(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_66),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_86),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_96),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_59),
.B1(n_74),
.B2(n_71),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_54),
.B1(n_62),
.B2(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_53),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_25),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_52),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_108),
.B(n_7),
.Y(n_137)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_98),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_114),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_94),
.B(n_66),
.Y(n_107)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_75),
.C(n_73),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_60),
.B1(n_61),
.B2(n_75),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_30),
.B1(n_14),
.B2(n_17),
.Y(n_142)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_89),
.Y(n_114)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_93),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_116),
.B(n_105),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_118),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_100),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_10),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_4),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_114),
.B(n_27),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_11),
.C(n_18),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_139),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_135),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_4),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_5),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_109),
.B(n_6),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_140),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_137),
.A2(n_142),
.B(n_11),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_8),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_9),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_19),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_31),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_149),
.C(n_153),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_133),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_147),
.B(n_155),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_154),
.C(n_28),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_32),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_20),
.B1(n_22),
.B2(n_24),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_142),
.B(n_143),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_127),
.C(n_126),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_167)
);

NOR3xp33_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_137),
.C(n_131),
.Y(n_164)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_164),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_145),
.C(n_159),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_161),
.C(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_171),
.C(n_168),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_160),
.C(n_150),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_146),
.B(n_151),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_143),
.A3(n_158),
.B1(n_35),
.B2(n_39),
.C1(n_44),
.C2(n_29),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_33),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_138),
.B1(n_46),
.B2(n_49),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);


endmodule