module fake_ariane_2629_n_1114 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1114);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1114;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_952;
wire n_864;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_445;
wire n_379;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_210;
wire n_1090;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_218;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_658;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_741;
wire n_747;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_215;
wire n_664;
wire n_629;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_991;
wire n_834;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_895;
wire n_304;
wire n_862;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_967;
wire n_999;
wire n_998;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_976;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_211;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_50),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_150),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_68),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_184),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_58),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_87),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_197),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_205),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_107),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_102),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_104),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_196),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_8),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_154),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_52),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_123),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_202),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_137),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_144),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_207),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_161),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_192),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_76),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_96),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_22),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_187),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_8),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_151),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_38),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_209),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_118),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_30),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_157),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_112),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_67),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_44),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_163),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_94),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_60),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_19),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_85),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_32),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_99),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_182),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_179),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_66),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_131),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_93),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_210),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_221),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_220),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_235),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_241),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_225),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_233),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_231),
.Y(n_295)
);

INVxp33_ASAP7_75t_L g296 ( 
.A(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_254),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_235),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_263),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_275),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_222),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_266),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_267),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_271),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_259),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_234),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_278),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_211),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_243),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_256),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_213),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_214),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_261),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_215),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_212),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_276),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_222),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_274),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_324),
.B(n_237),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_325),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_289),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_249),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_325),
.Y(n_335)
);

OA21x2_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_219),
.B(n_217),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_274),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_289),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_289),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_319),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_307),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_280),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_281),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_289),
.Y(n_346)
);

CKINVDCx8_ASAP7_75t_R g347 ( 
.A(n_288),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_321),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_286),
.A2(n_279),
.B1(n_273),
.B2(n_270),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_300),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

NAND2xp33_ASAP7_75t_L g352 ( 
.A(n_283),
.B(n_212),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_240),
.B1(n_265),
.B2(n_262),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_320),
.A2(n_236),
.B1(n_258),
.B2(n_251),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_300),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_323),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_303),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_286),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_328),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_298),
.B(n_227),
.Y(n_364)
);

AND2x4_ASAP7_75t_L g365 ( 
.A(n_310),
.B(n_228),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_229),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_329),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_293),
.A2(n_230),
.B1(n_238),
.B2(n_244),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_284),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_287),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_294),
.B(n_245),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

AOI22x1_ASAP7_75t_SL g375 ( 
.A1(n_293),
.A2(n_246),
.B1(n_247),
.B2(n_248),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_299),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_301),
.B(n_212),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_212),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_305),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_306),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_308),
.Y(n_383)
);

AND2x4_ASAP7_75t_L g384 ( 
.A(n_309),
.B(n_0),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_353),
.B(n_316),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_335),
.Y(n_388)
);

AND2x2_ASAP7_75t_SL g389 ( 
.A(n_384),
.B(n_313),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_365),
.B(n_322),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_335),
.Y(n_391)
);

BUFx6f_ASAP7_75t_SL g392 ( 
.A(n_365),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_365),
.B(n_322),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_366),
.B(n_311),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_339),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g396 ( 
.A(n_343),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_366),
.B(n_312),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_332),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_341),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_341),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_343),
.B(n_315),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_376),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_355),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

OR2x2_ASAP7_75t_L g409 ( 
.A(n_337),
.B(n_285),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_370),
.B(n_282),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_359),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_369),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_332),
.Y(n_414)
);

NAND3xp33_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_320),
.C(n_290),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_360),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_362),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_369),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_367),
.Y(n_420)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_382),
.Y(n_421)
);

CKINVDCx6p67_ASAP7_75t_R g422 ( 
.A(n_342),
.Y(n_422)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_369),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_376),
.B(n_290),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_212),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_334),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_366),
.B(n_212),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_360),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_354),
.B(n_272),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g432 ( 
.A1(n_379),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_367),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_374),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_374),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_373),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_381),
.B(n_272),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_L g439 ( 
.A(n_377),
.B(n_272),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_374),
.B(n_272),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

CKINVDCx6p67_ASAP7_75t_R g442 ( 
.A(n_333),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_383),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_347),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_336),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_333),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_383),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_364),
.B(n_384),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_383),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_347),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_340),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_364),
.B(n_272),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_351),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_340),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_453),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_407),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

OR2x2_ASAP7_75t_SL g465 ( 
.A(n_415),
.B(n_375),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_330),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_368),
.Y(n_467)
);

BUFx6f_ASAP7_75t_SL g468 ( 
.A(n_389),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_407),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_450),
.B(n_330),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_410),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

INVxp33_ASAP7_75t_SL g474 ( 
.A(n_444),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_412),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_412),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_456),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_396),
.B(n_372),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_456),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_438),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_442),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_378),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_442),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_394),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_387),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_438),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_389),
.B(n_384),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_387),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_389),
.B(n_336),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_417),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_375),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_396),
.B(n_349),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_417),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_418),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_418),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_411),
.B(n_344),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_409),
.B(n_361),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_436),
.B(n_411),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_409),
.B(n_436),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_422),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_386),
.B(n_345),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_420),
.Y(n_506)
);

OR2x6_ASAP7_75t_L g507 ( 
.A(n_447),
.B(n_358),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_400),
.B(n_336),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_433),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_395),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_391),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_404),
.B(n_382),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_397),
.B(n_358),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_390),
.B(n_358),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_393),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_430),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_430),
.B(n_416),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_431),
.B(n_346),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_428),
.B(n_350),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_395),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_441),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_399),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_391),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_R g527 ( 
.A(n_426),
.B(n_340),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_392),
.B(n_443),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_R g529 ( 
.A(n_437),
.B(n_356),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_401),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_392),
.B(n_382),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_401),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_402),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_392),
.B(n_382),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_400),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_437),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_403),
.B(n_406),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_R g541 ( 
.A(n_443),
.B(n_357),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_466),
.B(n_470),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_466),
.B(n_441),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_470),
.B(n_451),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_499),
.B(n_502),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_468),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_505),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_500),
.B(n_358),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_479),
.B(n_502),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_499),
.A2(n_445),
.B1(n_451),
.B2(n_435),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_479),
.B(n_451),
.Y(n_552)
);

OAI22xp33_ASAP7_75t_L g553 ( 
.A1(n_488),
.A2(n_432),
.B1(n_455),
.B2(n_363),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_500),
.B(n_363),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_505),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_494),
.B(n_452),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_468),
.A2(n_445),
.B1(n_419),
.B2(n_448),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_483),
.B(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_460),
.B(n_413),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_462),
.Y(n_560)
);

OAI22xp33_ASAP7_75t_L g561 ( 
.A1(n_488),
.A2(n_494),
.B1(n_478),
.B2(n_480),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_SL g562 ( 
.A(n_482),
.B(n_423),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_509),
.B(n_413),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_507),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_505),
.B(n_454),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_467),
.B(n_419),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_474),
.B(n_519),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_485),
.B(n_424),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_498),
.B(n_363),
.Y(n_570)
);

O2A1O1Ixp5_ASAP7_75t_L g571 ( 
.A1(n_514),
.A2(n_459),
.B(n_398),
.C(n_408),
.Y(n_571)
);

O2A1O1Ixp5_ASAP7_75t_L g572 ( 
.A1(n_514),
.A2(n_459),
.B(n_398),
.C(n_408),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_486),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_519),
.B(n_434),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_489),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_507),
.B(n_363),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_504),
.B(n_434),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_484),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_538),
.B(n_434),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_507),
.B(n_424),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_490),
.A2(n_429),
.B1(n_435),
.B2(n_448),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_518),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_429),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_539),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_490),
.A2(n_352),
.B1(n_439),
.B2(n_351),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_516),
.B(n_398),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_539),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_515),
.B(n_398),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_503),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_481),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_529),
.A2(n_440),
.B1(n_338),
.B2(n_408),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_487),
.B(n_492),
.Y(n_593)
);

INVx4_ASAP7_75t_L g594 ( 
.A(n_523),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_495),
.B(n_408),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_496),
.B(n_414),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_528),
.B(n_414),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_497),
.B(n_414),
.Y(n_598)
);

AO22x1_ASAP7_75t_L g599 ( 
.A1(n_528),
.A2(n_458),
.B1(n_457),
.B2(n_446),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_517),
.A2(n_338),
.B1(n_446),
.B2(n_414),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_501),
.B(n_446),
.Y(n_601)
);

NAND2xp33_ASAP7_75t_SL g602 ( 
.A(n_506),
.B(n_446),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_457),
.Y(n_603)
);

INVxp33_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_L g605 ( 
.A(n_511),
.B(n_449),
.C(n_421),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_536),
.A2(n_338),
.B1(n_457),
.B2(n_458),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_537),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_540),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_521),
.B(n_458),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_338),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_546),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_547),
.B(n_563),
.Y(n_612)
);

BUFx4f_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_546),
.B(n_520),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_569),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_543),
.B(n_522),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_550),
.B(n_465),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g618 ( 
.A(n_594),
.B(n_531),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_579),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_590),
.Y(n_620)
);

BUFx4f_ASAP7_75t_SL g621 ( 
.A(n_547),
.Y(n_621)
);

AND3x1_ASAP7_75t_SL g622 ( 
.A(n_591),
.B(n_1),
.C(n_2),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_585),
.B(n_524),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_564),
.Y(n_624)
);

NOR2x1p5_ASAP7_75t_L g625 ( 
.A(n_594),
.B(n_607),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_566),
.B(n_525),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_566),
.B(n_530),
.Y(n_628)
);

CKINVDCx8_ASAP7_75t_R g629 ( 
.A(n_563),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_560),
.Y(n_630)
);

NOR3xp33_ASAP7_75t_SL g631 ( 
.A(n_553),
.B(n_527),
.C(n_531),
.Y(n_631)
);

NAND2xp33_ASAP7_75t_SL g632 ( 
.A(n_567),
.B(n_541),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_561),
.B(n_535),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g634 ( 
.A(n_564),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_556),
.B(n_542),
.Y(n_635)
);

CKINVDCx20_ASAP7_75t_R g636 ( 
.A(n_563),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_568),
.B(n_532),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_573),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_588),
.B(n_533),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_555),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_561),
.A2(n_535),
.B1(n_472),
.B2(n_471),
.Y(n_641)
);

INVx3_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_575),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_578),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_556),
.B(n_464),
.C(n_463),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_568),
.B(n_534),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_469),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_570),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_R g649 ( 
.A(n_548),
.B(n_510),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_555),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_607),
.A2(n_526),
.B1(n_513),
.B2(n_475),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_555),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_SL g653 ( 
.A(n_553),
.B(n_510),
.C(n_476),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_R g654 ( 
.A(n_548),
.B(n_473),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_609),
.A2(n_477),
.B1(n_449),
.B2(n_421),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

BUFx4f_ASAP7_75t_L g657 ( 
.A(n_576),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_593),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

NOR3xp33_ASAP7_75t_SL g660 ( 
.A(n_601),
.B(n_3),
.C(n_4),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_558),
.Y(n_661)
);

BUFx4f_ASAP7_75t_L g662 ( 
.A(n_549),
.Y(n_662)
);

INVx1_ASAP7_75t_SL g663 ( 
.A(n_554),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_584),
.B(n_421),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_552),
.B(n_423),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_610),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g668 ( 
.A(n_604),
.B(n_421),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_602),
.B(n_423),
.Y(n_669)
);

NAND3xp33_ASAP7_75t_SL g670 ( 
.A(n_600),
.B(n_4),
.C(n_5),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_595),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_545),
.Y(n_672)
);

AOI21xp33_ASAP7_75t_L g673 ( 
.A1(n_633),
.A2(n_551),
.B(n_584),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_635),
.A2(n_565),
.B(n_571),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_611),
.B(n_551),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_650),
.Y(n_676)
);

AO31x2_ASAP7_75t_L g677 ( 
.A1(n_647),
.A2(n_601),
.A3(n_589),
.B(n_587),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_589),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_616),
.B(n_557),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_616),
.B(n_557),
.Y(n_680)
);

BUFx6f_ASAP7_75t_SL g681 ( 
.A(n_612),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_634),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_627),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_619),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_658),
.B(n_587),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_617),
.A2(n_577),
.B(n_597),
.C(n_580),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_666),
.A2(n_572),
.B(n_582),
.Y(n_687)
);

OAI21x1_ASAP7_75t_L g688 ( 
.A1(n_672),
.A2(n_647),
.B(n_582),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_672),
.A2(n_574),
.B(n_596),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_614),
.A2(n_598),
.B1(n_606),
.B2(n_586),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_663),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_661),
.B(n_562),
.Y(n_692)
);

AND3x4_ASAP7_75t_L g693 ( 
.A(n_660),
.B(n_605),
.C(n_5),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_637),
.B(n_599),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_612),
.B(n_592),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_613),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_664),
.A2(n_423),
.B(n_272),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_638),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_625),
.B(n_423),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_645),
.A2(n_423),
.B(n_449),
.Y(n_700)
);

OAI21x1_ASAP7_75t_L g701 ( 
.A1(n_623),
.A2(n_449),
.B(n_33),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_624),
.B(n_6),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_624),
.B(n_6),
.Y(n_703)
);

OAI21x1_ASAP7_75t_L g704 ( 
.A1(n_623),
.A2(n_639),
.B(n_641),
.Y(n_704)
);

OAI21xp5_ASAP7_75t_L g705 ( 
.A1(n_653),
.A2(n_7),
.B(n_9),
.Y(n_705)
);

AO31x2_ASAP7_75t_L g706 ( 
.A1(n_639),
.A2(n_110),
.A3(n_204),
.B(n_201),
.Y(n_706)
);

INVxp67_ASAP7_75t_SL g707 ( 
.A(n_662),
.Y(n_707)
);

O2A1O1Ixp33_ASAP7_75t_L g708 ( 
.A1(n_670),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_646),
.B(n_10),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_630),
.Y(n_710)
);

CKINVDCx6p67_ASAP7_75t_R g711 ( 
.A(n_615),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_613),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_653),
.A2(n_11),
.B(n_12),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_11),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_671),
.A2(n_36),
.B(n_31),
.Y(n_715)
);

AOI21xp33_ASAP7_75t_L g716 ( 
.A1(n_626),
.A2(n_12),
.B(n_13),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_643),
.Y(n_717)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_665),
.A2(n_39),
.B(n_37),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_632),
.A2(n_41),
.B(n_40),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_644),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_648),
.B(n_13),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_620),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_642),
.A2(n_652),
.B(n_618),
.Y(n_723)
);

NOR2x1_ASAP7_75t_SL g724 ( 
.A(n_640),
.B(n_14),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_14),
.Y(n_725)
);

AO21x2_ASAP7_75t_L g726 ( 
.A1(n_649),
.A2(n_43),
.B(n_42),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_654),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_650),
.Y(n_728)
);

OAI21x1_ASAP7_75t_L g729 ( 
.A1(n_642),
.A2(n_46),
.B(n_45),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_631),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_730)
);

AO31x2_ASAP7_75t_L g731 ( 
.A1(n_659),
.A2(n_120),
.A3(n_200),
.B(n_199),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_683),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_674),
.A2(n_704),
.B(n_673),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_673),
.A2(n_670),
.B(n_669),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_722),
.B(n_621),
.Y(n_735)
);

INVx1_ASAP7_75t_SL g736 ( 
.A(n_691),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_682),
.B(n_652),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_705),
.A2(n_662),
.B1(n_636),
.B2(n_668),
.Y(n_738)
);

OA21x2_ASAP7_75t_L g739 ( 
.A1(n_697),
.A2(n_631),
.B(n_660),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_712),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_702),
.B(n_657),
.Y(n_741)
);

BUFx4_ASAP7_75t_SL g742 ( 
.A(n_696),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_710),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_701),
.A2(n_651),
.B(n_655),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_678),
.B(n_657),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_685),
.B(n_695),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_695),
.B(n_640),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_676),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_705),
.A2(n_640),
.B(n_667),
.Y(n_749)
);

OAI21x1_ASAP7_75t_L g750 ( 
.A1(n_687),
.A2(n_622),
.B(n_629),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_691),
.B(n_15),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_727),
.B(n_16),
.Y(n_752)
);

A2O1A1Ixp33_ASAP7_75t_L g753 ( 
.A1(n_713),
.A2(n_17),
.B(n_18),
.C(n_20),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_711),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_714),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_713),
.A2(n_18),
.B(n_20),
.Y(n_756)
);

OAI21x1_ASAP7_75t_L g757 ( 
.A1(n_688),
.A2(n_122),
.B(n_198),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_719),
.A2(n_21),
.B(n_22),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_689),
.A2(n_124),
.B(n_194),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_709),
.B(n_21),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_725),
.B(n_23),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_692),
.A2(n_23),
.B(n_24),
.Y(n_762)
);

AOI21xp33_ASAP7_75t_L g763 ( 
.A1(n_679),
.A2(n_24),
.B(n_25),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_675),
.B(n_25),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_708),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_765)
);

AO31x2_ASAP7_75t_L g766 ( 
.A1(n_679),
.A2(n_680),
.A3(n_690),
.B(n_686),
.Y(n_766)
);

AOI21x1_ASAP7_75t_L g767 ( 
.A1(n_680),
.A2(n_126),
.B(n_193),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_690),
.A2(n_27),
.B(n_28),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_693),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_769)
);

AO31x2_ASAP7_75t_L g770 ( 
.A1(n_720),
.A2(n_128),
.A3(n_49),
.B(n_51),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_703),
.B(n_29),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_698),
.Y(n_772)
);

AOI21x1_ASAP7_75t_L g773 ( 
.A1(n_694),
.A2(n_53),
.B(n_54),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_SL g774 ( 
.A1(n_730),
.A2(n_55),
.B(n_56),
.Y(n_774)
);

AOI221x1_ASAP7_75t_L g775 ( 
.A1(n_716),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.C(n_63),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_729),
.A2(n_64),
.B(n_65),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_684),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_717),
.A2(n_69),
.A3(n_70),
.B(n_71),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_676),
.B(n_73),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_700),
.A2(n_208),
.B(n_75),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_721),
.B(n_74),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_715),
.A2(n_77),
.B(n_79),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_718),
.B(n_80),
.Y(n_783)
);

AND2x4_ASAP7_75t_L g784 ( 
.A(n_707),
.B(n_81),
.Y(n_784)
);

OAI22x1_ASAP7_75t_L g785 ( 
.A1(n_699),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_699),
.B(n_86),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_716),
.A2(n_88),
.B(n_89),
.Y(n_787)
);

OAI21x1_ASAP7_75t_L g788 ( 
.A1(n_723),
.A2(n_90),
.B(n_91),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_676),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_677),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_728),
.B(n_92),
.Y(n_791)
);

BUFx4_ASAP7_75t_SL g792 ( 
.A(n_681),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_726),
.A2(n_190),
.B(n_97),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_728),
.B(n_189),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_732),
.Y(n_795)
);

INVx2_ASAP7_75t_R g796 ( 
.A(n_792),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_754),
.Y(n_797)
);

BUFx8_ASAP7_75t_SL g798 ( 
.A(n_777),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_736),
.B(n_677),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_734),
.A2(n_726),
.B(n_724),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_753),
.A2(n_681),
.B1(n_728),
.B2(n_677),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_SL g802 ( 
.A1(n_756),
.A2(n_731),
.B1(n_706),
.B2(n_100),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_743),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_706),
.B1(n_731),
.B2(n_101),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_736),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_766),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_746),
.A2(n_706),
.B1(n_98),
.B2(n_103),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_745),
.B(n_95),
.Y(n_809)
);

INVx6_ASAP7_75t_L g810 ( 
.A(n_748),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_742),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_764),
.B(n_105),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_766),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_740),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_733),
.A2(n_106),
.B(n_108),
.Y(n_815)
);

BUFx4f_ASAP7_75t_SL g816 ( 
.A(n_789),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_766),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_768),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_737),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_790),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_755),
.B(n_114),
.Y(n_821)
);

OAI22xp33_ASAP7_75t_L g822 ( 
.A1(n_769),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_822)
);

BUFx2_ASAP7_75t_L g823 ( 
.A(n_748),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_758),
.A2(n_782),
.B(n_793),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_751),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_770),
.Y(n_826)
);

OAI22xp33_ASAP7_75t_L g827 ( 
.A1(n_760),
.A2(n_119),
.B1(n_121),
.B2(n_125),
.Y(n_827)
);

BUFx4f_ASAP7_75t_SL g828 ( 
.A(n_741),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_786),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_735),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_770),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_761),
.A2(n_127),
.B1(n_129),
.B2(n_130),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_787),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_833)
);

BUFx4f_ASAP7_75t_SL g834 ( 
.A(n_747),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_770),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_786),
.B(n_136),
.Y(n_836)
);

BUFx8_ASAP7_75t_L g837 ( 
.A(n_771),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_752),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_765),
.A2(n_138),
.B1(n_140),
.B2(n_141),
.Y(n_839)
);

INVx6_ASAP7_75t_L g840 ( 
.A(n_784),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_778),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_778),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_784),
.Y(n_843)
);

OAI22xp33_ASAP7_75t_L g844 ( 
.A1(n_775),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_781),
.B(n_146),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_750),
.B(n_147),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_791),
.Y(n_847)
);

INVxp67_ASAP7_75t_SL g848 ( 
.A(n_739),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_843),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_795),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_839),
.A2(n_774),
.B1(n_762),
.B2(n_749),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_803),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_843),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_804),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_806),
.B(n_763),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_799),
.B(n_739),
.Y(n_856)
);

OAI21x1_ASAP7_75t_L g857 ( 
.A1(n_800),
.A2(n_757),
.B(n_767),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_826),
.A2(n_835),
.B(n_831),
.Y(n_858)
);

OAI21x1_ASAP7_75t_L g859 ( 
.A1(n_824),
.A2(n_744),
.B(n_759),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_820),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_807),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_819),
.B(n_785),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_814),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_840),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_830),
.B(n_811),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_829),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_813),
.Y(n_867)
);

INVx3_ASAP7_75t_L g868 ( 
.A(n_840),
.Y(n_868)
);

INVx4_ASAP7_75t_L g869 ( 
.A(n_823),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_841),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_842),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_828),
.Y(n_873)
);

BUFx3_ASAP7_75t_L g874 ( 
.A(n_816),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_848),
.B(n_773),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_810),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_825),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_838),
.Y(n_878)
);

OR2x2_ASAP7_75t_L g879 ( 
.A(n_801),
.B(n_794),
.Y(n_879)
);

OAI21x1_ASAP7_75t_L g880 ( 
.A1(n_805),
.A2(n_788),
.B(n_776),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_846),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_829),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_829),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_801),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_802),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_836),
.Y(n_886)
);

HB1xp67_ASAP7_75t_SL g887 ( 
.A(n_837),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_821),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_812),
.Y(n_889)
);

NAND4xp25_ASAP7_75t_SL g890 ( 
.A(n_832),
.B(n_780),
.C(n_783),
.D(n_779),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_810),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_809),
.Y(n_892)
);

BUFx3_ASAP7_75t_L g893 ( 
.A(n_874),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_857),
.Y(n_894)
);

AO21x2_ASAP7_75t_L g895 ( 
.A1(n_875),
.A2(n_844),
.B(n_815),
.Y(n_895)
);

OAI21x1_ASAP7_75t_L g896 ( 
.A1(n_857),
.A2(n_808),
.B(n_839),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_867),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_860),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_849),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_856),
.B(n_796),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_856),
.B(n_836),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_867),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_870),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_850),
.B(n_832),
.Y(n_904)
);

CKINVDCx11_ASAP7_75t_R g905 ( 
.A(n_874),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_870),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_873),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_860),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_859),
.A2(n_818),
.B(n_833),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_861),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_850),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_861),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_852),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_871),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_852),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_854),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_873),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_858),
.A2(n_818),
.B(n_783),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_854),
.B(n_845),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_871),
.Y(n_920)
);

HB1xp67_ASAP7_75t_L g921 ( 
.A(n_875),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_878),
.Y(n_922)
);

AOI21x1_ASAP7_75t_L g923 ( 
.A1(n_855),
.A2(n_847),
.B(n_837),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_877),
.B(n_827),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_899),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_895),
.A2(n_885),
.B1(n_884),
.B2(n_851),
.Y(n_926)
);

NOR3xp33_ASAP7_75t_L g927 ( 
.A(n_924),
.B(n_889),
.C(n_892),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_922),
.B(n_889),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_921),
.B(n_900),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_897),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_900),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_916),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_897),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_921),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_905),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_916),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_893),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_910),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_922),
.B(n_904),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_893),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_901),
.B(n_869),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_897),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_901),
.B(n_869),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_904),
.B(n_888),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_901),
.B(n_863),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_910),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_898),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_919),
.B(n_853),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_928),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_935),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_907),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_931),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_930),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_947),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_932),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_926),
.A2(n_885),
.B1(n_895),
.B2(n_904),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_936),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_935),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_931),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_930),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_939),
.B(n_898),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_937),
.B(n_893),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_944),
.B(n_919),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_927),
.B(n_908),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_951),
.B(n_945),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_962),
.B(n_945),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_962),
.B(n_941),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_956),
.B(n_908),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_963),
.B(n_929),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_956),
.B(n_938),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_950),
.B(n_941),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_952),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_949),
.B(n_929),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_959),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_964),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_953),
.Y(n_976)
);

INVx1_ASAP7_75t_SL g977 ( 
.A(n_958),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_966),
.B(n_950),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_SL g979 ( 
.A(n_977),
.B(n_950),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_975),
.Y(n_980)
);

INVxp67_ASAP7_75t_L g981 ( 
.A(n_972),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_973),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_968),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_SL g984 ( 
.A1(n_977),
.A2(n_954),
.B(n_964),
.C(n_957),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_965),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_978),
.B(n_935),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_985),
.B(n_950),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_983),
.B(n_974),
.Y(n_989)
);

AO221x2_ASAP7_75t_L g990 ( 
.A1(n_982),
.A2(n_935),
.B1(n_887),
.B2(n_958),
.C(n_968),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_980),
.B(n_958),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_981),
.Y(n_992)
);

OAI221xp5_ASAP7_75t_L g993 ( 
.A1(n_984),
.A2(n_970),
.B1(n_976),
.B2(n_923),
.C(n_892),
.Y(n_993)
);

NAND2xp33_ASAP7_75t_L g994 ( 
.A(n_988),
.B(n_958),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_987),
.B(n_967),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_992),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_990),
.B(n_935),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_989),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_993),
.B(n_969),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_991),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_955),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_992),
.A2(n_986),
.B(n_979),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_992),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_992),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_996),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_1003),
.Y(n_1006)
);

OAI22xp33_ASAP7_75t_SL g1007 ( 
.A1(n_999),
.A2(n_970),
.B1(n_979),
.B2(n_1000),
.Y(n_1007)
);

AOI221xp5_ASAP7_75t_L g1008 ( 
.A1(n_1002),
.A2(n_984),
.B1(n_924),
.B2(n_895),
.C(n_822),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_1004),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_1001),
.Y(n_1010)
);

AOI31xp33_ASAP7_75t_L g1011 ( 
.A1(n_997),
.A2(n_865),
.A3(n_971),
.B(n_940),
.Y(n_1011)
);

AOI31xp33_ASAP7_75t_L g1012 ( 
.A1(n_1000),
.A2(n_940),
.A3(n_798),
.B(n_797),
.Y(n_1012)
);

OA21x2_ASAP7_75t_L g1013 ( 
.A1(n_998),
.A2(n_961),
.B(n_960),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_1005),
.Y(n_1014)
);

AOI322xp5_ASAP7_75t_L g1015 ( 
.A1(n_1008),
.A2(n_1010),
.A3(n_1006),
.B1(n_1009),
.B2(n_1007),
.C1(n_994),
.C2(n_1013),
.Y(n_1015)
);

OAI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_1013),
.A2(n_994),
.B1(n_923),
.B2(n_995),
.C(n_917),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_1012),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1011),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1010),
.B(n_961),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1005),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_1005),
.Y(n_1021)
);

OAI221xp5_ASAP7_75t_L g1022 ( 
.A1(n_1008),
.A2(n_907),
.B1(n_917),
.B2(n_918),
.C(n_862),
.Y(n_1022)
);

OAI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_1022),
.A2(n_907),
.B1(n_917),
.B2(n_879),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_1015),
.A2(n_896),
.B(n_909),
.C(n_880),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_1018),
.A2(n_896),
.B(n_909),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_1017),
.B(n_797),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1016),
.A2(n_1021),
.B1(n_1020),
.B2(n_1014),
.Y(n_1027)
);

AOI221xp5_ASAP7_75t_L g1028 ( 
.A1(n_1019),
.A2(n_895),
.B1(n_894),
.B2(n_890),
.C(n_960),
.Y(n_1028)
);

AOI321xp33_ASAP7_75t_L g1029 ( 
.A1(n_1022),
.A2(n_884),
.A3(n_879),
.B1(n_881),
.B2(n_953),
.C(n_919),
.Y(n_1029)
);

OAI211xp5_ASAP7_75t_L g1030 ( 
.A1(n_1015),
.A2(n_934),
.B(n_925),
.C(n_899),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1026),
.Y(n_1031)
);

INVxp33_ASAP7_75t_SL g1032 ( 
.A(n_1027),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1030),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1024),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1025),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_1029),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1023),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_1028),
.Y(n_1038)
);

NOR4xp25_ASAP7_75t_L g1039 ( 
.A(n_1031),
.B(n_946),
.C(n_938),
.D(n_920),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1035),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1036),
.Y(n_1041)
);

NAND3xp33_ASAP7_75t_L g1042 ( 
.A(n_1033),
.B(n_894),
.C(n_918),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_1034),
.B(n_896),
.C(n_909),
.Y(n_1043)
);

NAND3xp33_ASAP7_75t_L g1044 ( 
.A(n_1037),
.B(n_894),
.C(n_918),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_1032),
.B(n_891),
.Y(n_1045)
);

NOR2x1_ASAP7_75t_L g1046 ( 
.A(n_1041),
.B(n_1036),
.Y(n_1046)
);

AOI211x1_ASAP7_75t_L g1047 ( 
.A1(n_1040),
.A2(n_1038),
.B(n_948),
.C(n_946),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_1045),
.B(n_1042),
.C(n_1043),
.Y(n_1048)
);

NOR4xp25_ASAP7_75t_L g1049 ( 
.A(n_1044),
.B(n_920),
.C(n_913),
.D(n_915),
.Y(n_1049)
);

AOI211xp5_ASAP7_75t_L g1050 ( 
.A1(n_1039),
.A2(n_894),
.B(n_911),
.C(n_913),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1041),
.B(n_894),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_1051),
.A2(n_894),
.B1(n_911),
.B2(n_915),
.C(n_933),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_1046),
.A2(n_918),
.B(n_891),
.C(n_876),
.Y(n_1053)
);

NAND4xp75_ASAP7_75t_L g1054 ( 
.A(n_1047),
.B(n_918),
.C(n_948),
.D(n_881),
.Y(n_1054)
);

AOI21xp33_ASAP7_75t_SL g1055 ( 
.A1(n_1048),
.A2(n_148),
.B(n_149),
.Y(n_1055)
);

OAI211xp5_ASAP7_75t_SL g1056 ( 
.A1(n_1050),
.A2(n_925),
.B(n_876),
.C(n_899),
.Y(n_1056)
);

NAND3xp33_ASAP7_75t_L g1057 ( 
.A(n_1049),
.B(n_894),
.C(n_886),
.Y(n_1057)
);

NAND4xp25_ASAP7_75t_SL g1058 ( 
.A(n_1046),
.B(n_925),
.C(n_943),
.D(n_869),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_1046),
.B(n_943),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_1046),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_L g1061 ( 
.A(n_1055),
.B(n_876),
.C(n_864),
.Y(n_1061)
);

OAI221xp5_ASAP7_75t_L g1062 ( 
.A1(n_1060),
.A2(n_886),
.B1(n_942),
.B2(n_933),
.C(n_914),
.Y(n_1062)
);

NAND4xp25_ASAP7_75t_SL g1063 ( 
.A(n_1059),
.B(n_943),
.C(n_942),
.D(n_882),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1060),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_1058),
.B(n_899),
.Y(n_1065)
);

NOR2x1_ASAP7_75t_L g1066 ( 
.A(n_1054),
.B(n_849),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1053),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_1057),
.B(n_914),
.Y(n_1068)
);

NAND3x1_ASAP7_75t_L g1069 ( 
.A(n_1052),
.B(n_853),
.C(n_864),
.Y(n_1069)
);

NAND3x1_ASAP7_75t_L g1070 ( 
.A(n_1064),
.B(n_1056),
.C(n_853),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1067),
.B(n_886),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_1065),
.B(n_849),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1068),
.Y(n_1073)
);

NOR3xp33_ASAP7_75t_L g1074 ( 
.A(n_1063),
.B(n_868),
.C(n_864),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_1061),
.B(n_886),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_1066),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1062),
.B(n_886),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1069),
.Y(n_1078)
);

NAND4xp75_ASAP7_75t_L g1079 ( 
.A(n_1064),
.B(n_914),
.C(n_912),
.D(n_910),
.Y(n_1079)
);

NAND4xp75_ASAP7_75t_L g1080 ( 
.A(n_1064),
.B(n_912),
.C(n_883),
.D(n_882),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1067),
.B(n_912),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1064),
.Y(n_1082)
);

NAND5xp2_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_152),
.C(n_153),
.D(n_155),
.E(n_156),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1076),
.Y(n_1084)
);

INVxp67_ASAP7_75t_SL g1085 ( 
.A(n_1073),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1081),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_SL g1087 ( 
.A1(n_1071),
.A2(n_834),
.B1(n_880),
.B2(n_868),
.Y(n_1087)
);

AOI221x1_ASAP7_75t_L g1088 ( 
.A1(n_1078),
.A2(n_868),
.B1(n_872),
.B2(n_866),
.C(n_883),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_1070),
.Y(n_1089)
);

AO22x2_ASAP7_75t_L g1090 ( 
.A1(n_1072),
.A2(n_1080),
.B1(n_1075),
.B2(n_1079),
.Y(n_1090)
);

AOI22x1_ASAP7_75t_L g1091 ( 
.A1(n_1077),
.A2(n_866),
.B1(n_159),
.B2(n_160),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1085),
.Y(n_1092)
);

BUFx8_ASAP7_75t_L g1093 ( 
.A(n_1084),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1091),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1089),
.A2(n_1074),
.B1(n_866),
.B2(n_859),
.Y(n_1095)
);

AOI31xp33_ASAP7_75t_L g1096 ( 
.A1(n_1086),
.A2(n_158),
.A3(n_162),
.B(n_165),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1090),
.Y(n_1097)
);

AO22x2_ASAP7_75t_L g1098 ( 
.A1(n_1092),
.A2(n_1088),
.B1(n_1083),
.B2(n_1087),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1097),
.A2(n_166),
.B(n_169),
.Y(n_1099)
);

XNOR2xp5_ASAP7_75t_L g1100 ( 
.A(n_1094),
.B(n_1093),
.Y(n_1100)
);

OAI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1099),
.A2(n_1095),
.B1(n_1096),
.B2(n_866),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_1101),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1102),
.A2(n_1100),
.B(n_1098),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1102),
.A2(n_170),
.B(n_171),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1103),
.A2(n_866),
.B1(n_903),
.B2(n_902),
.Y(n_1105)
);

OAI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1104),
.A2(n_903),
.B1(n_902),
.B2(n_906),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1103),
.A2(n_872),
.B1(n_903),
.B2(n_902),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1105),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1107),
.B(n_172),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_1106),
.B(n_173),
.Y(n_1110)
);

OR2x6_ASAP7_75t_L g1111 ( 
.A(n_1108),
.B(n_1110),
.Y(n_1111)
);

OR2x6_ASAP7_75t_L g1112 ( 
.A(n_1109),
.B(n_174),
.Y(n_1112)
);

AOI221xp5_ASAP7_75t_L g1113 ( 
.A1(n_1111),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.C(n_178),
.Y(n_1113)
);

AOI211xp5_ASAP7_75t_L g1114 ( 
.A1(n_1113),
.A2(n_1112),
.B(n_180),
.C(n_181),
.Y(n_1114)
);


endmodule