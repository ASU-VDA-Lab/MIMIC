module fake_jpeg_7011_n_124 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_124);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_25),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_27),
.A2(n_16),
.B1(n_21),
.B2(n_3),
.Y(n_50)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_21),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_22),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_40),
.Y(n_54)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_1),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_26),
.B1(n_23),
.B2(n_13),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_16),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_26),
.B1(n_23),
.B2(n_13),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_14),
.B1(n_20),
.B2(n_18),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_29),
.A2(n_14),
.B1(n_20),
.B2(n_18),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_57),
.B1(n_11),
.B2(n_4),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_3),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_39),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_4),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_35),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_31),
.C(n_36),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_72),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_66),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_31),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_68),
.Y(n_87)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_38),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_78),
.B(n_54),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_50),
.B(n_56),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_89),
.B(n_70),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_51),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_58),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_73),
.B1(n_64),
.B2(n_67),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_41),
.B(n_48),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_84),
.B(n_85),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_65),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_98),
.Y(n_102)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_71),
.B1(n_66),
.B2(n_64),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_99),
.B1(n_89),
.B2(n_86),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_96),
.A2(n_82),
.B(n_86),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

OAI32xp33_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_74),
.A3(n_57),
.B1(n_36),
.B2(n_61),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_100),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_106),
.B1(n_60),
.B2(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_108),
.A2(n_79),
.B(n_101),
.Y(n_110)
);

A2O1A1O1Ixp25_ASAP7_75t_L g109 ( 
.A1(n_106),
.A2(n_93),
.B(n_99),
.C(n_101),
.D(n_97),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_110),
.Y(n_117)
);

AO221x1_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_100),
.B1(n_91),
.B2(n_94),
.C(n_75),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_113),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_103),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_100),
.C(n_87),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_80),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_102),
.B1(n_60),
.B2(n_104),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_114),
.B(n_117),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_119),
.A2(n_116),
.B(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_120),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_121),
.B(n_11),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_123),
.B(n_68),
.Y(n_124)
);


endmodule