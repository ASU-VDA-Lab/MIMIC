module fake_jpeg_10399_n_57 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_57);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx11_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

INVx3_ASAP7_75t_SL g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_10),
.B1(n_9),
.B2(n_12),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_19),
.B1(n_12),
.B2(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_21),
.A2(n_20),
.B(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_13),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_8),
.B1(n_13),
.B2(n_17),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_33),
.B1(n_0),
.B2(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_6),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_24),
.A2(n_8),
.B1(n_1),
.B2(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_37),
.B(n_3),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_35),
.B1(n_38),
.B2(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_33),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_42),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_30),
.C(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_44),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_45),
.B(n_3),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.Y(n_51)
);

A2O1A1O1Ixp25_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_37),
.B(n_34),
.C(n_29),
.D(n_7),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_44),
.B1(n_43),
.B2(n_34),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_46),
.B1(n_47),
.B2(n_29),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_52),
.A2(n_53),
.B(n_51),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_17),
.C(n_4),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_54),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_51),
.C(n_4),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_17),
.Y(n_57)
);


endmodule