module fake_jpeg_21042_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_34),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_56),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_27),
.B(n_16),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_17),
.B(n_23),
.C(n_29),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_35),
.B(n_18),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_50),
.B(n_23),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_55),
.B1(n_20),
.B2(n_31),
.Y(n_81)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g92 ( 
.A(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_42),
.A2(n_25),
.B1(n_26),
.B2(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_60),
.B(n_19),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_18),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_26),
.B1(n_25),
.B2(n_32),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_62),
.A2(n_31),
.B1(n_20),
.B2(n_29),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_30),
.Y(n_84)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_89),
.B1(n_93),
.B2(n_57),
.Y(n_102)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx2_ASAP7_75t_SL g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_70),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_71),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_84),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_31),
.B1(n_20),
.B2(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_73),
.A2(n_81),
.B1(n_83),
.B2(n_97),
.Y(n_101)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_88),
.Y(n_100)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_46),
.B(n_56),
.C(n_59),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_95),
.C(n_30),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_82),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_60),
.B(n_33),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_86),
.Y(n_118)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_91),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_47),
.A2(n_28),
.B(n_22),
.C(n_17),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_17),
.B1(n_30),
.B2(n_21),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_30),
.C(n_21),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_23),
.B1(n_30),
.B2(n_17),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_102),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_103),
.A2(n_115),
.B1(n_92),
.B2(n_45),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_107),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g106 ( 
.A1(n_68),
.A2(n_57),
.B1(n_66),
.B2(n_48),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_74),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_75),
.A2(n_48),
.B(n_51),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_109),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_110),
.B(n_112),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_81),
.A2(n_66),
.B1(n_58),
.B2(n_63),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_116),
.B(n_0),
.Y(n_152)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_94),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_58),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_58),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_45),
.B(n_63),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_66),
.C(n_24),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_126),
.Y(n_164)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_109),
.A2(n_95),
.B1(n_79),
.B2(n_96),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_130),
.A2(n_133),
.B1(n_136),
.B2(n_150),
.Y(n_166)
);

INVxp33_ASAP7_75t_SL g131 ( 
.A(n_108),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_146),
.Y(n_159)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_80),
.B1(n_88),
.B2(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_106),
.C(n_115),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_45),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_106),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_105),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_140),
.B(n_148),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_77),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_142),
.B(n_103),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_106),
.B(n_69),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_92),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_143),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_117),
.Y(n_145)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_93),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_111),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_67),
.B1(n_92),
.B2(n_69),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_151),
.A2(n_153),
.B1(n_114),
.B2(n_119),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_154),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_103),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_0),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_121),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_121),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_124),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_157),
.B(n_162),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_161),
.B(n_167),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_155),
.A2(n_103),
.B1(n_110),
.B2(n_116),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_126),
.Y(n_162)
);

AND2x6_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_98),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_163),
.B(n_170),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_102),
.B1(n_101),
.B2(n_115),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_120),
.B(n_114),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_168),
.A2(n_1),
.B(n_2),
.Y(n_218)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

XNOR2x1_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_118),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_173),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_120),
.B(n_106),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_174),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_111),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_135),
.C(n_113),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_176),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_139),
.B(n_101),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_179),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_151),
.B1(n_147),
.B2(n_154),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_183),
.B1(n_133),
.B2(n_146),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_147),
.A2(n_106),
.B(n_45),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_R g193 ( 
.A(n_186),
.B(n_142),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_113),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_160),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_197),
.B(n_218),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_164),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_211),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_133),
.B(n_141),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_200),
.A2(n_203),
.B1(n_206),
.B2(n_217),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_183),
.B1(n_179),
.B2(n_163),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_132),
.B1(n_138),
.B2(n_140),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_213),
.Y(n_221)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_171),
.A2(n_127),
.B(n_156),
.C(n_152),
.D(n_137),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_205),
.B(n_160),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_172),
.B1(n_166),
.B2(n_187),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_165),
.B(n_119),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_210),
.B(n_185),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_212),
.B(n_195),
.C(n_197),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_166),
.A2(n_161),
.B1(n_158),
.B2(n_159),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_113),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_209),
.B(n_198),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_207),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_145),
.B1(n_90),
.B2(n_10),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_172),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_168),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_219),
.B(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_225),
.C(n_244),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_173),
.C(n_177),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_159),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_239),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_227),
.A2(n_242),
.B(n_2),
.Y(n_258)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_228),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_178),
.B1(n_184),
.B2(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_229),
.A2(n_207),
.B1(n_205),
.B2(n_202),
.Y(n_252)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_233),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_234),
.B(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_236),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_217),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_160),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_238),
.B(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_241),
.Y(n_261)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_212),
.C(n_206),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_203),
.B1(n_199),
.B2(n_209),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_204),
.C(n_219),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_253),
.C(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_238),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_225),
.B(n_218),
.C(n_192),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_15),
.C(n_13),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_230),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_231),
.B1(n_236),
.B2(n_242),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_258),
.A2(n_260),
.B(n_264),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_2),
.B(n_3),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_227),
.A2(n_10),
.B(n_11),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_226),
.C(n_221),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_253),
.C(n_250),
.Y(n_285)
);

OAI322xp33_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_239),
.A3(n_243),
.B1(n_233),
.B2(n_235),
.C1(n_223),
.C2(n_232),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_279),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_221),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_230),
.Y(n_272)
);

OAI321xp33_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_275),
.A3(n_231),
.B1(n_260),
.B2(n_276),
.C(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_229),
.Y(n_274)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_274),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_255),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_228),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_286),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_254),
.C(n_248),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_266),
.B(n_248),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_293),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_264),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_279),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_303),
.Y(n_307)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_261),
.B(n_265),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_272),
.Y(n_300)
);

NAND3xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_276),
.C(n_269),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_301),
.A2(n_305),
.B1(n_293),
.B2(n_11),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_294),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_283),
.A2(n_257),
.B(n_220),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_295),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_306),
.Y(n_317)
);

AO22x1_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_296),
.A2(n_285),
.B(n_292),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_309),
.A2(n_311),
.B(n_313),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_302),
.A2(n_281),
.B(n_289),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_4),
.Y(n_316)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_12),
.C2(n_298),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_300),
.B(n_298),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_316),
.B(n_307),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_318),
.B(n_7),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_319),
.B(n_320),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_314),
.C(n_317),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_7),
.B1(n_310),
.B2(n_322),
.Y(n_324)
);


endmodule