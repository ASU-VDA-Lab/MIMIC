module fake_ariane_1145_n_2251 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_236, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_54, n_25, n_2251);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_236;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2251;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2116;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_928;
wire n_253;
wire n_1153;
wire n_271;
wire n_465;
wire n_1103;
wire n_825;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_180),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_26),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_142),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_137),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_169),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_26),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_234),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_82),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_146),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_128),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_179),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_92),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_158),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_184),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_160),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_149),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_176),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_65),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_124),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_159),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_97),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_213),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_22),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_50),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_42),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_229),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_195),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_157),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_78),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_235),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_1),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_173),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_126),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_116),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_102),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_215),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_220),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_15),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g294 ( 
.A(n_2),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_141),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_204),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_162),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_27),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_53),
.Y(n_299)
);

BUFx8_ASAP7_75t_SL g300 ( 
.A(n_241),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_75),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_203),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_163),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_40),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_15),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_181),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_206),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_196),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_55),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_103),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_71),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_61),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_34),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_7),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_22),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_178),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_0),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_170),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_165),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_4),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_86),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_49),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_41),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_192),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_152),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_31),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_190),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_95),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_25),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_139),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_39),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_44),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_81),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_49),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_81),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_117),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_12),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_230),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_38),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_138),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_30),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_185),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_211),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_19),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_145),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_154),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_112),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_140),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_65),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_12),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_221),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_48),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_66),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_0),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_212),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_57),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_177),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_130),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_205),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_42),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_119),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_71),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_150),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_111),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_29),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_189),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_156),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_46),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_121),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_219),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_60),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_69),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_171),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_231),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_233),
.Y(n_376)
);

BUFx10_ASAP7_75t_L g377 ( 
.A(n_84),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_64),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_59),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_151),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_54),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_45),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_238),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_75),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_9),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_23),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_110),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_73),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_57),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_21),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_115),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_77),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_9),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_187),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_5),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_232),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_73),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_147),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_80),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_67),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_58),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_39),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_85),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_132),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_34),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_175),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_107),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_193),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_23),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_174),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_109),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_68),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_41),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_68),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_222),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_32),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_167),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_19),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_72),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_118),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_240),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_70),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_134),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_101),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_38),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_122),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_30),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_218),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_166),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_199),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_24),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_58),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_55),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_125),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_228),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_133),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_56),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_88),
.Y(n_438)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_191),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_31),
.Y(n_440)
);

BUFx10_ASAP7_75t_L g441 ( 
.A(n_99),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_197),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g443 ( 
.A(n_108),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_93),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_67),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_28),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_50),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_70),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_64),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_182),
.Y(n_450)
);

CKINVDCx14_ASAP7_75t_R g451 ( 
.A(n_96),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_237),
.Y(n_452)
);

BUFx2_ASAP7_75t_SL g453 ( 
.A(n_4),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_87),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_148),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_236),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_66),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_217),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_74),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_129),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_226),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_51),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_201),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_183),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_63),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_91),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_62),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_188),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_106),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_63),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_168),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_46),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_300),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_248),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_248),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_250),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_309),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_255),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_255),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_259),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_313),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_401),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_254),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_258),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_278),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_259),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_344),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_260),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_260),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_348),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_267),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_452),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_469),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_265),
.Y(n_496)
);

INVxp33_ASAP7_75t_SL g497 ( 
.A(n_412),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_267),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_249),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_244),
.Y(n_500)
);

INVxp33_ASAP7_75t_L g501 ( 
.A(n_418),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_400),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_244),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_251),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_270),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_270),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_257),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_244),
.Y(n_509)
);

CKINVDCx16_ASAP7_75t_R g510 ( 
.A(n_377),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_273),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_274),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_273),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_275),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_244),
.Y(n_515)
);

BUFx10_ASAP7_75t_L g516 ( 
.A(n_368),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_279),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_279),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_299),
.Y(n_519)
);

INVxp33_ASAP7_75t_SL g520 ( 
.A(n_453),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_304),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_286),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_312),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_314),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_307),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_307),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_317),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_443),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_329),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_443),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_331),
.Y(n_531)
);

INVxp67_ASAP7_75t_SL g532 ( 
.A(n_244),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_272),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_332),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_333),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_286),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_290),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_335),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_345),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_290),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_301),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_303),
.Y(n_542)
);

BUFx6f_ASAP7_75t_SL g543 ( 
.A(n_377),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_303),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_328),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_328),
.Y(n_546)
);

INVxp33_ASAP7_75t_SL g547 ( 
.A(n_453),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_339),
.Y(n_548)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_272),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_351),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_339),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_346),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_346),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_347),
.Y(n_554)
);

INVxp33_ASAP7_75t_SL g555 ( 
.A(n_353),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_347),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_354),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_355),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_358),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_358),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_320),
.Y(n_561)
);

CKINVDCx14_ASAP7_75t_R g562 ( 
.A(n_439),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_360),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_360),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_374),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_374),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_376),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_376),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_282),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_383),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_357),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_383),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_361),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_366),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_387),
.Y(n_575)
);

INVxp33_ASAP7_75t_SL g576 ( 
.A(n_369),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_280),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_387),
.Y(n_578)
);

INVxp33_ASAP7_75t_L g579 ( 
.A(n_294),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_391),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_391),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_280),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_291),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_291),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_377),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_394),
.Y(n_587)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_377),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_398),
.Y(n_589)
);

INVx1_ASAP7_75t_SL g590 ( 
.A(n_386),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_373),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_398),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_420),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_420),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_378),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_379),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_426),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_402),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_282),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_382),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_426),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_384),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_440),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_434),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_405),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_503),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_569),
.B(n_451),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_562),
.B(n_434),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_569),
.B(n_298),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_475),
.B(n_405),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_579),
.A2(n_445),
.B1(n_315),
.B2(n_416),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_509),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_500),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_500),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_510),
.B(n_438),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_599),
.B(n_298),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_515),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_515),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_496),
.A2(n_305),
.B1(n_322),
.B2(n_293),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_541),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_489),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_542),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_311),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_542),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_577),
.B(n_311),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_556),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_492),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_494),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_556),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_568),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_473),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_549),
.B(n_585),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_568),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_592),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_588),
.B(n_390),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_543),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_592),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_597),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_525),
.B(n_438),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_597),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_476),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_476),
.A2(n_456),
.B(n_455),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_480),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_526),
.B(n_390),
.Y(n_646)
);

OA21x2_ASAP7_75t_L g647 ( 
.A1(n_480),
.A2(n_456),
.B(n_455),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_481),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_481),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_528),
.B(n_295),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_482),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_482),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_488),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_488),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_495),
.B(n_407),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_490),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_530),
.B(n_458),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_490),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_555),
.B(n_458),
.Y(n_659)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_561),
.B(n_385),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_491),
.B(n_425),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_491),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_493),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_R g664 ( 
.A(n_499),
.B(n_242),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_493),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_477),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_498),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_498),
.Y(n_668)
);

NOR2x1_ASAP7_75t_L g669 ( 
.A(n_505),
.B(n_276),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_505),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_506),
.B(n_511),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_506),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_511),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_513),
.B(n_425),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_485),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_513),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_517),
.Y(n_677)
);

OAI21x1_ASAP7_75t_L g678 ( 
.A1(n_517),
.A2(n_463),
.B(n_461),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_518),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_518),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_522),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_478),
.Y(n_682)
);

CKINVDCx11_ASAP7_75t_R g683 ( 
.A(n_603),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_522),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_536),
.B(n_407),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_536),
.B(n_246),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_537),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_537),
.B(n_461),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_540),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_483),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_SL g691 ( 
.A(n_543),
.B(n_407),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_516),
.Y(n_692)
);

BUFx8_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_544),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_L g697 ( 
.A(n_504),
.B(n_508),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_545),
.B(n_546),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_545),
.B(n_463),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_546),
.B(n_246),
.Y(n_700)
);

AND2x6_ASAP7_75t_L g701 ( 
.A(n_548),
.B(n_284),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_548),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_486),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_643),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_608),
.B(n_576),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_659),
.A2(n_520),
.B1(n_547),
.B2(n_497),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_623),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_645),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_623),
.Y(n_709)
);

BUFx4f_ASAP7_75t_L g710 ( 
.A(n_643),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_623),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_664),
.B(n_512),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_693),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_623),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_633),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_620),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_685),
.B(n_533),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_648),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_649),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_R g720 ( 
.A(n_621),
.B(n_629),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_643),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_649),
.Y(n_722)
);

AND3x2_ASAP7_75t_L g723 ( 
.A(n_691),
.B(n_507),
.C(n_479),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_692),
.B(n_514),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_623),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_651),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_630),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_671),
.B(n_551),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_703),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_623),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_634),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_634),
.B(n_590),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_643),
.Y(n_733)
);

BUFx6f_ASAP7_75t_SL g734 ( 
.A(n_638),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_628),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_628),
.Y(n_736)
);

NOR2xp67_ASAP7_75t_L g737 ( 
.A(n_692),
.B(n_519),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_685),
.B(n_551),
.Y(n_738)
);

BUFx10_ASAP7_75t_L g739 ( 
.A(n_650),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_693),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_628),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_671),
.B(n_552),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_637),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_628),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_643),
.Y(n_745)
);

AOI22xp33_ASAP7_75t_L g746 ( 
.A1(n_657),
.A2(n_507),
.B1(n_502),
.B2(n_474),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_643),
.B(n_521),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_692),
.B(n_523),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_663),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_692),
.B(n_524),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_637),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_671),
.B(n_552),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_663),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_683),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_693),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_606),
.B(n_553),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_666),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_606),
.B(n_553),
.Y(n_758)
);

INVx5_ASAP7_75t_L g759 ( 
.A(n_663),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_628),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_615),
.B(n_527),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_628),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_691),
.A2(n_529),
.B1(n_534),
.B2(n_531),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_631),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_619),
.B(n_416),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_651),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_612),
.B(n_622),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_631),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_631),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_653),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_653),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_660),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_663),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_663),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_663),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_671),
.B(n_554),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_692),
.B(n_535),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_668),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_668),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_668),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_631),
.Y(n_781)
);

CKINVDCx6p67_ASAP7_75t_R g782 ( 
.A(n_692),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_612),
.B(n_554),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_626),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_668),
.B(n_656),
.Y(n_785)
);

OAI22xp33_ASAP7_75t_SL g786 ( 
.A1(n_611),
.A2(n_598),
.B1(n_484),
.B2(n_462),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_654),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_559),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_L g789 ( 
.A(n_655),
.B(n_539),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_607),
.B(n_550),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_698),
.B(n_559),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_658),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_658),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_698),
.B(n_560),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_662),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_607),
.B(n_557),
.Y(n_796)
);

NAND3xp33_ASAP7_75t_L g797 ( 
.A(n_697),
.B(n_573),
.C(n_558),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_631),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_675),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_698),
.B(n_661),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_605),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_693),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_638),
.B(n_591),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_631),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_638),
.B(n_595),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_662),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_605),
.B(n_582),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_672),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_638),
.B(n_596),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_635),
.Y(n_810)
);

INVx5_ASAP7_75t_L g811 ( 
.A(n_668),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_661),
.B(n_560),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_660),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_672),
.B(n_602),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_668),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_673),
.B(n_571),
.Y(n_816)
);

AND3x2_ASAP7_75t_L g817 ( 
.A(n_682),
.B(n_600),
.C(n_574),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_656),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_605),
.B(n_583),
.Y(n_819)
);

AND2x6_ASAP7_75t_L g820 ( 
.A(n_673),
.B(n_681),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_656),
.Y(n_821)
);

INVx3_ASAP7_75t_L g822 ( 
.A(n_635),
.Y(n_822)
);

AND2x6_ASAP7_75t_L g823 ( 
.A(n_681),
.B(n_466),
.Y(n_823)
);

CKINVDCx20_ASAP7_75t_R g824 ( 
.A(n_690),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_635),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_609),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_609),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_667),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_635),
.Y(n_829)
);

BUFx10_ASAP7_75t_L g830 ( 
.A(n_605),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_610),
.B(n_516),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_684),
.B(n_516),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_610),
.B(n_563),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_635),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_611),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_635),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_667),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_636),
.Y(n_838)
);

INVx8_ASAP7_75t_L g839 ( 
.A(n_686),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_667),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_686),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_667),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_SL g843 ( 
.A(n_684),
.B(n_563),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_610),
.A2(n_501),
.B1(n_565),
.B2(n_564),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_636),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_678),
.A2(n_565),
.B(n_564),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_636),
.Y(n_847)
);

AO21x2_ASAP7_75t_L g848 ( 
.A1(n_678),
.A2(n_699),
.B(n_688),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_687),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_644),
.A2(n_567),
.B(n_566),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_687),
.B(n_566),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_610),
.B(n_567),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_636),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_636),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_632),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_632),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_689),
.Y(n_857)
);

INVxp67_ASAP7_75t_SL g858 ( 
.A(n_636),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_689),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_632),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_644),
.Y(n_861)
);

NAND3xp33_ASAP7_75t_L g862 ( 
.A(n_627),
.B(n_604),
.C(n_572),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_652),
.Y(n_863)
);

NAND2xp33_ASAP7_75t_SL g864 ( 
.A(n_694),
.B(n_570),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_652),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_652),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_830),
.B(n_694),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_849),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_860),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_801),
.B(n_627),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_728),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_802),
.B(n_665),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_784),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_784),
.B(n_616),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_830),
.B(n_696),
.Y(n_875)
);

BUFx6f_ASAP7_75t_SL g876 ( 
.A(n_715),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_801),
.B(n_696),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_860),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_761),
.B(n_616),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_830),
.B(n_665),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_731),
.B(n_624),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_814),
.B(n_624),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_705),
.B(n_641),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_738),
.B(n_665),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_863),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_L g887 ( 
.A(n_820),
.B(n_670),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_728),
.B(n_670),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_843),
.A2(n_669),
.B1(n_676),
.B2(n_670),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_796),
.B(n_619),
.C(n_462),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_843),
.A2(n_669),
.B1(n_677),
.B2(n_676),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_743),
.B(n_676),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_857),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_743),
.B(n_677),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_863),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_732),
.B(n_646),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_742),
.B(n_677),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_742),
.B(n_679),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_752),
.B(n_679),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_818),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_752),
.B(n_679),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_818),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_776),
.B(n_680),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_821),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_723),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_864),
.A2(n_680),
.B1(n_702),
.B2(n_695),
.Y(n_906)
);

INVx3_ASAP7_75t_L g907 ( 
.A(n_842),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_864),
.A2(n_680),
.B1(n_702),
.B2(n_695),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_706),
.A2(n_695),
.B1(n_702),
.B2(n_389),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_720),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_765),
.A2(n_647),
.B1(n_644),
.B2(n_572),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_751),
.B(n_646),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_776),
.B(n_674),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_763),
.B(n_739),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_791),
.B(n_674),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_791),
.B(n_625),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_812),
.B(n_832),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_821),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_820),
.B(n_686),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_751),
.B(n_625),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_863),
.Y(n_921)
);

NAND2xp33_ASAP7_75t_L g922 ( 
.A(n_820),
.B(n_686),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_827),
.B(n_487),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_812),
.B(n_639),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_717),
.B(n_639),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_842),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_828),
.Y(n_927)
);

OR2x2_ASAP7_75t_L g928 ( 
.A(n_729),
.B(n_584),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_739),
.B(n_640),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_713),
.B(n_570),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_717),
.B(n_640),
.Y(n_931)
);

OAI221xp5_ASAP7_75t_L g932 ( 
.A1(n_844),
.A2(n_342),
.B1(n_340),
.B2(n_393),
.C(n_293),
.Y(n_932)
);

INVxp67_ASAP7_75t_L g933 ( 
.A(n_757),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_739),
.B(n_642),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_713),
.B(n_575),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_828),
.B(n_471),
.Y(n_936)
);

NOR2xp67_ASAP7_75t_L g937 ( 
.A(n_802),
.B(n_642),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_717),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_837),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_789),
.A2(n_700),
.B1(n_701),
.B2(n_686),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_837),
.B(n_471),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_716),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_820),
.A2(n_686),
.B1(n_701),
.B2(n_700),
.Y(n_943)
);

NAND2xp33_ASAP7_75t_L g944 ( 
.A(n_820),
.B(n_686),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_716),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_820),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_727),
.B(n_575),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_865),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_727),
.B(n_388),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_800),
.B(n_578),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_816),
.A2(n_800),
.B1(n_819),
.B2(n_807),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_840),
.B(n_578),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_794),
.B(n_580),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_826),
.B(n_580),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_840),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_790),
.B(n_767),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_L g957 ( 
.A(n_823),
.B(n_686),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_710),
.B(n_581),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_708),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_807),
.B(n_581),
.Y(n_960)
);

AND2x6_ASAP7_75t_L g961 ( 
.A(n_740),
.B(n_284),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_L g962 ( 
.A1(n_765),
.A2(n_647),
.B1(n_644),
.B2(n_587),
.Y(n_962)
);

OAI22xp33_ASAP7_75t_L g963 ( 
.A1(n_765),
.A2(n_587),
.B1(n_589),
.B2(n_586),
.Y(n_963)
);

OAI22xp33_ASAP7_75t_L g964 ( 
.A1(n_765),
.A2(n_589),
.B1(n_593),
.B2(n_586),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_865),
.Y(n_965)
);

INVx1_ASAP7_75t_SL g966 ( 
.A(n_757),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_799),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_807),
.B(n_593),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_866),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_819),
.B(n_594),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_866),
.Y(n_971)
);

INVxp67_ASAP7_75t_L g972 ( 
.A(n_799),
.Y(n_972)
);

INVx8_ASAP7_75t_L g973 ( 
.A(n_734),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_797),
.B(n_397),
.C(n_395),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_819),
.B(n_594),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_762),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_831),
.B(n_399),
.Y(n_977)
);

AND2x6_ASAP7_75t_SL g978 ( 
.A(n_754),
.B(n_305),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_746),
.A2(n_326),
.B1(n_323),
.B2(n_322),
.C(n_419),
.Y(n_979)
);

OR2x6_ASAP7_75t_L g980 ( 
.A(n_740),
.B(n_601),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_710),
.B(n_601),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_862),
.B(n_409),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_855),
.Y(n_983)
);

OAI22xp33_ASAP7_75t_L g984 ( 
.A1(n_835),
.A2(n_851),
.B1(n_604),
.B2(n_758),
.Y(n_984)
);

OAI21xp33_ASAP7_75t_L g985 ( 
.A1(n_718),
.A2(n_414),
.B(n_413),
.Y(n_985)
);

AND2x2_ASAP7_75t_SL g986 ( 
.A(n_785),
.B(n_647),
.Y(n_986)
);

INVx8_ASAP7_75t_L g987 ( 
.A(n_734),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_719),
.Y(n_988)
);

OAI221xp5_ASAP7_75t_L g989 ( 
.A1(n_833),
.A2(n_334),
.B1(n_393),
.B2(n_381),
.C(n_372),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_L g990 ( 
.A(n_823),
.B(n_700),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_722),
.B(n_647),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_747),
.A2(n_701),
.B1(n_700),
.B2(n_436),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_726),
.B(n_700),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_766),
.B(n_700),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_770),
.B(n_700),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_771),
.B(n_700),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_787),
.B(n_701),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_753),
.Y(n_998)
);

NAND3xp33_ASAP7_75t_L g999 ( 
.A(n_747),
.B(n_433),
.C(n_422),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_715),
.B(n_323),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_792),
.B(n_701),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_793),
.B(n_701),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_855),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_795),
.B(n_701),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_806),
.B(n_701),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_737),
.B(n_437),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_823),
.A2(n_372),
.B1(n_427),
.B2(n_431),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_808),
.B(n_446),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_859),
.B(n_618),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_715),
.B(n_326),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_856),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_835),
.B(n_334),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_756),
.B(n_618),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_783),
.B(n_618),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_788),
.B(n_618),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_813),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_852),
.B(n_454),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_754),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_710),
.B(n_436),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_712),
.B(n_449),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_823),
.B(n_337),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_762),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_823),
.B(n_337),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_753),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_SL g1025 ( 
.A(n_803),
.B(n_457),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_805),
.A2(n_459),
.B1(n_472),
.B2(n_465),
.Y(n_1026)
);

INVx2_ASAP7_75t_SL g1027 ( 
.A(n_755),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_823),
.B(n_338),
.Y(n_1028)
);

O2A1O1Ixp5_ASAP7_75t_L g1029 ( 
.A1(n_753),
.A2(n_245),
.B(n_404),
.C(n_350),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_724),
.B(n_467),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_900),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_884),
.B(n_755),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_923),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_884),
.B(n_782),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_983),
.Y(n_1035)
);

BUFx8_ASAP7_75t_L g1036 ( 
.A(n_876),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_902),
.Y(n_1037)
);

AND2x2_ASAP7_75t_SL g1038 ( 
.A(n_890),
.B(n_785),
.Y(n_1038)
);

AOI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_890),
.A2(n_824),
.B1(n_750),
.B2(n_777),
.Y(n_1039)
);

BUFx8_ASAP7_75t_L g1040 ( 
.A(n_876),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_871),
.A2(n_824),
.B1(n_748),
.B2(n_809),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_917),
.B(n_782),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_1012),
.A2(n_861),
.B1(n_786),
.B2(n_848),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_SL g1044 ( 
.A1(n_945),
.A2(n_772),
.B1(n_350),
.B2(n_363),
.Y(n_1044)
);

BUFx4f_ASAP7_75t_L g1045 ( 
.A(n_980),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_869),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_904),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_880),
.B(n_848),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_871),
.B(n_883),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_956),
.B(n_929),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_956),
.B(n_778),
.Y(n_1051)
);

INVx2_ASAP7_75t_SL g1052 ( 
.A(n_942),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_951),
.B(n_778),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_967),
.B(n_363),
.C(n_338),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_918),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_879),
.Y(n_1056)
);

INVx3_ASAP7_75t_L g1057 ( 
.A(n_946),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_947),
.B(n_419),
.C(n_381),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_1003),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_927),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1011),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_946),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_874),
.B(n_817),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_929),
.B(n_848),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_947),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_939),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_934),
.B(n_920),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_882),
.B(n_850),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_955),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_910),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_946),
.B(n_759),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_980),
.B(n_778),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_959),
.Y(n_1073)
);

BUFx4f_ASAP7_75t_L g1074 ( 
.A(n_980),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_963),
.B(n_759),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_938),
.B(n_861),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_973),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_930),
.B(n_861),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_886),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_934),
.B(n_822),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_895),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_973),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_907),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_973),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_921),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_984),
.A2(n_839),
.B1(n_408),
.B2(n_441),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_914),
.B(n_873),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_984),
.A2(n_839),
.B1(n_408),
.B2(n_441),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_896),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_988),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1009),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_979),
.A2(n_839),
.B1(n_408),
.B2(n_441),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_948),
.Y(n_1093)
);

A2O1A1Ixp33_ASAP7_75t_SL g1094 ( 
.A1(n_907),
.A2(n_845),
.B(n_853),
.C(n_822),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_966),
.B(n_431),
.C(n_427),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_965),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_926),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_926),
.B(n_841),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_920),
.B(n_822),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_870),
.B(n_845),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_924),
.Y(n_1101)
);

INVx5_ASAP7_75t_L g1102 ( 
.A(n_987),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_928),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_868),
.B(n_845),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_925),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_930),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1007),
.A2(n_932),
.B1(n_962),
.B2(n_911),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_892),
.B(n_853),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_931),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_969),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_935),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_963),
.B(n_759),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_SL g1113 ( 
.A1(n_933),
.A2(n_447),
.B1(n_448),
.B2(n_432),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_972),
.B(n_853),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_964),
.A2(n_721),
.B1(n_733),
.B2(n_704),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_964),
.A2(n_733),
.B1(n_745),
.B2(n_721),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_971),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_912),
.A2(n_749),
.B1(n_773),
.B2(n_745),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_976),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_1018),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_986),
.B(n_976),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_1000),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1007),
.A2(n_839),
.B1(n_408),
.B2(n_441),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_976),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_888),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_892),
.B(n_854),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1024),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_911),
.A2(n_407),
.B1(n_447),
.B2(n_432),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_998),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_SL g1130 ( 
.A(n_986),
.B(n_759),
.Y(n_1130)
);

OAI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_960),
.A2(n_448),
.B1(n_470),
.B2(n_779),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_912),
.A2(n_773),
.B1(n_815),
.B2(n_749),
.Y(n_1132)
);

NOR2x2_ASAP7_75t_L g1133 ( 
.A(n_949),
.B(n_336),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_894),
.B(n_854),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_L g1135 ( 
.A(n_877),
.B(n_854),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_976),
.B(n_759),
.Y(n_1136)
);

NOR3xp33_ASAP7_75t_SL g1137 ( 
.A(n_1025),
.B(n_470),
.C(n_247),
.Y(n_1137)
);

BUFx3_ASAP7_75t_L g1138 ( 
.A(n_987),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_894),
.B(n_774),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_1022),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_935),
.B(n_841),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_950),
.B(n_774),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_897),
.A2(n_780),
.B(n_775),
.C(n_779),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_1027),
.B(n_841),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_998),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_898),
.Y(n_1146)
);

NOR2x2_ASAP7_75t_L g1147 ( 
.A(n_978),
.B(n_336),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_899),
.Y(n_1148)
);

NOR2x1p5_ASAP7_75t_L g1149 ( 
.A(n_1010),
.B(n_846),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_954),
.B(n_775),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_901),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_SL g1152 ( 
.A(n_974),
.B(n_252),
.C(n_243),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1022),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1022),
.Y(n_1154)
);

AOI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1020),
.A2(n_780),
.B1(n_815),
.B2(n_858),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_991),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_1016),
.B(n_707),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_968),
.B(n_707),
.Y(n_1158)
);

NOR3xp33_ASAP7_75t_SL g1159 ( 
.A(n_1008),
.B(n_256),
.C(n_253),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_970),
.B(n_709),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_975),
.B(n_709),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_893),
.B(n_711),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_L g1163 ( 
.A1(n_993),
.A2(n_846),
.B(n_714),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_867),
.B(n_841),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_903),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_SL g1166 ( 
.A(n_962),
.B(n_811),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1020),
.A2(n_847),
.B1(n_838),
.B2(n_836),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_913),
.B(n_711),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_915),
.B(n_714),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_994),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_905),
.B(n_725),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_916),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1008),
.B(n_725),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_953),
.B(n_730),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_878),
.B(n_885),
.Y(n_1175)
);

OR2x6_ASAP7_75t_L g1176 ( 
.A(n_987),
.B(n_730),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_SL g1177 ( 
.A(n_867),
.B(n_811),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_961),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_952),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_961),
.Y(n_1180)
);

AOI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_875),
.A2(n_847),
.B1(n_735),
.B2(n_838),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_982),
.A2(n_741),
.B1(n_836),
.B2(n_834),
.Y(n_1182)
);

AOI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_875),
.A2(n_769),
.B1(n_834),
.B2(n_736),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_982),
.B(n_1030),
.Y(n_1184)
);

NAND2xp33_ASAP7_75t_L g1185 ( 
.A(n_974),
.B(n_762),
.Y(n_1185)
);

AO22x1_ASAP7_75t_L g1186 ( 
.A1(n_961),
.A2(n_841),
.B1(n_352),
.B2(n_415),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1030),
.B(n_735),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_909),
.B(n_736),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_961),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_887),
.B(n_734),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_952),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_977),
.B(n_741),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_961),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_906),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_1021),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1023),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_995),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_908),
.Y(n_1198)
);

AND3x1_ASAP7_75t_L g1199 ( 
.A(n_977),
.B(n_760),
.C(n_744),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_996),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_937),
.B(n_760),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_889),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_997),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_985),
.B(n_764),
.Y(n_1204)
);

INVx2_ASAP7_75t_SL g1205 ( 
.A(n_1028),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1017),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_891),
.A2(n_769),
.B(n_764),
.C(n_768),
.Y(n_1207)
);

NOR2xp67_ASAP7_75t_L g1208 ( 
.A(n_872),
.B(n_781),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1013),
.Y(n_1209)
);

AOI21xp33_ASAP7_75t_L g1210 ( 
.A1(n_1001),
.A2(n_1004),
.B(n_1002),
.Y(n_1210)
);

OR2x4_ASAP7_75t_L g1211 ( 
.A(n_1005),
.B(n_762),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_881),
.A2(n_798),
.B(n_781),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1050),
.B(n_1026),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1045),
.B(n_999),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1120),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_SL g1216 ( 
.A(n_1065),
.B(n_881),
.Y(n_1216)
);

O2A1O1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1067),
.A2(n_936),
.B(n_941),
.C(n_1006),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1103),
.B(n_936),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1034),
.A2(n_981),
.B(n_958),
.Y(n_1219)
);

AO32x1_ASAP7_75t_L g1220 ( 
.A1(n_1173),
.A2(n_810),
.A3(n_804),
.B1(n_798),
.B2(n_614),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1082),
.B(n_958),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1049),
.B(n_1014),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1163),
.A2(n_810),
.B(n_804),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_SL g1224 ( 
.A(n_1045),
.B(n_989),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1073),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1175),
.A2(n_1048),
.B(n_1064),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_L g1227 ( 
.A1(n_1184),
.A2(n_1019),
.B(n_941),
.C(n_981),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_R g1228 ( 
.A(n_1070),
.B(n_1082),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_1032),
.B(n_1087),
.Y(n_1229)
);

OR2x6_ASAP7_75t_SL g1230 ( 
.A(n_1036),
.B(n_261),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1036),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1087),
.B(n_1015),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1108),
.A2(n_922),
.B(n_919),
.Y(n_1233)
);

AOI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1166),
.A2(n_1019),
.B(n_614),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1172),
.B(n_940),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1074),
.B(n_943),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1040),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1126),
.A2(n_944),
.B(n_957),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1176),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1040),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_SL g1241 ( 
.A(n_1074),
.B(n_1077),
.Y(n_1241)
);

BUFx6f_ASAP7_75t_L g1242 ( 
.A(n_1084),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1138),
.B(n_811),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1044),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_1103),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1090),
.Y(n_1246)
);

CKINVDCx16_ASAP7_75t_R g1247 ( 
.A(n_1138),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1059),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1212),
.A2(n_1029),
.B(n_992),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1106),
.B(n_762),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1089),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1031),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1037),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1052),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_SL g1255 ( 
.A(n_1041),
.B(n_825),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1047),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1089),
.B(n_613),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_SL g1258 ( 
.A(n_1042),
.B(n_825),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1055),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1061),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1111),
.B(n_1078),
.Y(n_1261)
);

O2A1O1Ixp5_ASAP7_75t_L g1262 ( 
.A1(n_1177),
.A2(n_614),
.B(n_613),
.C(n_617),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1078),
.B(n_825),
.Y(n_1263)
);

NOR2x1_ASAP7_75t_L g1264 ( 
.A(n_1077),
.B(n_990),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1134),
.A2(n_811),
.B(n_825),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1060),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1101),
.B(n_829),
.Y(n_1267)
);

NOR3xp33_ASAP7_75t_SL g1268 ( 
.A(n_1095),
.B(n_263),
.C(n_262),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1106),
.B(n_829),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1099),
.A2(n_829),
.B(n_352),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1122),
.B(n_613),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1105),
.B(n_829),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1139),
.A2(n_411),
.B(n_349),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1176),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1051),
.A2(n_415),
.B(n_411),
.C(n_349),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_R g1276 ( 
.A(n_1084),
.B(n_264),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1033),
.B(n_617),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1084),
.B(n_617),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1053),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1051),
.A2(n_435),
.B(n_428),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1080),
.A2(n_435),
.B(n_428),
.Y(n_1281)
);

O2A1O1Ixp33_ASAP7_75t_L g1282 ( 
.A1(n_1125),
.A2(n_276),
.B(n_330),
.C(n_444),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1066),
.Y(n_1283)
);

AOI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1166),
.A2(n_444),
.B(n_330),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_R g1285 ( 
.A(n_1084),
.B(n_266),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1063),
.B(n_1),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1102),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1094),
.A2(n_1142),
.B(n_1210),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1094),
.A2(n_435),
.B(n_428),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1069),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1035),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1109),
.B(n_2),
.Y(n_1292)
);

OR2x6_ASAP7_75t_L g1293 ( 
.A(n_1141),
.B(n_428),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1058),
.B(n_268),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1168),
.A2(n_428),
.B(n_435),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1192),
.A2(n_468),
.B(n_464),
.C(n_460),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1146),
.B(n_3),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1169),
.A2(n_435),
.B(n_442),
.Y(n_1298)
);

O2A1O1Ixp5_ASAP7_75t_SL g1299 ( 
.A1(n_1121),
.A2(n_450),
.B(n_430),
.C(n_429),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1192),
.A2(n_424),
.B(n_423),
.C(n_421),
.Y(n_1300)
);

INVx8_ASAP7_75t_L g1301 ( 
.A(n_1102),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1072),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1157),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1046),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1148),
.A2(n_3),
.B(n_5),
.C(n_6),
.Y(n_1305)
);

NOR2xp33_ASAP7_75t_L g1306 ( 
.A(n_1039),
.B(n_269),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_1046),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1053),
.A2(n_417),
.B(n_410),
.C(n_406),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1107),
.A2(n_403),
.B1(n_396),
.B2(n_380),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1151),
.B(n_6),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1056),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1121),
.A2(n_375),
.B(n_371),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1056),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_1102),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1206),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1165),
.B(n_7),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1128),
.A2(n_370),
.B1(n_367),
.B2(n_365),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1079),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1143),
.A2(n_364),
.B(n_362),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1079),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1156),
.A2(n_105),
.B(n_227),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1209),
.B(n_8),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1202),
.B(n_8),
.Y(n_1323)
);

BUFx12f_ASAP7_75t_L g1324 ( 
.A(n_1102),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1072),
.B(n_10),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1150),
.B(n_10),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1054),
.Y(n_1327)
);

A2O1A1Ixp33_ASAP7_75t_L g1328 ( 
.A1(n_1086),
.A2(n_359),
.B(n_356),
.C(n_343),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1195),
.B(n_1092),
.Y(n_1329)
);

AO32x2_ASAP7_75t_L g1330 ( 
.A1(n_1196),
.A2(n_11),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_1330)
);

INVx4_ASAP7_75t_L g1331 ( 
.A(n_1176),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1128),
.A2(n_341),
.B1(n_327),
.B2(n_325),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1038),
.B(n_271),
.Y(n_1333)
);

INVxp67_ASAP7_75t_SL g1334 ( 
.A(n_1119),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1092),
.B(n_11),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1086),
.A2(n_324),
.B1(n_321),
.B2(n_319),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1038),
.A2(n_292),
.B1(n_316),
.B2(n_310),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1091),
.B(n_13),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1143),
.A2(n_288),
.B(n_308),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1068),
.B(n_14),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1123),
.A2(n_318),
.B1(n_306),
.B2(n_302),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_SL g1342 ( 
.A(n_1141),
.B(n_297),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1076),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1187),
.A2(n_289),
.B(n_287),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1057),
.B(n_296),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1081),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1081),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1149),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1152),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1349)
);

NOR2xp33_ASAP7_75t_SL g1350 ( 
.A(n_1189),
.B(n_277),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1083),
.B(n_281),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1194),
.B(n_17),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1057),
.B(n_18),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1085),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1123),
.A2(n_285),
.B1(n_283),
.B2(n_24),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1198),
.B(n_20),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1171),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1211),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1100),
.A2(n_20),
.B(n_21),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1131),
.B(n_25),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1174),
.A2(n_27),
.B(n_28),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1054),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1131),
.B(n_29),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_SL g1364 ( 
.A(n_1113),
.B(n_32),
.C(n_33),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1088),
.A2(n_1043),
.B1(n_1205),
.B2(n_1156),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1130),
.A2(n_33),
.B(n_35),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1043),
.B(n_35),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1254),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1279),
.B(n_1179),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1223),
.A2(n_1199),
.B(n_1130),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1213),
.A2(n_1279),
.B1(n_1229),
.B2(n_1088),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1288),
.A2(n_1207),
.B(n_1188),
.Y(n_1372)
);

NOR3xp33_ASAP7_75t_L g1373 ( 
.A(n_1349),
.B(n_1185),
.C(n_1114),
.Y(n_1373)
);

AOI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1288),
.A2(n_1177),
.B(n_1186),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1228),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1251),
.B(n_1137),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1232),
.B(n_1191),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_SL g1378 ( 
.A1(n_1219),
.A2(n_1132),
.B(n_1118),
.Y(n_1378)
);

BUFx10_ASAP7_75t_L g1379 ( 
.A(n_1237),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1251),
.B(n_1119),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1225),
.Y(n_1381)
);

NAND2x1_ASAP7_75t_L g1382 ( 
.A(n_1242),
.B(n_1124),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1222),
.B(n_1226),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1265),
.A2(n_1197),
.B(n_1200),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1324),
.Y(n_1385)
);

NOR2xp67_ASAP7_75t_L g1386 ( 
.A(n_1215),
.B(n_1062),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1226),
.A2(n_1136),
.B(n_1112),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1233),
.A2(n_1136),
.B(n_1112),
.Y(n_1388)
);

INVx4_ASAP7_75t_L g1389 ( 
.A(n_1301),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1245),
.B(n_1137),
.Y(n_1390)
);

OAI21xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1333),
.A2(n_1075),
.B(n_1135),
.Y(n_1391)
);

BUFx4f_ASAP7_75t_SL g1392 ( 
.A(n_1240),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1265),
.A2(n_1281),
.B(n_1295),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1281),
.A2(n_1170),
.B(n_1197),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1238),
.A2(n_1207),
.B(n_1071),
.Y(n_1395)
);

INVx4_ASAP7_75t_L g1396 ( 
.A(n_1301),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1360),
.A2(n_1159),
.B1(n_1115),
.B2(n_1116),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1303),
.B(n_1083),
.Y(n_1398)
);

NAND2x1_ASAP7_75t_L g1399 ( 
.A(n_1242),
.B(n_1124),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1306),
.A2(n_1159),
.B(n_1155),
.C(n_1204),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1218),
.B(n_1097),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1217),
.A2(n_1204),
.B(n_1135),
.C(n_1104),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1295),
.A2(n_1167),
.B(n_1208),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1217),
.A2(n_1104),
.B(n_1162),
.C(n_1062),
.Y(n_1404)
);

AO21x1_ASAP7_75t_L g1405 ( 
.A1(n_1275),
.A2(n_1162),
.B(n_1071),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1315),
.B(n_1357),
.Y(n_1406)
);

INVxp67_ASAP7_75t_L g1407 ( 
.A(n_1286),
.Y(n_1407)
);

AOI211x1_ASAP7_75t_L g1408 ( 
.A1(n_1363),
.A2(n_1158),
.B(n_1160),
.C(n_1161),
.Y(n_1408)
);

O2A1O1Ixp33_ASAP7_75t_SL g1409 ( 
.A1(n_1340),
.A2(n_1129),
.B(n_1145),
.C(n_1097),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1302),
.B(n_1093),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1349),
.A2(n_1145),
.B(n_1127),
.C(n_1110),
.Y(n_1411)
);

AOI211x1_ASAP7_75t_L g1412 ( 
.A1(n_1335),
.A2(n_1201),
.B(n_1133),
.C(n_43),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1234),
.A2(n_1170),
.B(n_1203),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1348),
.B(n_1153),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1280),
.A2(n_1119),
.B(n_1140),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_SL g1416 ( 
.A(n_1224),
.B(n_1140),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1289),
.A2(n_1182),
.B(n_1181),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1365),
.B(n_1154),
.Y(n_1418)
);

OAI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1227),
.A2(n_1183),
.B(n_1182),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1275),
.A2(n_1193),
.B(n_1178),
.C(n_1180),
.Y(n_1420)
);

A2O1A1Ixp33_ASAP7_75t_L g1421 ( 
.A1(n_1294),
.A2(n_1193),
.B(n_1093),
.C(n_1096),
.Y(n_1421)
);

INVx3_ASAP7_75t_SL g1422 ( 
.A(n_1247),
.Y(n_1422)
);

AOI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1284),
.A2(n_1127),
.B(n_1096),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1325),
.B(n_1110),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1246),
.B(n_1117),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1331),
.B(n_1144),
.Y(n_1426)
);

AO31x2_ASAP7_75t_L g1427 ( 
.A1(n_1298),
.A2(n_1117),
.A3(n_1211),
.B(n_1164),
.Y(n_1427)
);

AO22x2_ASAP7_75t_L g1428 ( 
.A1(n_1367),
.A2(n_1147),
.B1(n_1144),
.B2(n_1190),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1249),
.A2(n_1164),
.B(n_1098),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1235),
.A2(n_1098),
.B(n_1190),
.Y(n_1430)
);

OA21x2_ASAP7_75t_L g1431 ( 
.A1(n_1227),
.A2(n_225),
.B(n_223),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1321),
.A2(n_214),
.B(n_210),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1262),
.A2(n_208),
.B(n_207),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1252),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1319),
.A2(n_36),
.B(n_40),
.Y(n_1435)
);

NOR2xp67_ASAP7_75t_SL g1436 ( 
.A(n_1231),
.B(n_36),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1355),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1253),
.Y(n_1438)
);

OAI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1319),
.A2(n_47),
.B(n_48),
.Y(n_1439)
);

O2A1O1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1364),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1440)
);

A2O1A1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1282),
.A2(n_52),
.B(n_54),
.C(n_56),
.Y(n_1441)
);

NAND3xp33_ASAP7_75t_L g1442 ( 
.A(n_1305),
.B(n_59),
.C(n_60),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1301),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1339),
.A2(n_61),
.B(n_62),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1257),
.B(n_69),
.Y(n_1445)
);

AO21x1_ASAP7_75t_L g1446 ( 
.A1(n_1282),
.A2(n_72),
.B(n_74),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_SL g1447 ( 
.A1(n_1339),
.A2(n_76),
.B(n_77),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1256),
.B(n_76),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1267),
.A2(n_114),
.B(n_198),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1323),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_1450)
);

A2O1A1Ixp33_ASAP7_75t_L g1451 ( 
.A1(n_1352),
.A2(n_79),
.B(n_82),
.C(n_83),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1262),
.A2(n_127),
.B(n_89),
.Y(n_1452)
);

O2A1O1Ixp5_ASAP7_75t_SL g1453 ( 
.A1(n_1258),
.A2(n_83),
.B(n_90),
.C(n_94),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1276),
.Y(n_1454)
);

A2O1A1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1356),
.A2(n_98),
.B(n_100),
.C(n_113),
.Y(n_1455)
);

AOI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1270),
.A2(n_123),
.B(n_131),
.Y(n_1456)
);

AO31x2_ASAP7_75t_L g1457 ( 
.A1(n_1298),
.A2(n_136),
.A3(n_153),
.B(n_155),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1270),
.A2(n_161),
.B(n_172),
.Y(n_1458)
);

AOI21xp5_ASAP7_75t_L g1459 ( 
.A1(n_1272),
.A2(n_186),
.B(n_202),
.Y(n_1459)
);

A2O1A1Ixp33_ASAP7_75t_L g1460 ( 
.A1(n_1305),
.A2(n_1328),
.B(n_1308),
.C(n_1322),
.Y(n_1460)
);

NAND2x1p5_ASAP7_75t_L g1461 ( 
.A(n_1331),
.B(n_1242),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1259),
.B(n_1266),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1273),
.A2(n_1299),
.B(n_1274),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1273),
.A2(n_1274),
.B(n_1239),
.Y(n_1464)
);

OAI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1338),
.A2(n_1310),
.B(n_1316),
.Y(n_1465)
);

O2A1O1Ixp33_ASAP7_75t_SL g1466 ( 
.A1(n_1296),
.A2(n_1300),
.B(n_1297),
.C(n_1326),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_L g1467 ( 
.A(n_1287),
.B(n_1264),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1239),
.A2(n_1255),
.B(n_1366),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1325),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1283),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1285),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_L g1472 ( 
.A1(n_1336),
.A2(n_1292),
.B1(n_1353),
.B2(n_1290),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1271),
.B(n_1241),
.Y(n_1473)
);

NAND3xp33_ASAP7_75t_L g1474 ( 
.A(n_1361),
.B(n_1359),
.C(n_1337),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1248),
.B(n_1260),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1327),
.A2(n_1362),
.B1(n_1214),
.B2(n_1244),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1329),
.B(n_1347),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1366),
.A2(n_1361),
.B(n_1312),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1353),
.Y(n_1479)
);

NAND3x1_ASAP7_75t_L g1480 ( 
.A(n_1230),
.B(n_1351),
.C(n_1277),
.Y(n_1480)
);

NOR2xp67_ASAP7_75t_L g1481 ( 
.A(n_1358),
.B(n_1243),
.Y(n_1481)
);

AOI221xp5_ASAP7_75t_SL g1482 ( 
.A1(n_1344),
.A2(n_1309),
.B1(n_1341),
.B2(n_1332),
.C(n_1317),
.Y(n_1482)
);

BUFx10_ASAP7_75t_L g1483 ( 
.A(n_1243),
.Y(n_1483)
);

INVx5_ASAP7_75t_L g1484 ( 
.A(n_1293),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1318),
.A2(n_1354),
.B(n_1346),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1304),
.B(n_1311),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1344),
.A2(n_1220),
.B(n_1263),
.Y(n_1487)
);

INVx2_ASAP7_75t_SL g1488 ( 
.A(n_1314),
.Y(n_1488)
);

AOI21xp5_ASAP7_75t_L g1489 ( 
.A1(n_1220),
.A2(n_1216),
.B(n_1334),
.Y(n_1489)
);

INVx2_ASAP7_75t_SL g1490 ( 
.A(n_1287),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1313),
.B(n_1320),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1343),
.B(n_1307),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1268),
.B(n_1291),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1250),
.B(n_1269),
.Y(n_1494)
);

AO21x1_ASAP7_75t_L g1495 ( 
.A1(n_1236),
.A2(n_1350),
.B(n_1345),
.Y(n_1495)
);

NOR2xp67_ASAP7_75t_SL g1496 ( 
.A(n_1287),
.B(n_1342),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1221),
.A2(n_1261),
.B(n_1278),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1221),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1278),
.A2(n_1330),
.B(n_1293),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_L g1500 ( 
.A1(n_1330),
.A2(n_1067),
.B(n_1050),
.Y(n_1500)
);

INVx1_ASAP7_75t_SL g1501 ( 
.A(n_1330),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1303),
.Y(n_1502)
);

AOI21xp5_ASAP7_75t_L g1503 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_L g1504 ( 
.A(n_1229),
.B(n_727),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1223),
.A2(n_1265),
.B(n_1281),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1225),
.Y(n_1506)
);

BUFx12f_ASAP7_75t_L g1507 ( 
.A(n_1240),
.Y(n_1507)
);

AOI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1213),
.A2(n_757),
.B1(n_799),
.B2(n_727),
.Y(n_1508)
);

OAI21x1_ASAP7_75t_L g1509 ( 
.A1(n_1223),
.A2(n_1265),
.B(n_1281),
.Y(n_1509)
);

AOI21xp5_ASAP7_75t_L g1510 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1213),
.A2(n_1050),
.B1(n_1067),
.B2(n_1049),
.Y(n_1511)
);

NOR2x1_ASAP7_75t_SL g1512 ( 
.A(n_1242),
.B(n_1287),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1223),
.A2(n_1265),
.B(n_1281),
.Y(n_1513)
);

INVx5_ASAP7_75t_L g1514 ( 
.A(n_1301),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1279),
.B(n_1050),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1324),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1279),
.B(n_1050),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1279),
.B(n_1050),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1521)
);

AOI21xp5_ASAP7_75t_L g1522 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1279),
.B(n_1050),
.Y(n_1523)
);

AOI22xp33_ASAP7_75t_L g1524 ( 
.A1(n_1367),
.A2(n_890),
.B1(n_835),
.B2(n_765),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1226),
.A2(n_1067),
.B(n_1050),
.Y(n_1525)
);

OA21x2_ASAP7_75t_L g1526 ( 
.A1(n_1288),
.A2(n_1289),
.B(n_1226),
.Y(n_1526)
);

AOI221xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1213),
.A2(n_1305),
.B1(n_1349),
.B2(n_1361),
.C(n_1359),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1223),
.A2(n_1265),
.B(n_1281),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1504),
.A2(n_1508),
.B1(n_1371),
.B2(n_1511),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1507),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1462),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1462),
.Y(n_1532)
);

AO32x2_ASAP7_75t_L g1533 ( 
.A1(n_1371),
.A2(n_1511),
.A3(n_1472),
.B1(n_1397),
.B2(n_1450),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1381),
.Y(n_1534)
);

AO21x2_ASAP7_75t_L g1535 ( 
.A1(n_1383),
.A2(n_1487),
.B(n_1489),
.Y(n_1535)
);

AOI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1503),
.A2(n_1515),
.B(n_1510),
.Y(n_1536)
);

A2O1A1Ixp33_ASAP7_75t_L g1537 ( 
.A1(n_1391),
.A2(n_1400),
.B(n_1435),
.C(n_1439),
.Y(n_1537)
);

OAI21x1_ASAP7_75t_L g1538 ( 
.A1(n_1528),
.A2(n_1393),
.B(n_1423),
.Y(n_1538)
);

NAND2x1p5_ASAP7_75t_L g1539 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1539)
);

OAI21x1_ASAP7_75t_L g1540 ( 
.A1(n_1395),
.A2(n_1478),
.B(n_1388),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1484),
.B(n_1497),
.Y(n_1541)
);

OAI21x1_ASAP7_75t_SL g1542 ( 
.A1(n_1465),
.A2(n_1439),
.B(n_1435),
.Y(n_1542)
);

AOI221xp5_ASAP7_75t_SL g1543 ( 
.A1(n_1440),
.A2(n_1450),
.B1(n_1451),
.B2(n_1437),
.C(n_1397),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1500),
.A2(n_1387),
.B(n_1383),
.Y(n_1544)
);

CKINVDCx6p67_ASAP7_75t_R g1545 ( 
.A(n_1422),
.Y(n_1545)
);

OAI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1518),
.A2(n_1522),
.B(n_1521),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1419),
.A2(n_1370),
.B(n_1525),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1516),
.A2(n_1519),
.B1(n_1523),
.B2(n_1520),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1434),
.Y(n_1549)
);

INVx4_ASAP7_75t_L g1550 ( 
.A(n_1375),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1485),
.Y(n_1552)
);

A2O1A1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1444),
.A2(n_1527),
.B(n_1465),
.C(n_1474),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1438),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1415),
.A2(n_1394),
.B(n_1429),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1520),
.A2(n_1523),
.B1(n_1524),
.B2(n_1460),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1526),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1463),
.A2(n_1384),
.B(n_1417),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1413),
.A2(n_1464),
.B(n_1452),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1433),
.A2(n_1374),
.B(n_1432),
.Y(n_1560)
);

CKINVDCx8_ASAP7_75t_R g1561 ( 
.A(n_1454),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1470),
.Y(n_1562)
);

NAND3xp33_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1442),
.C(n_1444),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1468),
.Y(n_1564)
);

OAI21x1_ASAP7_75t_L g1565 ( 
.A1(n_1456),
.A2(n_1458),
.B(n_1419),
.Y(n_1565)
);

BUFx3_ASAP7_75t_L g1566 ( 
.A(n_1471),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1431),
.A2(n_1378),
.B(n_1453),
.Y(n_1567)
);

OAI21xp5_ASAP7_75t_L g1568 ( 
.A1(n_1402),
.A2(n_1404),
.B(n_1482),
.Y(n_1568)
);

OAI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1482),
.A2(n_1377),
.B(n_1472),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1372),
.A2(n_1430),
.B(n_1459),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1407),
.A2(n_1376),
.B1(n_1390),
.B2(n_1494),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1372),
.Y(n_1572)
);

INVxp67_ASAP7_75t_SL g1573 ( 
.A(n_1405),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1412),
.A2(n_1501),
.B1(n_1466),
.B2(n_1476),
.C(n_1441),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1409),
.A2(n_1373),
.B(n_1494),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1369),
.B(n_1469),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1449),
.A2(n_1411),
.B(n_1416),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1506),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1428),
.A2(n_1501),
.B1(n_1446),
.B2(n_1493),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1392),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1424),
.B(n_1498),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1582)
);

AOI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1477),
.A2(n_1418),
.B(n_1495),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1369),
.A2(n_1445),
.B1(n_1448),
.B2(n_1484),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1427),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1420),
.A2(n_1421),
.B(n_1403),
.Y(n_1586)
);

AO31x2_ASAP7_75t_L g1587 ( 
.A1(n_1418),
.A2(n_1477),
.A3(n_1486),
.B(n_1491),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1428),
.B(n_1398),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1497),
.B(n_1426),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1406),
.B(n_1401),
.Y(n_1590)
);

OR2x6_ASAP7_75t_L g1591 ( 
.A(n_1473),
.B(n_1408),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1496),
.B(n_1455),
.C(n_1436),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1426),
.B(n_1481),
.Y(n_1593)
);

BUFx3_ASAP7_75t_L g1594 ( 
.A(n_1385),
.Y(n_1594)
);

AO21x2_ASAP7_75t_L g1595 ( 
.A1(n_1486),
.A2(n_1491),
.B(n_1447),
.Y(n_1595)
);

OAI22x1_ASAP7_75t_L g1596 ( 
.A1(n_1502),
.A2(n_1480),
.B1(n_1380),
.B2(n_1488),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1386),
.A2(n_1414),
.B1(n_1502),
.B2(n_1443),
.Y(n_1597)
);

NAND3xp33_ASAP7_75t_L g1598 ( 
.A(n_1467),
.B(n_1410),
.C(n_1425),
.Y(n_1598)
);

BUFx2_ASAP7_75t_SL g1599 ( 
.A(n_1368),
.Y(n_1599)
);

BUFx12f_ASAP7_75t_L g1600 ( 
.A(n_1379),
.Y(n_1600)
);

OAI21xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1499),
.A2(n_1396),
.B(n_1389),
.Y(n_1601)
);

NAND2x1_ASAP7_75t_L g1602 ( 
.A(n_1443),
.B(n_1389),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1483),
.A2(n_1517),
.B1(n_1385),
.B2(n_1492),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_L g1604 ( 
.A1(n_1382),
.A2(n_1399),
.B(n_1490),
.Y(n_1604)
);

BUFx4f_ASAP7_75t_L g1605 ( 
.A(n_1385),
.Y(n_1605)
);

NAND2x1p5_ASAP7_75t_L g1606 ( 
.A(n_1514),
.B(n_1396),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1427),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1514),
.B(n_1517),
.Y(n_1608)
);

HB1xp67_ASAP7_75t_L g1609 ( 
.A(n_1427),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_SL g1610 ( 
.A1(n_1483),
.A2(n_1475),
.B1(n_1512),
.B2(n_1517),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1457),
.Y(n_1611)
);

AOI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1457),
.A2(n_1461),
.B(n_1379),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1457),
.B(n_1215),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1462),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_SL g1617 ( 
.A1(n_1504),
.A2(n_1213),
.B(n_1439),
.C(n_1435),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1462),
.Y(n_1618)
);

OAI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1371),
.A2(n_1279),
.B1(n_765),
.B2(n_1360),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1371),
.A2(n_890),
.B1(n_765),
.B2(n_1524),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1508),
.A2(n_890),
.B1(n_884),
.B2(n_1371),
.C(n_1184),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1526),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1485),
.Y(n_1625)
);

OAI21x1_ASAP7_75t_SL g1626 ( 
.A1(n_1465),
.A2(n_1371),
.B(n_1435),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1462),
.Y(n_1627)
);

OAI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1504),
.A2(n_1213),
.B1(n_1508),
.B2(n_1371),
.Y(n_1628)
);

OAI21x1_ASAP7_75t_L g1629 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_SL g1630 ( 
.A1(n_1511),
.A2(n_1460),
.B(n_1400),
.C(n_1371),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1503),
.A2(n_1515),
.B(n_1510),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1504),
.A2(n_1213),
.B1(n_1508),
.B2(n_1371),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1371),
.A2(n_1213),
.B(n_1184),
.Y(n_1633)
);

INVx1_ASAP7_75t_SL g1634 ( 
.A(n_1422),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1479),
.Y(n_1635)
);

O2A1O1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1371),
.A2(n_1511),
.B(n_1213),
.C(n_1184),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1503),
.A2(n_1515),
.B(n_1510),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1503),
.A2(n_1515),
.B(n_1510),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1485),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_1514),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1507),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1485),
.Y(n_1643)
);

OAI21x1_ASAP7_75t_L g1644 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1462),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1407),
.B(n_1286),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1488),
.B(n_1215),
.Y(n_1647)
);

NAND2x1p5_ASAP7_75t_L g1648 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1648)
);

NAND2x1p5_ASAP7_75t_L g1649 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1649)
);

NOR2xp33_ASAP7_75t_L g1650 ( 
.A(n_1371),
.B(n_1504),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1371),
.A2(n_890),
.B1(n_765),
.B2(n_1524),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1383),
.A2(n_1487),
.B(n_1226),
.Y(n_1652)
);

INVx6_ASAP7_75t_L g1653 ( 
.A(n_1483),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_SL g1655 ( 
.A1(n_1371),
.A2(n_1367),
.B1(n_835),
.B2(n_619),
.Y(n_1655)
);

AOI21xp33_ASAP7_75t_L g1656 ( 
.A1(n_1527),
.A2(n_1184),
.B(n_1306),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1484),
.B(n_1497),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1375),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1371),
.A2(n_890),
.B1(n_765),
.B2(n_1524),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1462),
.Y(n_1660)
);

AO31x2_ASAP7_75t_L g1661 ( 
.A1(n_1383),
.A2(n_1226),
.A3(n_1405),
.B(n_1487),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1485),
.Y(n_1662)
);

AOI22xp33_ASAP7_75t_L g1663 ( 
.A1(n_1371),
.A2(n_890),
.B1(n_765),
.B2(n_1524),
.Y(n_1663)
);

AOI221xp5_ASAP7_75t_L g1664 ( 
.A1(n_1371),
.A2(n_890),
.B1(n_884),
.B2(n_1113),
.C(n_1511),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1665)
);

AO31x2_ASAP7_75t_L g1666 ( 
.A1(n_1383),
.A2(n_1226),
.A3(n_1405),
.B(n_1487),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1484),
.B(n_1497),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1485),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1371),
.A2(n_1367),
.B1(n_835),
.B2(n_619),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1485),
.Y(n_1672)
);

AOI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1423),
.A2(n_1289),
.B(n_1487),
.Y(n_1673)
);

OAI21x1_ASAP7_75t_SL g1674 ( 
.A1(n_1465),
.A2(n_1371),
.B(n_1435),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1676)
);

OA21x2_ASAP7_75t_L g1677 ( 
.A1(n_1393),
.A2(n_1509),
.B(n_1505),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1369),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1485),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1479),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1485),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1393),
.A2(n_1509),
.B(n_1505),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1375),
.Y(n_1686)
);

INVx4_ASAP7_75t_L g1687 ( 
.A(n_1422),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1507),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1516),
.B(n_1519),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1407),
.B(n_1286),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1407),
.B(n_1286),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1504),
.A2(n_1371),
.B1(n_890),
.B2(n_1224),
.Y(n_1692)
);

NAND2x1_ASAP7_75t_L g1693 ( 
.A(n_1443),
.B(n_1378),
.Y(n_1693)
);

OAI21x1_ASAP7_75t_L g1694 ( 
.A1(n_1505),
.A2(n_1513),
.B(n_1509),
.Y(n_1694)
);

AOI222xp33_ASAP7_75t_L g1695 ( 
.A1(n_1524),
.A2(n_619),
.B1(n_835),
.B2(n_611),
.C1(n_1044),
.C2(n_1113),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1504),
.A2(n_1213),
.B1(n_1508),
.B2(n_1371),
.Y(n_1696)
);

NAND2x1p5_ASAP7_75t_L g1697 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1484),
.B(n_1497),
.Y(n_1698)
);

O2A1O1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1371),
.A2(n_1511),
.B(n_1213),
.C(n_1184),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1504),
.A2(n_1213),
.B1(n_1508),
.B2(n_1371),
.Y(n_1700)
);

XNOR2xp5_ASAP7_75t_L g1701 ( 
.A(n_1476),
.B(n_620),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1503),
.A2(n_1515),
.B(n_1510),
.Y(n_1702)
);

NAND2x1p5_ASAP7_75t_L g1703 ( 
.A(n_1484),
.B(n_1514),
.Y(n_1703)
);

INVx3_ASAP7_75t_SL g1704 ( 
.A(n_1422),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1534),
.Y(n_1706)
);

BUFx2_ASAP7_75t_L g1707 ( 
.A(n_1566),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1615),
.B(n_1616),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1665),
.B(n_1668),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1675),
.B(n_1689),
.Y(n_1711)
);

AND2x2_ASAP7_75t_SL g1712 ( 
.A(n_1650),
.B(n_1664),
.Y(n_1712)
);

AND2x4_ASAP7_75t_L g1713 ( 
.A(n_1541),
.B(n_1657),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1650),
.B(n_1590),
.Y(n_1714)
);

AND2x4_ASAP7_75t_L g1715 ( 
.A(n_1541),
.B(n_1657),
.Y(n_1715)
);

AOI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1628),
.A2(n_1632),
.B(n_1700),
.C(n_1696),
.Y(n_1716)
);

AND2x2_ASAP7_75t_SL g1717 ( 
.A(n_1692),
.B(n_1622),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1572),
.Y(n_1718)
);

AOI21x1_ASAP7_75t_SL g1719 ( 
.A1(n_1564),
.A2(n_1690),
.B(n_1646),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1667),
.B(n_1698),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1566),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1536),
.A2(n_1637),
.B(n_1631),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1678),
.B(n_1633),
.Y(n_1723)
);

OR2x6_ASAP7_75t_L g1724 ( 
.A(n_1667),
.B(n_1698),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1588),
.B(n_1691),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1576),
.B(n_1571),
.Y(n_1726)
);

AOI31xp33_ASAP7_75t_L g1727 ( 
.A1(n_1655),
.A2(n_1671),
.A3(n_1529),
.B(n_1695),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1655),
.A2(n_1671),
.B1(n_1623),
.B2(n_1663),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1622),
.A2(n_1651),
.B1(n_1659),
.B2(n_1663),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1678),
.B(n_1531),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1580),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1572),
.Y(n_1732)
);

INVx8_ASAP7_75t_L g1733 ( 
.A(n_1593),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1636),
.B(n_1699),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1549),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1635),
.B(n_1682),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1636),
.B(n_1699),
.Y(n_1737)
);

O2A1O1Ixp33_ASAP7_75t_L g1738 ( 
.A1(n_1617),
.A2(n_1619),
.B(n_1630),
.C(n_1656),
.Y(n_1738)
);

BUFx3_ASAP7_75t_L g1739 ( 
.A(n_1608),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1532),
.B(n_1614),
.Y(n_1740)
);

OA21x2_ASAP7_75t_L g1741 ( 
.A1(n_1536),
.A2(n_1637),
.B(n_1631),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1579),
.B(n_1554),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1661),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1579),
.B(n_1562),
.Y(n_1744)
);

OA21x2_ASAP7_75t_L g1745 ( 
.A1(n_1639),
.A2(n_1702),
.B(n_1540),
.Y(n_1745)
);

OAI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1651),
.A2(n_1659),
.B1(n_1619),
.B2(n_1537),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1533),
.B(n_1578),
.Y(n_1747)
);

NOR2xp67_ASAP7_75t_L g1748 ( 
.A(n_1550),
.B(n_1687),
.Y(n_1748)
);

O2A1O1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1630),
.A2(n_1537),
.B(n_1553),
.C(n_1674),
.Y(n_1749)
);

O2A1O1Ixp5_ASAP7_75t_L g1750 ( 
.A1(n_1568),
.A2(n_1553),
.B(n_1569),
.C(n_1563),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1556),
.A2(n_1592),
.B1(n_1574),
.B2(n_1658),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1618),
.B(n_1627),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1686),
.A2(n_1550),
.B1(n_1591),
.B2(n_1634),
.Y(n_1753)
);

INVxp67_ASAP7_75t_L g1754 ( 
.A(n_1647),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1645),
.B(n_1660),
.Y(n_1755)
);

OAI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1591),
.A2(n_1584),
.B1(n_1561),
.B2(n_1701),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1543),
.A2(n_1577),
.B(n_1573),
.C(n_1533),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1591),
.A2(n_1584),
.B1(n_1704),
.B2(n_1545),
.Y(n_1758)
);

AND2x4_ASAP7_75t_L g1759 ( 
.A(n_1589),
.B(n_1613),
.Y(n_1759)
);

AOI21x1_ASAP7_75t_SL g1760 ( 
.A1(n_1557),
.A2(n_1624),
.B(n_1704),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_SL g1761 ( 
.A1(n_1539),
.A2(n_1703),
.B(n_1697),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1599),
.Y(n_1762)
);

AOI21x1_ASAP7_75t_SL g1763 ( 
.A1(n_1600),
.A2(n_1626),
.B(n_1687),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1612),
.B(n_1641),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1598),
.B(n_1603),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1575),
.A2(n_1693),
.B1(n_1605),
.B2(n_1533),
.Y(n_1766)
);

AOI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1542),
.A2(n_1583),
.B1(n_1596),
.B2(n_1546),
.C(n_1611),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1533),
.B(n_1594),
.Y(n_1768)
);

OA21x2_ASAP7_75t_L g1769 ( 
.A1(n_1538),
.A2(n_1586),
.B(n_1558),
.Y(n_1769)
);

O2A1O1Ixp33_ASAP7_75t_L g1770 ( 
.A1(n_1575),
.A2(n_1597),
.B(n_1594),
.C(n_1608),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_SL g1771 ( 
.A(n_1641),
.B(n_1595),
.Y(n_1771)
);

AOI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1565),
.A2(n_1586),
.B(n_1652),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1539),
.A2(n_1703),
.B(n_1697),
.Y(n_1773)
);

O2A1O1Ixp33_ASAP7_75t_L g1774 ( 
.A1(n_1602),
.A2(n_1601),
.B(n_1606),
.C(n_1604),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1605),
.B(n_1595),
.Y(n_1775)
);

O2A1O1Ixp5_ASAP7_75t_L g1776 ( 
.A1(n_1673),
.A2(n_1640),
.B(n_1643),
.C(n_1662),
.Y(n_1776)
);

INVxp67_ASAP7_75t_SL g1777 ( 
.A(n_1547),
.Y(n_1777)
);

O2A1O1Ixp5_ASAP7_75t_L g1778 ( 
.A1(n_1552),
.A2(n_1625),
.B(n_1683),
.C(n_1672),
.Y(n_1778)
);

OAI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1606),
.A2(n_1653),
.B1(n_1610),
.B2(n_1530),
.Y(n_1779)
);

HB1xp67_ASAP7_75t_L g1780 ( 
.A(n_1666),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1653),
.A2(n_1610),
.B1(n_1642),
.B2(n_1547),
.Y(n_1781)
);

AOI21x1_ASAP7_75t_SL g1782 ( 
.A1(n_1585),
.A2(n_1607),
.B(n_1609),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1570),
.A2(n_1567),
.B(n_1607),
.C(n_1585),
.Y(n_1783)
);

O2A1O1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1547),
.A2(n_1609),
.B(n_1535),
.C(n_1652),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1582),
.A2(n_1649),
.B1(n_1648),
.B2(n_1688),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1587),
.B(n_1666),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1582),
.A2(n_1648),
.B1(n_1649),
.B2(n_1544),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1677),
.A2(n_1684),
.B1(n_1679),
.B2(n_1672),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1677),
.A2(n_1684),
.B(n_1694),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1560),
.A2(n_1559),
.B(n_1555),
.C(n_1552),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1666),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1677),
.B(n_1684),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1625),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1629),
.B(n_1638),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1670),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1644),
.B(n_1654),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1669),
.A2(n_1676),
.B(n_1680),
.C(n_1681),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1685),
.B(n_1581),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1801)
);

BUFx8_ASAP7_75t_L g1802 ( 
.A(n_1688),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1590),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1580),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1534),
.Y(n_1808)
);

OAI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1650),
.A2(n_1692),
.B1(n_1664),
.B2(n_1671),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1633),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_SL g1811 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1537),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_SL g1812 ( 
.A1(n_1551),
.A2(n_1376),
.B(n_1390),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_L g1813 ( 
.A1(n_1650),
.A2(n_1692),
.B1(n_1664),
.B2(n_1671),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1814)
);

AOI21x1_ASAP7_75t_SL g1815 ( 
.A1(n_1551),
.A2(n_1376),
.B(n_1390),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1817)
);

NOR2xp67_ASAP7_75t_L g1818 ( 
.A(n_1550),
.B(n_1687),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1534),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1820)
);

OAI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1650),
.A2(n_1692),
.B1(n_1664),
.B2(n_1671),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_SL g1823 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1537),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1633),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1534),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1534),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1541),
.B(n_1657),
.Y(n_1829)
);

AOI21xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1537),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1581),
.B(n_1590),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1534),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1534),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_SL g1834 ( 
.A1(n_1650),
.A2(n_1671),
.B1(n_1655),
.B2(n_1628),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1572),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1636),
.A2(n_1699),
.B(n_1633),
.Y(n_1836)
);

BUFx3_ASAP7_75t_L g1837 ( 
.A(n_1566),
.Y(n_1837)
);

OAI22xp5_ASAP7_75t_L g1838 ( 
.A1(n_1650),
.A2(n_1692),
.B1(n_1664),
.B2(n_1671),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1839)
);

O2A1O1Ixp5_ASAP7_75t_L g1840 ( 
.A1(n_1650),
.A2(n_1633),
.B(n_1628),
.C(n_1632),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1650),
.A2(n_1692),
.B1(n_1664),
.B2(n_1671),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1572),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1551),
.B(n_1615),
.Y(n_1844)
);

O2A1O1Ixp5_ASAP7_75t_L g1845 ( 
.A1(n_1650),
.A2(n_1633),
.B(n_1628),
.C(n_1632),
.Y(n_1845)
);

AOI21x1_ASAP7_75t_SL g1846 ( 
.A1(n_1551),
.A2(n_1376),
.B(n_1390),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1548),
.B(n_1551),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1848)
);

OAI31xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1650),
.A2(n_1632),
.A3(n_1696),
.B(n_1628),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1533),
.B(n_1534),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1786),
.B(n_1743),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1747),
.B(n_1843),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1706),
.Y(n_1853)
);

OR2x6_ASAP7_75t_L g1854 ( 
.A(n_1724),
.B(n_1759),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1712),
.Y(n_1855)
);

AOI21x1_ASAP7_75t_L g1856 ( 
.A1(n_1789),
.A2(n_1813),
.B(n_1809),
.Y(n_1856)
);

AO21x2_ASAP7_75t_L g1857 ( 
.A1(n_1772),
.A2(n_1783),
.B(n_1757),
.Y(n_1857)
);

AO21x2_ASAP7_75t_L g1858 ( 
.A1(n_1783),
.A2(n_1757),
.B(n_1777),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1718),
.Y(n_1859)
);

AO21x2_ASAP7_75t_L g1860 ( 
.A1(n_1788),
.A2(n_1784),
.B(n_1790),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1759),
.B(n_1713),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1713),
.B(n_1715),
.Y(n_1862)
);

BUFx3_ASAP7_75t_L g1863 ( 
.A(n_1721),
.Y(n_1863)
);

OA21x2_ASAP7_75t_L g1864 ( 
.A1(n_1776),
.A2(n_1790),
.B(n_1767),
.Y(n_1864)
);

INVx3_ASAP7_75t_L g1865 ( 
.A(n_1792),
.Y(n_1865)
);

AOI222xp33_ASAP7_75t_L g1866 ( 
.A1(n_1834),
.A2(n_1728),
.B1(n_1821),
.B2(n_1841),
.C1(n_1838),
.C2(n_1712),
.Y(n_1866)
);

INVx2_ASAP7_75t_SL g1867 ( 
.A(n_1775),
.Y(n_1867)
);

INVx3_ASAP7_75t_L g1868 ( 
.A(n_1794),
.Y(n_1868)
);

OAI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1716),
.A2(n_1727),
.B1(n_1714),
.B2(n_1737),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1732),
.Y(n_1870)
);

INVx3_ASAP7_75t_L g1871 ( 
.A(n_1795),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1705),
.B(n_1814),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1735),
.Y(n_1873)
);

INVx1_ASAP7_75t_SL g1874 ( 
.A(n_1721),
.Y(n_1874)
);

AOI222xp33_ASAP7_75t_L g1875 ( 
.A1(n_1717),
.A2(n_1729),
.B1(n_1746),
.B2(n_1734),
.C1(n_1804),
.C2(n_1751),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1816),
.B(n_1820),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1732),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1780),
.B(n_1747),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1808),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1843),
.B(n_1848),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_L g1881 ( 
.A(n_1824),
.B(n_1825),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1819),
.Y(n_1882)
);

AO21x2_ASAP7_75t_L g1883 ( 
.A1(n_1810),
.A2(n_1826),
.B(n_1836),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1839),
.B(n_1847),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1827),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1848),
.B(n_1850),
.Y(n_1886)
);

INVx3_ASAP7_75t_L g1887 ( 
.A(n_1797),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1778),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1717),
.A2(n_1756),
.B1(n_1726),
.B2(n_1768),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1850),
.B(n_1835),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1828),
.Y(n_1891)
);

INVx1_ASAP7_75t_SL g1892 ( 
.A(n_1837),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1832),
.Y(n_1893)
);

AO21x2_ASAP7_75t_L g1894 ( 
.A1(n_1811),
.A2(n_1823),
.B(n_1830),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1791),
.B(n_1799),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1723),
.B(n_1849),
.Y(n_1896)
);

AO21x2_ASAP7_75t_L g1897 ( 
.A1(n_1811),
.A2(n_1823),
.B(n_1771),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1833),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1842),
.B(n_1730),
.Y(n_1899)
);

AOI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1742),
.A2(n_1744),
.B1(n_1725),
.B2(n_1765),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1791),
.B(n_1722),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1722),
.B(n_1741),
.Y(n_1902)
);

OA21x2_ASAP7_75t_L g1903 ( 
.A1(n_1750),
.A2(n_1845),
.B(n_1840),
.Y(n_1903)
);

BUFx3_ASAP7_75t_L g1904 ( 
.A(n_1707),
.Y(n_1904)
);

OA21x2_ASAP7_75t_L g1905 ( 
.A1(n_1798),
.A2(n_1793),
.B(n_1796),
.Y(n_1905)
);

AOI21x1_ASAP7_75t_L g1906 ( 
.A1(n_1781),
.A2(n_1758),
.B(n_1766),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1740),
.Y(n_1907)
);

AO21x2_ASAP7_75t_L g1908 ( 
.A1(n_1738),
.A2(n_1787),
.B(n_1749),
.Y(n_1908)
);

AO21x2_ASAP7_75t_L g1909 ( 
.A1(n_1764),
.A2(n_1753),
.B(n_1709),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1762),
.B(n_1731),
.Y(n_1910)
);

AO21x2_ASAP7_75t_L g1911 ( 
.A1(n_1764),
.A2(n_1708),
.B(n_1711),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1752),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1755),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_1741),
.Y(n_1914)
);

BUFx2_ASAP7_75t_L g1915 ( 
.A(n_1764),
.Y(n_1915)
);

OA21x2_ASAP7_75t_L g1916 ( 
.A1(n_1796),
.A2(n_1829),
.B(n_1720),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1769),
.Y(n_1917)
);

AO21x2_ASAP7_75t_L g1918 ( 
.A1(n_1770),
.A2(n_1782),
.B(n_1779),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1844),
.B(n_1710),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1745),
.B(n_1805),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1745),
.B(n_1803),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1774),
.Y(n_1922)
);

INVx2_ASAP7_75t_SL g1923 ( 
.A(n_1904),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1880),
.B(n_1801),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1870),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1880),
.B(n_1806),
.Y(n_1926)
);

OR2x6_ASAP7_75t_L g1927 ( 
.A(n_1854),
.B(n_1773),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1886),
.B(n_1920),
.Y(n_1928)
);

INVx3_ASAP7_75t_SL g1929 ( 
.A(n_1855),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1870),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1886),
.B(n_1800),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1886),
.B(n_1817),
.Y(n_1932)
);

OAI221xp5_ASAP7_75t_L g1933 ( 
.A1(n_1866),
.A2(n_1754),
.B1(n_1818),
.B2(n_1748),
.C(n_1785),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1869),
.A2(n_1831),
.B1(n_1822),
.B2(n_1736),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1920),
.B(n_1760),
.Y(n_1935)
);

AOI33xp33_ASAP7_75t_L g1936 ( 
.A1(n_1889),
.A2(n_1815),
.A3(n_1812),
.B1(n_1846),
.B2(n_1763),
.B3(n_1719),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1881),
.B(n_1739),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1881),
.B(n_1739),
.Y(n_1938)
);

INVx4_ASAP7_75t_L g1939 ( 
.A(n_1894),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1877),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1869),
.A2(n_1733),
.B1(n_1731),
.B2(n_1807),
.Y(n_1941)
);

NAND4xp25_ASAP7_75t_L g1942 ( 
.A(n_1866),
.B(n_1875),
.C(n_1896),
.D(n_1884),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1890),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1890),
.Y(n_1944)
);

BUFx5_ASAP7_75t_L g1945 ( 
.A(n_1901),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1872),
.B(n_1761),
.Y(n_1946)
);

BUFx3_ASAP7_75t_L g1947 ( 
.A(n_1863),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1859),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1859),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1876),
.B(n_1733),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1921),
.B(n_1761),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1855),
.B(n_1807),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1878),
.B(n_1802),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1853),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1878),
.B(n_1802),
.Y(n_1955)
);

AO21x2_ASAP7_75t_L g1956 ( 
.A1(n_1888),
.A2(n_1802),
.B(n_1917),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1876),
.B(n_1884),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1861),
.B(n_1862),
.Y(n_1958)
);

AND2x4_ASAP7_75t_L g1959 ( 
.A(n_1861),
.B(n_1862),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1883),
.B(n_1896),
.Y(n_1960)
);

OAI211xp5_ASAP7_75t_L g1961 ( 
.A1(n_1875),
.A2(n_1855),
.B(n_1856),
.C(n_1903),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1883),
.B(n_1911),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1878),
.B(n_1852),
.Y(n_1963)
);

AOI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1883),
.A2(n_1889),
.B1(n_1900),
.B2(n_1922),
.C(n_1855),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_SL g1965 ( 
.A(n_1894),
.B(n_1897),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_L g1966 ( 
.A(n_1960),
.B(n_1922),
.C(n_1903),
.Y(n_1966)
);

AOI33xp33_ASAP7_75t_L g1967 ( 
.A1(n_1964),
.A2(n_1900),
.A3(n_1913),
.B1(n_1912),
.B2(n_1882),
.B3(n_1879),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1957),
.B(n_1883),
.Y(n_1968)
);

NAND3xp33_ASAP7_75t_L g1969 ( 
.A(n_1961),
.B(n_1903),
.C(n_1864),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1953),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1942),
.A2(n_1894),
.B1(n_1908),
.B2(n_1903),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1958),
.Y(n_1972)
);

BUFx3_ASAP7_75t_L g1973 ( 
.A(n_1953),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1963),
.B(n_1865),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1963),
.B(n_1928),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1942),
.A2(n_1894),
.B1(n_1908),
.B2(n_1918),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1925),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1958),
.B(n_1862),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1925),
.Y(n_1979)
);

OAI31xp33_ASAP7_75t_L g1980 ( 
.A1(n_1934),
.A2(n_1851),
.A3(n_1856),
.B(n_1915),
.Y(n_1980)
);

NAND2xp33_ASAP7_75t_SL g1981 ( 
.A(n_1929),
.B(n_1897),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1930),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1955),
.Y(n_1983)
);

OAI33xp33_ASAP7_75t_L g1984 ( 
.A1(n_1934),
.A2(n_1919),
.A3(n_1907),
.B1(n_1899),
.B2(n_1912),
.B3(n_1913),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1956),
.A2(n_1908),
.B1(n_1918),
.B2(n_1909),
.Y(n_1985)
);

CKINVDCx20_ASAP7_75t_R g1986 ( 
.A(n_1955),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1930),
.Y(n_1987)
);

BUFx3_ASAP7_75t_L g1988 ( 
.A(n_1947),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1946),
.Y(n_1989)
);

AOI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1962),
.A2(n_1897),
.B(n_1903),
.Y(n_1990)
);

NOR2x1_ASAP7_75t_SL g1991 ( 
.A(n_1927),
.B(n_1897),
.Y(n_1991)
);

OAI22xp33_ASAP7_75t_L g1992 ( 
.A1(n_1946),
.A2(n_1906),
.B1(n_1916),
.B2(n_1854),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1937),
.B(n_1904),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1940),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1940),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1938),
.B(n_1910),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1924),
.B(n_1911),
.Y(n_1997)
);

OAI211xp5_ASAP7_75t_L g1998 ( 
.A1(n_1941),
.A2(n_1906),
.B(n_1864),
.C(n_1905),
.Y(n_1998)
);

AOI22xp33_ASAP7_75t_L g1999 ( 
.A1(n_1956),
.A2(n_1908),
.B1(n_1918),
.B2(n_1909),
.Y(n_1999)
);

OAI211xp5_ASAP7_75t_L g2000 ( 
.A1(n_1941),
.A2(n_1864),
.B(n_1905),
.C(n_1902),
.Y(n_2000)
);

AOI211xp5_ASAP7_75t_SL g2001 ( 
.A1(n_1933),
.A2(n_1871),
.B(n_1887),
.C(n_1868),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1943),
.Y(n_2002)
);

AND2x4_ASAP7_75t_L g2003 ( 
.A(n_1958),
.B(n_1862),
.Y(n_2003)
);

AOI221xp5_ASAP7_75t_SL g2004 ( 
.A1(n_1935),
.A2(n_1874),
.B1(n_1892),
.B2(n_1895),
.C(n_1893),
.Y(n_2004)
);

AOI22xp33_ASAP7_75t_L g2005 ( 
.A1(n_1956),
.A2(n_1918),
.B1(n_1909),
.B2(n_1857),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1928),
.B(n_1865),
.Y(n_2006)
);

NAND4xp25_ASAP7_75t_L g2007 ( 
.A(n_1936),
.B(n_1935),
.C(n_1949),
.D(n_1948),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1950),
.B(n_1919),
.Y(n_2008)
);

BUFx3_ASAP7_75t_L g2009 ( 
.A(n_1947),
.Y(n_2009)
);

NOR2x1_ASAP7_75t_L g2010 ( 
.A(n_1952),
.B(n_1863),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1956),
.A2(n_1857),
.B1(n_1858),
.B2(n_1867),
.Y(n_2011)
);

AO21x2_ASAP7_75t_L g2012 ( 
.A1(n_1965),
.A2(n_1888),
.B(n_1860),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1951),
.A2(n_1857),
.B1(n_1858),
.B2(n_1867),
.Y(n_2013)
);

AOI33xp33_ASAP7_75t_L g2014 ( 
.A1(n_1944),
.A2(n_1882),
.A3(n_1885),
.B1(n_1898),
.B2(n_1873),
.B3(n_1891),
.Y(n_2014)
);

OA21x2_ASAP7_75t_L g2015 ( 
.A1(n_1990),
.A2(n_1917),
.B(n_1914),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1977),
.Y(n_2016)
);

HB1xp67_ASAP7_75t_L g2017 ( 
.A(n_1977),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1979),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1979),
.Y(n_2019)
);

NAND3xp33_ASAP7_75t_SL g2020 ( 
.A(n_1971),
.B(n_1939),
.C(n_1892),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1982),
.Y(n_2021)
);

HB1xp67_ASAP7_75t_L g2022 ( 
.A(n_1982),
.Y(n_2022)
);

INVx4_ASAP7_75t_L g2023 ( 
.A(n_1988),
.Y(n_2023)
);

INVx3_ASAP7_75t_L g2024 ( 
.A(n_1972),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_SL g2025 ( 
.A1(n_1969),
.A2(n_1965),
.B(n_1905),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1978),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1968),
.B(n_1944),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_1981),
.Y(n_2028)
);

AOI21xp33_ASAP7_75t_SL g2029 ( 
.A1(n_1970),
.A2(n_1929),
.B(n_1923),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1975),
.B(n_2006),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1987),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1975),
.B(n_1945),
.Y(n_2032)
);

BUFx2_ASAP7_75t_L g2033 ( 
.A(n_1981),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_2014),
.B(n_1954),
.Y(n_2034)
);

AOI21xp5_ASAP7_75t_SL g2035 ( 
.A1(n_1998),
.A2(n_1905),
.B(n_1939),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_1988),
.Y(n_2036)
);

AOI21xp33_ASAP7_75t_SL g2037 ( 
.A1(n_1970),
.A2(n_1929),
.B(n_1923),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2006),
.B(n_1945),
.Y(n_2038)
);

INVx4_ASAP7_75t_L g2039 ( 
.A(n_2009),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1986),
.Y(n_2040)
);

AO21x2_ASAP7_75t_L g2041 ( 
.A1(n_1966),
.A2(n_1860),
.B(n_1858),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_2003),
.B(n_1959),
.Y(n_2042)
);

HB1xp67_ASAP7_75t_L g2043 ( 
.A(n_1994),
.Y(n_2043)
);

AND3x2_ASAP7_75t_L g2044 ( 
.A(n_2035),
.B(n_1980),
.C(n_1989),
.Y(n_2044)
);

AOI31xp33_ASAP7_75t_L g2045 ( 
.A1(n_2020),
.A2(n_1976),
.A3(n_2000),
.B(n_2001),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2032),
.B(n_2004),
.Y(n_2046)
);

NOR2x1_ASAP7_75t_L g2047 ( 
.A(n_2023),
.B(n_2007),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_2017),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2034),
.B(n_1997),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_2034),
.B(n_1995),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2017),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2030),
.B(n_1974),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_2041),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_2030),
.B(n_1974),
.Y(n_2054)
);

BUFx2_ASAP7_75t_SL g2055 ( 
.A(n_2040),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_2041),
.A2(n_1999),
.B1(n_1985),
.B2(n_2005),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_2030),
.B(n_2003),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2022),
.B(n_1967),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_2038),
.B(n_2003),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_2041),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_2022),
.Y(n_2061)
);

HB1xp67_ASAP7_75t_L g2062 ( 
.A(n_2043),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2043),
.Y(n_2063)
);

INVx1_ASAP7_75t_SL g2064 ( 
.A(n_2040),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2016),
.Y(n_2065)
);

AND2x2_ASAP7_75t_L g2066 ( 
.A(n_2038),
.B(n_1993),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2016),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_2041),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2016),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2041),
.A2(n_2013),
.B1(n_1984),
.B2(n_1858),
.Y(n_2070)
);

NAND4xp25_ASAP7_75t_L g2071 ( 
.A(n_2036),
.B(n_2010),
.C(n_2011),
.D(n_1973),
.Y(n_2071)
);

INVxp67_ASAP7_75t_L g2072 ( 
.A(n_2036),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2015),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_2018),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2018),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2015),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2026),
.B(n_1983),
.Y(n_2077)
);

BUFx3_ASAP7_75t_L g2078 ( 
.A(n_2028),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2018),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_2027),
.B(n_2002),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2019),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2061),
.Y(n_2082)
);

NOR2x1_ASAP7_75t_L g2083 ( 
.A(n_2078),
.B(n_2023),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2058),
.B(n_2027),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_2057),
.B(n_2042),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2053),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2057),
.B(n_2042),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2072),
.B(n_2008),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2053),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2057),
.B(n_2042),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2053),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2061),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2077),
.B(n_2042),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2072),
.B(n_1926),
.Y(n_2094)
);

INVxp67_ASAP7_75t_SL g2095 ( 
.A(n_2078),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2077),
.B(n_2042),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2062),
.Y(n_2097)
);

NAND2x1_ASAP7_75t_L g2098 ( 
.A(n_2047),
.B(n_2026),
.Y(n_2098)
);

NOR2x1_ASAP7_75t_L g2099 ( 
.A(n_2078),
.B(n_2023),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2062),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2050),
.B(n_1931),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_2050),
.B(n_2064),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_2077),
.B(n_2042),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2064),
.B(n_2058),
.Y(n_2104)
);

INVx1_ASAP7_75t_SL g2105 ( 
.A(n_2055),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2070),
.B(n_1931),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2047),
.B(n_2023),
.Y(n_2107)
);

OAI21xp5_ASAP7_75t_SL g2108 ( 
.A1(n_2044),
.A2(n_2020),
.B(n_2029),
.Y(n_2108)
);

OAI21xp5_ASAP7_75t_L g2109 ( 
.A1(n_2045),
.A2(n_2025),
.B(n_2028),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2065),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2052),
.B(n_2023),
.Y(n_2111)
);

AOI21xp5_ASAP7_75t_L g2112 ( 
.A1(n_2045),
.A2(n_1992),
.B(n_2028),
.Y(n_2112)
);

NOR2xp67_ASAP7_75t_L g2113 ( 
.A(n_2071),
.B(n_2026),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_2078),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2070),
.B(n_1932),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2049),
.B(n_2027),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_2048),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2052),
.B(n_2039),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_SL g2119 ( 
.A1(n_2044),
.A2(n_2033),
.B(n_1991),
.Y(n_2119)
);

OR2x2_ASAP7_75t_L g2120 ( 
.A(n_2049),
.B(n_2019),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2052),
.B(n_2039),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2065),
.Y(n_2122)
);

NOR2x1_ASAP7_75t_L g2123 ( 
.A(n_2055),
.B(n_2039),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2067),
.Y(n_2124)
);

NOR4xp25_ASAP7_75t_L g2125 ( 
.A(n_2071),
.B(n_2024),
.C(n_2031),
.D(n_2021),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2110),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2110),
.Y(n_2127)
);

AND2x2_ASAP7_75t_L g2128 ( 
.A(n_2111),
.B(n_2054),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_2125),
.B(n_2048),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2114),
.Y(n_2130)
);

INVx1_ASAP7_75t_SL g2131 ( 
.A(n_2105),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2122),
.Y(n_2132)
);

AOI221xp5_ASAP7_75t_L g2133 ( 
.A1(n_2112),
.A2(n_2056),
.B1(n_2049),
.B2(n_2053),
.C(n_2068),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_L g2134 ( 
.A(n_2088),
.B(n_1986),
.Y(n_2134)
);

HB1xp67_ASAP7_75t_L g2135 ( 
.A(n_2114),
.Y(n_2135)
);

INVx1_ASAP7_75t_SL g2136 ( 
.A(n_2123),
.Y(n_2136)
);

INVx3_ASAP7_75t_SL g2137 ( 
.A(n_2107),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2122),
.Y(n_2138)
);

INVx1_ASAP7_75t_SL g2139 ( 
.A(n_2123),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2095),
.B(n_2104),
.Y(n_2140)
);

OA21x2_ASAP7_75t_L g2141 ( 
.A1(n_2109),
.A2(n_2068),
.B(n_2060),
.Y(n_2141)
);

AND2x4_ASAP7_75t_L g2142 ( 
.A(n_2083),
.B(n_2059),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2102),
.B(n_2054),
.Y(n_2143)
);

INVx3_ASAP7_75t_L g2144 ( 
.A(n_2098),
.Y(n_2144)
);

AOI22xp5_ASAP7_75t_L g2145 ( 
.A1(n_2113),
.A2(n_2056),
.B1(n_2068),
.B2(n_2060),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2111),
.B(n_2054),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2118),
.B(n_2121),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2124),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2106),
.A2(n_2068),
.B1(n_2060),
.B2(n_2073),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2086),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2094),
.B(n_2046),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2117),
.B(n_2082),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_2083),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2118),
.B(n_2121),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2124),
.Y(n_2155)
);

AOI21xp33_ASAP7_75t_L g2156 ( 
.A1(n_2129),
.A2(n_2084),
.B(n_2108),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_2131),
.B(n_2085),
.Y(n_2157)
);

O2A1O1Ixp33_ASAP7_75t_L g2158 ( 
.A1(n_2129),
.A2(n_2108),
.B(n_2098),
.C(n_2082),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2142),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2131),
.B(n_2092),
.Y(n_2160)
);

OAI211xp5_ASAP7_75t_L g2161 ( 
.A1(n_2140),
.A2(n_2153),
.B(n_2139),
.C(n_2136),
.Y(n_2161)
);

OR2x2_ASAP7_75t_L g2162 ( 
.A(n_2143),
.B(n_2084),
.Y(n_2162)
);

OAI211xp5_ASAP7_75t_L g2163 ( 
.A1(n_2153),
.A2(n_2099),
.B(n_2119),
.C(n_2113),
.Y(n_2163)
);

OAI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_2151),
.A2(n_2119),
.B1(n_2046),
.B2(n_2115),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2147),
.B(n_2085),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2135),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2130),
.Y(n_2167)
);

AOI22xp33_ASAP7_75t_L g2168 ( 
.A1(n_2133),
.A2(n_2076),
.B1(n_2073),
.B2(n_2086),
.Y(n_2168)
);

NAND2x1p5_ASAP7_75t_L g2169 ( 
.A(n_2144),
.B(n_2099),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2130),
.Y(n_2170)
);

OAI322xp33_ASAP7_75t_L g2171 ( 
.A1(n_2145),
.A2(n_2116),
.A3(n_2092),
.B1(n_2100),
.B2(n_2097),
.C1(n_2120),
.C2(n_2107),
.Y(n_2171)
);

AOI22xp5_ASAP7_75t_L g2172 ( 
.A1(n_2145),
.A2(n_2076),
.B1(n_2073),
.B2(n_2012),
.Y(n_2172)
);

AOI21xp33_ASAP7_75t_SL g2173 ( 
.A1(n_2137),
.A2(n_2100),
.B(n_2097),
.Y(n_2173)
);

AOI22xp5_ASAP7_75t_L g2174 ( 
.A1(n_2134),
.A2(n_2076),
.B1(n_2073),
.B2(n_2012),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_2152),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_SL g2176 ( 
.A(n_2142),
.B(n_2029),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2130),
.Y(n_2177)
);

NAND3xp33_ASAP7_75t_SL g2178 ( 
.A(n_2136),
.B(n_2033),
.C(n_2046),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_2142),
.A2(n_2074),
.B(n_2033),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_2158),
.B(n_2144),
.Y(n_2180)
);

OAI21xp33_ASAP7_75t_L g2181 ( 
.A1(n_2156),
.A2(n_2154),
.B(n_2147),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2157),
.B(n_2137),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2165),
.B(n_2137),
.Y(n_2183)
);

CKINVDCx16_ASAP7_75t_R g2184 ( 
.A(n_2160),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2175),
.B(n_2128),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_2167),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_2162),
.B(n_2128),
.Y(n_2187)
);

NAND2xp5_ASAP7_75t_SL g2188 ( 
.A(n_2158),
.B(n_2142),
.Y(n_2188)
);

HB1xp67_ASAP7_75t_L g2189 ( 
.A(n_2170),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2177),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2159),
.B(n_2154),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2166),
.B(n_2178),
.Y(n_2192)
);

NOR2x1_ASAP7_75t_L g2193 ( 
.A(n_2161),
.B(n_2144),
.Y(n_2193)
);

AND2x2_ASAP7_75t_L g2194 ( 
.A(n_2176),
.B(n_2146),
.Y(n_2194)
);

OAI211xp5_ASAP7_75t_L g2195 ( 
.A1(n_2193),
.A2(n_2161),
.B(n_2163),
.C(n_2173),
.Y(n_2195)
);

NAND3xp33_ASAP7_75t_SL g2196 ( 
.A(n_2188),
.B(n_2163),
.C(n_2139),
.Y(n_2196)
);

NOR3xp33_ASAP7_75t_L g2197 ( 
.A(n_2184),
.B(n_2171),
.C(n_2164),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2191),
.B(n_2146),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2192),
.A2(n_2174),
.B1(n_2144),
.B2(n_2168),
.Y(n_2199)
);

AOI221xp5_ASAP7_75t_L g2200 ( 
.A1(n_2180),
.A2(n_2149),
.B1(n_2172),
.B2(n_2179),
.C(n_2155),
.Y(n_2200)
);

OAI21xp5_ASAP7_75t_SL g2201 ( 
.A1(n_2180),
.A2(n_2169),
.B(n_2096),
.Y(n_2201)
);

AOI21x1_ASAP7_75t_L g2202 ( 
.A1(n_2189),
.A2(n_2127),
.B(n_2126),
.Y(n_2202)
);

AOI322xp5_ASAP7_75t_L g2203 ( 
.A1(n_2189),
.A2(n_2076),
.A3(n_2150),
.B1(n_2155),
.B2(n_2127),
.C1(n_2126),
.C2(n_2132),
.Y(n_2203)
);

AOI21xp5_ASAP7_75t_L g2204 ( 
.A1(n_2187),
.A2(n_2169),
.B(n_2138),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2185),
.B(n_2101),
.Y(n_2205)
);

OAI21xp5_ASAP7_75t_L g2206 ( 
.A1(n_2181),
.A2(n_2138),
.B(n_2132),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2202),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2198),
.Y(n_2208)
);

AO21x1_ASAP7_75t_L g2209 ( 
.A1(n_2197),
.A2(n_2190),
.B(n_2186),
.Y(n_2209)
);

XNOR2xp5_ASAP7_75t_L g2210 ( 
.A(n_2196),
.B(n_2194),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2195),
.A2(n_2182),
.B1(n_2183),
.B2(n_2120),
.Y(n_2211)
);

OAI22xp5_ASAP7_75t_L g2212 ( 
.A1(n_2200),
.A2(n_2199),
.B1(n_2201),
.B2(n_2205),
.Y(n_2212)
);

AOI211xp5_ASAP7_75t_L g2213 ( 
.A1(n_2206),
.A2(n_2204),
.B(n_2148),
.C(n_2203),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2207),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_2210),
.B(n_2087),
.Y(n_2215)
);

NOR2xp33_ASAP7_75t_L g2216 ( 
.A(n_2211),
.B(n_2148),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2209),
.B(n_2074),
.Y(n_2217)
);

NOR2x1_ASAP7_75t_L g2218 ( 
.A(n_2208),
.B(n_2051),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2213),
.Y(n_2219)
);

HB1xp67_ASAP7_75t_L g2220 ( 
.A(n_2212),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2210),
.Y(n_2221)
);

INVx1_ASAP7_75t_SL g2222 ( 
.A(n_2215),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2217),
.A2(n_2141),
.B(n_2150),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2217),
.Y(n_2224)
);

NOR2xp33_ASAP7_75t_R g2225 ( 
.A(n_2221),
.B(n_2039),
.Y(n_2225)
);

OAI211xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2219),
.A2(n_2150),
.B(n_2116),
.C(n_2091),
.Y(n_2226)
);

NOR2x1_ASAP7_75t_SL g2227 ( 
.A(n_2214),
.B(n_2051),
.Y(n_2227)
);

NAND2xp33_ASAP7_75t_R g2228 ( 
.A(n_2216),
.B(n_2141),
.Y(n_2228)
);

OAI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_2222),
.A2(n_2220),
.B1(n_2218),
.B2(n_2063),
.Y(n_2229)
);

NAND3xp33_ASAP7_75t_L g2230 ( 
.A(n_2224),
.B(n_2141),
.C(n_2063),
.Y(n_2230)
);

NOR2x1_ASAP7_75t_L g2231 ( 
.A(n_2223),
.B(n_2039),
.Y(n_2231)
);

NAND3x1_ASAP7_75t_L g2232 ( 
.A(n_2225),
.B(n_2096),
.C(n_2093),
.Y(n_2232)
);

OR2x2_ASAP7_75t_L g2233 ( 
.A(n_2228),
.B(n_2093),
.Y(n_2233)
);

NOR3xp33_ASAP7_75t_L g2234 ( 
.A(n_2229),
.B(n_2226),
.C(n_2227),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2233),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_2230),
.Y(n_2236)
);

OAI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2235),
.A2(n_2231),
.B1(n_2232),
.B2(n_2141),
.Y(n_2237)
);

AOI322xp5_ASAP7_75t_L g2238 ( 
.A1(n_2234),
.A2(n_2236),
.A3(n_2089),
.B1(n_2091),
.B2(n_2103),
.C1(n_2090),
.C2(n_2087),
.Y(n_2238)
);

OAI21x1_ASAP7_75t_L g2239 ( 
.A1(n_2237),
.A2(n_2103),
.B(n_2090),
.Y(n_2239)
);

AND2x2_ASAP7_75t_SL g2240 ( 
.A(n_2238),
.B(n_2089),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2237),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2240),
.B(n_2239),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2241),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_2241),
.Y(n_2244)
);

OR2x2_ASAP7_75t_L g2245 ( 
.A(n_2244),
.B(n_2080),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2245),
.Y(n_2246)
);

BUFx2_ASAP7_75t_L g2247 ( 
.A(n_2246),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2247),
.A2(n_2243),
.B1(n_2244),
.B2(n_2242),
.Y(n_2248)
);

AOI322xp5_ASAP7_75t_L g2249 ( 
.A1(n_2248),
.A2(n_2081),
.A3(n_2079),
.B1(n_2067),
.B2(n_2069),
.C1(n_2075),
.C2(n_2066),
.Y(n_2249)
);

OAI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_2249),
.A2(n_2080),
.B1(n_2081),
.B2(n_2079),
.Y(n_2250)
);

AOI211xp5_ASAP7_75t_L g2251 ( 
.A1(n_2250),
.A2(n_2037),
.B(n_1996),
.C(n_2069),
.Y(n_2251)
);


endmodule