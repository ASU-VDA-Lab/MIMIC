module real_aes_2115_n_10 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_1, n_10);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_1;
output n_10;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_13;
wire n_34;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_35;
wire n_15;
wire n_27;
wire n_23;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
CKINVDCx16_ASAP7_75t_R g24 ( .A(n_0), .Y(n_24) );
INVx1_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
BUFx2_ASAP7_75t_L g25 ( .A(n_2), .Y(n_25) );
NAND2xp5_ASAP7_75t_SL g28 ( .A(n_3), .B(n_29), .Y(n_28) );
AOI222xp33_ASAP7_75t_L g10 ( .A1(n_4), .A2(n_6), .B1(n_11), .B2(n_26), .C1(n_27), .C2(n_33), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_5), .B(n_24), .Y(n_23) );
INVx1_ASAP7_75t_L g15 ( .A(n_7), .Y(n_15) );
OR2x6_ASAP7_75t_L g13 ( .A(n_8), .B(n_14), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g20 ( .A(n_9), .Y(n_20) );
INVx1_ASAP7_75t_SL g11 ( .A(n_12), .Y(n_11) );
NAND2xp5_ASAP7_75t_SL g12 ( .A(n_13), .B(n_17), .Y(n_12) );
OR2x2_ASAP7_75t_L g19 ( .A(n_13), .B(n_20), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g32 ( .A(n_13), .Y(n_32) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_15), .B(n_16), .Y(n_14) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_17), .Y(n_26) );
CKINVDCx16_ASAP7_75t_R g35 ( .A(n_17), .Y(n_35) );
NOR2x1_ASAP7_75t_L g17 ( .A(n_18), .B(n_21), .Y(n_17) );
INVx3_ASAP7_75t_L g18 ( .A(n_19), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_20), .B(n_32), .Y(n_31) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_22), .B(n_25), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_23), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_28), .Y(n_27) );
INVx1_ASAP7_75t_SL g29 ( .A(n_30), .Y(n_29) );
BUFx2_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx1_ASAP7_75t_L g33 ( .A(n_34), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_35), .Y(n_34) );
endmodule