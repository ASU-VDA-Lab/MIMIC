module fake_jpeg_29706_n_406 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_406);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_406;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_45),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx6p67_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_49),
.Y(n_116)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_56),
.A2(n_21),
.B1(n_40),
.B2(n_34),
.Y(n_96)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_62),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_43),
.B(n_6),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_28),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_72),
.Y(n_111)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_70),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_71),
.B(n_73),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_82),
.Y(n_125)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_75),
.B(n_76),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_78),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_79),
.B(n_80),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_81),
.B(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_20),
.B(n_6),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_84),
.B(n_85),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_32),
.B(n_7),
.C(n_12),
.Y(n_85)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_36),
.B1(n_23),
.B2(n_38),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_87),
.A2(n_98),
.B1(n_122),
.B2(n_22),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_71),
.A2(n_36),
.B1(n_17),
.B2(n_23),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_88),
.A2(n_91),
.B1(n_107),
.B2(n_117),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_36),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_89),
.B(n_93),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_28),
.B1(n_40),
.B2(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_41),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_22),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_41),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_97),
.B(n_99),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_46),
.A2(n_15),
.B1(n_37),
.B2(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_41),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_15),
.B1(n_37),
.B2(n_29),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_54),
.A2(n_34),
.B1(n_17),
.B2(n_15),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_134),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_37),
.B1(n_29),
.B2(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_133),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_69),
.A2(n_30),
.B1(n_24),
.B2(n_18),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_30),
.B1(n_24),
.B2(n_18),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_76),
.B1(n_72),
.B2(n_80),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_41),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_52),
.B(n_41),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_65),
.B(n_24),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_7),
.C(n_12),
.Y(n_166)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_65),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_151),
.Y(n_188)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_78),
.B1(n_77),
.B2(n_18),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_140),
.A2(n_144),
.B1(n_156),
.B2(n_104),
.Y(n_205)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_102),
.A2(n_78),
.B1(n_77),
.B2(n_49),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_145),
.Y(n_192)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_100),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_150),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_94),
.B(n_76),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_154),
.B1(n_103),
.B2(n_104),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_72),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_162),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_105),
.A2(n_45),
.B1(n_50),
.B2(n_22),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_155),
.A2(n_167),
.B1(n_176),
.B2(n_129),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_108),
.A2(n_115),
.B1(n_126),
.B2(n_110),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_175),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_100),
.Y(n_159)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_159),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_100),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_129),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_161),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_88),
.B(n_22),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_7),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_170),
.Y(n_221)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2x1p5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_0),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_103),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_105),
.A2(n_5),
.B1(n_11),
.B2(n_10),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_168),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_134),
.B(n_4),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_93),
.A2(n_4),
.B(n_9),
.C(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_173),
.B(n_174),
.Y(n_198)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

INVx11_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_124),
.A2(n_9),
.B1(n_14),
.B2(n_2),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_114),
.B(n_9),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_177),
.B(n_182),
.Y(n_223)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_179),
.B(n_180),
.Y(n_212)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_113),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_181),
.B(n_131),
.Y(n_196)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_138),
.B(n_130),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_200),
.Y(n_232)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_128),
.C(n_99),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_222),
.C(n_172),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_128),
.B(n_132),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_204),
.B(n_215),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_103),
.B(n_127),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_191),
.A2(n_165),
.B(n_159),
.Y(n_236)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_165),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_151),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_205),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_131),
.B1(n_119),
.B2(n_115),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_203),
.A2(n_206),
.B1(n_220),
.B2(n_159),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_137),
.A2(n_121),
.B(n_97),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_147),
.A2(n_124),
.B1(n_120),
.B2(n_101),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_153),
.B(n_101),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_160),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_218),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_112),
.B1(n_90),
.B2(n_2),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_182),
.B1(n_163),
.B2(n_168),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_90),
.B(n_112),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_148),
.A2(n_9),
.B(n_1),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_147),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_0),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_224),
.A2(n_247),
.B1(n_255),
.B2(n_206),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_228),
.B1(n_239),
.B2(n_205),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_220),
.A2(n_171),
.B1(n_178),
.B2(n_169),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_222),
.B(n_170),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_229),
.B(n_230),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_231),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_197),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_236),
.C(n_199),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_136),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_248),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_186),
.B(n_180),
.C(n_179),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_244),
.C(n_212),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_198),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_241),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_152),
.B1(n_174),
.B2(n_173),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_240),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_187),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_256),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_139),
.C(n_143),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_246),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_181),
.B1(n_145),
.B2(n_142),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_149),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_207),
.A2(n_157),
.B(n_146),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_249),
.A2(n_199),
.B(n_190),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_145),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_209),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_184),
.A2(n_161),
.B(n_142),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_252),
.A2(n_189),
.B(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_209),
.Y(n_253)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_253),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_1),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_187),
.A2(n_194),
.B1(n_219),
.B2(n_214),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_223),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_223),
.B(n_1),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_2),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_260),
.B(n_263),
.C(n_272),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_261),
.B(n_227),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_274),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_215),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_187),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_245),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_245),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_269),
.A2(n_279),
.B(n_286),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_188),
.C(n_199),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_188),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_275),
.A2(n_290),
.B1(n_226),
.B2(n_225),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_276),
.B(n_230),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_211),
.B(n_201),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_225),
.A2(n_203),
.B1(n_221),
.B2(n_216),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_224),
.B1(n_249),
.B2(n_250),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_244),
.B(n_221),
.C(n_195),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_233),
.C(n_229),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_232),
.B(n_195),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_287),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_210),
.B(n_202),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_232),
.B(n_210),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_256),
.B(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_289),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_235),
.B(n_213),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_255),
.A2(n_175),
.B1(n_192),
.B2(n_183),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_273),
.Y(n_296)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_296),
.Y(n_321)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_297),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_227),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_298),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_299),
.A2(n_312),
.B1(n_315),
.B2(n_269),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_301),
.B(n_316),
.C(n_260),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_263),
.B(n_236),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_299),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_281),
.Y(n_305)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_307),
.A2(n_264),
.B(n_286),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_259),
.B(n_228),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_278),
.Y(n_309)
);

OAI21xp33_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_314),
.B(n_287),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_261),
.B(n_258),
.Y(n_310)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_310),
.B(n_311),
.C(n_266),
.Y(n_327)
);

AOI21xp33_ASAP7_75t_L g311 ( 
.A1(n_268),
.A2(n_257),
.B(n_245),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_267),
.C(n_268),
.Y(n_337)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_279),
.A2(n_245),
.B1(n_225),
.B2(n_239),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_317),
.B(n_320),
.C(n_322),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_327),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_260),
.C(n_263),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_276),
.C(n_265),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_276),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_324),
.C(n_326),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_283),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_301),
.B(n_313),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_329),
.A2(n_307),
.B(n_270),
.Y(n_351)
);

AOI322xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_293),
.A3(n_274),
.B1(n_303),
.B2(n_292),
.C1(n_271),
.C2(n_259),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_304),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_329),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_283),
.C(n_272),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_334),
.C(n_337),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_267),
.C(n_264),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_335),
.B(n_320),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_303),
.B1(n_315),
.B2(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_340),
.A2(n_346),
.B1(n_348),
.B2(n_355),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_271),
.B(n_300),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_341),
.A2(n_350),
.B(n_351),
.Y(n_365)
);

AOI21x1_ASAP7_75t_L g342 ( 
.A1(n_338),
.A2(n_300),
.B(n_289),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_334),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_336),
.B(n_266),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_353),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_345),
.B(n_254),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_319),
.A2(n_275),
.B1(n_292),
.B2(n_290),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_347),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_335),
.A2(n_270),
.B1(n_262),
.B2(n_314),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_328),
.A2(n_307),
.B(n_330),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_304),
.C(n_288),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_354),
.B(n_356),
.C(n_333),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_330),
.A2(n_309),
.B1(n_306),
.B2(n_296),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_282),
.C(n_285),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_364),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_339),
.A2(n_324),
.B1(n_323),
.B2(n_321),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_363),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_360),
.B(n_345),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_322),
.C(n_337),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_370),
.C(n_344),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_354),
.B(n_328),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_285),
.Y(n_367)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_325),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_369),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_246),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_281),
.C(n_253),
.Y(n_370)
);

AOI31xp67_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_351),
.A3(n_340),
.B(n_352),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_371),
.B(n_375),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_370),
.Y(n_383)
);

NAND4xp25_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_344),
.C(n_247),
.D(n_356),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_377),
.Y(n_384)
);

OR2x2_ASAP7_75t_L g375 ( 
.A(n_367),
.B(n_346),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_366),
.A2(n_297),
.B1(n_277),
.B2(n_240),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_378),
.A2(n_240),
.B1(n_366),
.B2(n_192),
.Y(n_382)
);

AO21x1_ASAP7_75t_L g380 ( 
.A1(n_365),
.A2(n_251),
.B(n_231),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_380),
.A2(n_357),
.B(n_362),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_382),
.B(n_383),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_378),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_387),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_375),
.B(n_365),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_386),
.B(n_381),
.Y(n_392)
);

OR2x6_ASAP7_75t_SL g388 ( 
.A(n_380),
.B(n_364),
.Y(n_388)
);

AOI21x1_ASAP7_75t_L g394 ( 
.A1(n_388),
.A2(n_372),
.B(n_213),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_376),
.B(n_361),
.Y(n_390)
);

NOR4xp25_ASAP7_75t_L g393 ( 
.A(n_390),
.B(n_360),
.C(n_372),
.D(n_183),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_384),
.A2(n_373),
.B(n_379),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_391),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_392),
.B(n_395),
.C(n_389),
.Y(n_398)
);

NOR2x1_ASAP7_75t_L g401 ( 
.A(n_393),
.B(n_394),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_SL g395 ( 
.A(n_388),
.B(n_3),
.C(n_389),
.Y(n_395)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_398),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_385),
.C(n_388),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_399),
.A2(n_3),
.B1(n_397),
.B2(n_400),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_397),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_404),
.B(n_405),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_402),
.B(n_401),
.Y(n_405)
);


endmodule