module fake_jpeg_5972_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_219;
wire n_70;
wire n_102;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_0),
.B(n_14),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_SL g99 ( 
.A(n_45),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_2),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_53),
.Y(n_95)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_21),
.B(n_2),
.Y(n_53)
);

INVxp67_ASAP7_75t_SL g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_57),
.B1(n_34),
.B2(n_37),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_4),
.Y(n_56)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_38),
.Y(n_86)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_4),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_4),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_20),
.C(n_31),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_25),
.B1(n_32),
.B2(n_22),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_62),
.A2(n_85),
.B1(n_17),
.B2(n_19),
.Y(n_112)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_29),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_72),
.B(n_78),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_84),
.Y(n_120)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_59),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_57),
.B1(n_55),
.B2(n_22),
.Y(n_85)
);

OR2x4_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_27),
.Y(n_116)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

CKINVDCx12_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_89),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_34),
.B1(n_39),
.B2(n_37),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_35),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_104),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_35),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_105),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_31),
.C(n_20),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_114),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_63),
.B1(n_82),
.B2(n_81),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_77),
.A2(n_25),
.B1(n_41),
.B2(n_36),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_113),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_18),
.C(n_36),
.Y(n_114)
);

OA22x2_ASAP7_75t_L g115 ( 
.A1(n_90),
.A2(n_52),
.B1(n_35),
.B2(n_27),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_115),
.A2(n_124),
.B1(n_8),
.B2(n_9),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_126),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_19),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_121),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_27),
.B(n_26),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_98),
.A2(n_52),
.B1(n_13),
.B2(n_12),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_94),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_125),
.A2(n_132),
.B1(n_5),
.B2(n_7),
.Y(n_134)
);

AND2x2_ASAP7_75t_SL g126 ( 
.A(n_100),
.B(n_5),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_64),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_119),
.B1(n_126),
.B2(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_76),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_133),
.B(n_134),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_125),
.A2(n_63),
.B1(n_97),
.B2(n_81),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_146),
.B1(n_147),
.B2(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_139),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_69),
.Y(n_141)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_141),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_100),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_143),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_74),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_69),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_110),
.B(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_103),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_153),
.B(n_160),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_116),
.A2(n_70),
.B1(n_82),
.B2(n_91),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_161),
.Y(n_168)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_111),
.Y(n_159)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_93),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_165),
.Y(n_193)
);

CKINVDCx11_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_163),
.B(n_169),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_143),
.C(n_136),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_154),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_173),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_120),
.C(n_121),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_182),
.C(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_107),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_128),
.B1(n_106),
.B2(n_117),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_180),
.B1(n_105),
.B2(n_93),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_178),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_145),
.A2(n_107),
.B(n_128),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_139),
.B(n_151),
.Y(n_198)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_156),
.A2(n_106),
.B1(n_124),
.B2(n_70),
.Y(n_180)
);

MAJx2_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_118),
.C(n_99),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_184),
.B(n_91),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_152),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_189),
.C(n_192),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_172),
.A2(n_158),
.B1(n_145),
.B2(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_195),
.B1(n_198),
.B2(n_205),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_196),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_135),
.C(n_140),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_157),
.B1(n_134),
.B2(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_185),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_197),
.B(n_201),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_199),
.B(n_202),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_181),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_164),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_171),
.B(n_118),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_207),
.B(n_210),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_203),
.A2(n_169),
.B1(n_183),
.B2(n_166),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_206),
.C(n_198),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_175),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_214),
.B(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_162),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_187),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_221),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_164),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_222),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_201),
.B1(n_191),
.B2(n_176),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_195),
.Y(n_236)
);

XOR2x2_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_189),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_207),
.B1(n_220),
.B2(n_221),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_208),
.A2(n_192),
.B1(n_193),
.B2(n_188),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_232),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_220),
.C(n_210),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_219),
.A2(n_177),
.B1(n_166),
.B2(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_209),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_226),
.A2(n_217),
.B(n_219),
.C(n_211),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_235),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_239),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_228),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_237),
.A2(n_229),
.B(n_182),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_240),
.A2(n_241),
.B(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_177),
.B1(n_179),
.B2(n_234),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_249),
.C(n_237),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_234),
.B1(n_178),
.B2(n_224),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_231),
.B1(n_205),
.B2(n_218),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_239),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_254),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_248),
.B(n_179),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_255),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_230),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

AOI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_257),
.A2(n_258),
.B(n_212),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_252),
.A2(n_246),
.B(n_247),
.C(n_245),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_256),
.B(n_9),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_259),
.B(n_105),
.C(n_10),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_261),
.A2(n_102),
.B(n_122),
.Y(n_263)
);

XNOR2x2_ASAP7_75t_SL g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_102),
.Y(n_265)
);


endmodule