module real_aes_18055_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_502;
wire n_505;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_0), .Y(n_195) );
AND2x4_ASAP7_75t_L g114 ( .A(n_1), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_2), .A2(n_4), .B1(n_219), .B2(n_592), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_3), .A2(n_19), .B1(n_146), .B2(n_187), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_5), .A2(n_50), .B1(n_193), .B2(n_507), .Y(n_506) );
BUFx3_ASAP7_75t_L g261 ( .A(n_6), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_7), .A2(n_13), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_9), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_10), .B(n_237), .Y(n_236) );
BUFx2_ASAP7_75t_L g106 ( .A(n_11), .Y(n_106) );
OR2x2_ASAP7_75t_L g122 ( .A(n_11), .B(n_29), .Y(n_122) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_12), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_14), .B(n_150), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_15), .B(n_176), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_16), .A2(n_83), .B1(n_146), .B2(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_17), .A2(n_125), .B1(n_126), .B2(n_127), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_17), .Y(n_125) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_18), .A2(n_45), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_20), .B(n_187), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_21), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_22), .B(n_144), .Y(n_542) );
INVx4_ASAP7_75t_R g531 ( .A(n_23), .Y(n_531) );
AO32x1_ASAP7_75t_L g137 ( .A1(n_24), .A2(n_138), .A3(n_141), .B1(n_152), .B2(n_156), .Y(n_137) );
AO32x2_ASAP7_75t_L g269 ( .A1(n_24), .A2(n_138), .A3(n_141), .B1(n_152), .B2(n_156), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_25), .B(n_187), .Y(n_548) );
INVx1_ASAP7_75t_L g594 ( .A(n_26), .Y(n_594) );
A2O1A1Ixp33_ASAP7_75t_SL g574 ( .A1(n_27), .A2(n_151), .B(n_515), .C(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_28), .A2(n_42), .B1(n_148), .B2(n_515), .Y(n_582) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_30), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_31), .A2(n_48), .B1(n_187), .B2(n_188), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g145 ( .A1(n_32), .A2(n_88), .B1(n_146), .B2(n_148), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_33), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_34), .B(n_164), .Y(n_171) );
INVx1_ASAP7_75t_L g545 ( .A(n_35), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_36), .A2(n_65), .B1(n_148), .B2(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_37), .B(n_515), .Y(n_547) );
CKINVDCx5p33_ASAP7_75t_R g557 ( .A(n_38), .Y(n_557) );
INVx2_ASAP7_75t_L g813 ( .A(n_39), .Y(n_813) );
INVx1_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
BUFx3_ASAP7_75t_L g816 ( .A(n_40), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_41), .B(n_173), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_43), .A2(n_84), .B1(n_148), .B2(n_515), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g532 ( .A(n_44), .Y(n_532) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_46), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_47), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_49), .A2(n_77), .B1(n_164), .B2(n_196), .Y(n_247) );
CKINVDCx5p33_ASAP7_75t_R g521 ( .A(n_51), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_52), .A2(n_81), .B1(n_146), .B2(n_150), .Y(n_257) );
INVx1_ASAP7_75t_L g140 ( .A(n_53), .Y(n_140) );
AND2x4_ASAP7_75t_L g154 ( .A(n_54), .B(n_155), .Y(n_154) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_55), .A2(n_493), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_55), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_56), .A2(n_100), .B1(n_116), .B2(n_839), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_57), .A2(n_89), .B1(n_148), .B2(n_590), .Y(n_589) );
AO22x1_ASAP7_75t_L g502 ( .A1(n_58), .A2(n_71), .B1(n_503), .B2(n_504), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_59), .B(n_146), .Y(n_235) );
INVx1_ASAP7_75t_L g155 ( .A(n_60), .Y(n_155) );
AND2x2_ASAP7_75t_L g577 ( .A(n_61), .B(n_156), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_62), .B(n_156), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_63), .A2(n_168), .B(n_193), .C(n_194), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_64), .B(n_146), .C(n_240), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_66), .B(n_193), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_67), .Y(n_571) );
INVx1_ASAP7_75t_L g118 ( .A(n_68), .Y(n_118) );
AND2x2_ASAP7_75t_L g198 ( .A(n_69), .B(n_199), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_70), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g817 ( .A1(n_72), .A2(n_818), .B1(n_829), .B2(n_832), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_73), .B(n_187), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_74), .A2(n_93), .B1(n_150), .B2(n_196), .Y(n_249) );
INVx2_ASAP7_75t_L g144 ( .A(n_75), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_76), .B(n_224), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_78), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_79), .B(n_156), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_80), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_82), .B(n_178), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_85), .B(n_240), .Y(n_239) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_86), .A2(n_98), .B1(n_148), .B2(n_188), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_87), .B(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_90), .B(n_156), .Y(n_554) );
INVx1_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_91), .B(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_92), .B(n_176), .Y(n_175) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_94), .A2(n_191), .B(n_193), .C(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g534 ( .A(n_95), .B(n_199), .Y(n_534) );
NAND2xp33_ASAP7_75t_L g560 ( .A(n_96), .B(n_237), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g218 ( .A(n_97), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx8_ASAP7_75t_L g840 ( .A(n_101), .Y(n_840) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_107), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
NOR2x1p5_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
AND3x2_ASAP7_75t_L g120 ( .A(n_108), .B(n_112), .C(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g827 ( .A(n_109), .Y(n_827) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_114), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g490 ( .A(n_113), .Y(n_490) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_123), .Y(n_116) );
INVx1_ASAP7_75t_L g828 ( .A(n_117), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_121), .B(n_815), .Y(n_814) );
AND2x6_ASAP7_75t_SL g825 ( .A(n_121), .B(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_122), .B(n_816), .Y(n_838) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_809), .B(n_817), .Y(n_123) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AO22x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_488), .B1(n_491), .B2(n_493), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_375), .Y(n_128) );
AND4x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_284), .C(n_322), .D(n_360), .Y(n_129) );
NOR2x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_262), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_201), .B(n_212), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_157), .Y(n_133) );
NAND2xp5_ASAP7_75t_R g333 ( .A(n_134), .B(n_281), .Y(n_333) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g434 ( .A(n_136), .B(n_312), .Y(n_434) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OR2x2_ASAP7_75t_L g203 ( .A(n_137), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g295 ( .A(n_137), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_137), .B(n_204), .Y(n_309) );
INVx4_ASAP7_75t_L g156 ( .A(n_138), .Y(n_156) );
INVx2_ASAP7_75t_SL g160 ( .A(n_138), .Y(n_160) );
BUFx3_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_138), .B(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_138), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g549 ( .A(n_138), .B(n_228), .Y(n_549) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_145), .B1(n_149), .B2(n_151), .Y(n_141) );
O2A1O1Ixp5_ASAP7_75t_L g217 ( .A1(n_142), .A2(n_218), .B(n_219), .C(n_221), .Y(n_217) );
OAI21xp5_ASAP7_75t_L g569 ( .A1(n_142), .A2(n_570), .B(n_572), .Y(n_569) );
BUFx4f_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g240 ( .A(n_143), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_143), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx8_ASAP7_75t_L g151 ( .A(n_144), .Y(n_151) );
INVx2_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx1_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
INVx2_ASAP7_75t_SL g164 ( .A(n_146), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_146), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_147), .Y(n_148) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_147), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g193 ( .A(n_147), .Y(n_193) );
INVx1_ASAP7_75t_L g196 ( .A(n_147), .Y(n_196) );
INVx1_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_147), .Y(n_237) );
INVx1_ASAP7_75t_L g508 ( .A(n_147), .Y(n_508) );
INVx3_ASAP7_75t_L g515 ( .A(n_147), .Y(n_515) );
INVx2_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_148), .B(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g592 ( .A(n_148), .Y(n_592) );
INVx3_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
INVxp67_ASAP7_75t_SL g503 ( .A(n_150), .Y(n_503) );
INVx6_ASAP7_75t_L g174 ( .A(n_151), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_151), .A2(n_235), .B(n_236), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_151), .A2(n_174), .B1(n_257), .B2(n_258), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_151), .A2(n_502), .B(n_505), .C(n_510), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_151), .A2(n_560), .B(n_561), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_151), .B(n_502), .Y(n_606) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_152), .A2(n_162), .B(n_170), .Y(n_161) );
INVx2_ASAP7_75t_SL g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_SL g250 ( .A(n_153), .Y(n_250) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g197 ( .A(n_154), .Y(n_197) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_154), .A2(n_205), .A3(n_206), .B(n_210), .Y(n_204) );
BUFx10_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
BUFx10_ASAP7_75t_L g519 ( .A(n_154), .Y(n_519) );
INVx2_ASAP7_75t_L g255 ( .A(n_156), .Y(n_255) );
NOR2x1_ASAP7_75t_L g562 ( .A(n_156), .B(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_179), .Y(n_157) );
BUFx2_ASAP7_75t_L g202 ( .A(n_158), .Y(n_202) );
AND2x2_ASAP7_75t_L g267 ( .A(n_158), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g282 ( .A(n_158), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_158), .B(n_204), .Y(n_299) );
INVx3_ASAP7_75t_L g312 ( .A(n_158), .Y(n_312) );
AND2x2_ASAP7_75t_L g347 ( .A(n_158), .B(n_269), .Y(n_347) );
INVx2_ASAP7_75t_L g359 ( .A(n_158), .Y(n_359) );
INVx1_ASAP7_75t_L g363 ( .A(n_158), .Y(n_363) );
INVxp67_ASAP7_75t_L g400 ( .A(n_158), .Y(n_400) );
OR2x2_ASAP7_75t_L g413 ( .A(n_158), .B(n_296), .Y(n_413) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
OAI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_161), .B(n_175), .Y(n_159) );
AOI21x1_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_167), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_166), .A2(n_239), .B(n_241), .Y(n_238) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_167), .A2(n_174), .B1(n_207), .B2(n_209), .Y(n_206) );
OAI21x1_ASAP7_75t_L g505 ( .A1(n_167), .A2(n_506), .B(n_509), .Y(n_505) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_167), .A2(n_547), .B(n_548), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_167), .A2(n_174), .B1(n_581), .B2(n_582), .Y(n_580) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g225 ( .A(n_169), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_174), .Y(n_170) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_174), .A2(n_247), .B1(n_248), .B2(n_249), .Y(n_246) );
OAI22x1_ASAP7_75t_L g513 ( .A1(n_174), .A2(n_514), .B1(n_517), .B2(n_518), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_174), .A2(n_518), .B1(n_589), .B2(n_591), .Y(n_588) );
INVx2_ASAP7_75t_L g182 ( .A(n_176), .Y(n_182) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g200 ( .A(n_178), .Y(n_200) );
INVx2_ASAP7_75t_L g232 ( .A(n_178), .Y(n_232) );
OAI21xp33_ASAP7_75t_L g510 ( .A1(n_178), .A2(n_197), .B(n_509), .Y(n_510) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx1_ASAP7_75t_L g265 ( .A(n_180), .Y(n_265) );
INVx1_ASAP7_75t_L g352 ( .A(n_180), .Y(n_352) );
AND2x2_ASAP7_75t_L g367 ( .A(n_180), .B(n_204), .Y(n_367) );
INVx1_ASAP7_75t_L g382 ( .A(n_180), .Y(n_382) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g296 ( .A(n_181), .Y(n_296) );
AOI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_198), .Y(n_181) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_182), .A2(n_525), .B(n_534), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_192), .B(n_197), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_185), .B(n_190), .Y(n_184) );
OAI22xp5_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B1(n_188), .B2(n_189), .Y(n_185) );
INVx2_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_187), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g530 ( .A1(n_188), .A2(n_237), .B1(n_531), .B2(n_532), .Y(n_530) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_SL g248 ( .A(n_191), .Y(n_248) );
INVx1_ASAP7_75t_L g518 ( .A(n_191), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
INVx1_ASAP7_75t_L g504 ( .A(n_196), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_197), .A2(n_569), .B(n_574), .Y(n_568) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_200), .B(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_200), .B(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g567 ( .A(n_200), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_200), .B(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_200), .B(n_594), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_201), .A2(n_471), .B1(n_473), .B2(n_475), .Y(n_470) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_202), .B(n_351), .Y(n_428) );
BUFx2_ASAP7_75t_L g442 ( .A(n_202), .Y(n_442) );
AND2x2_ASAP7_75t_L g460 ( .A(n_202), .B(n_316), .Y(n_460) );
INVx2_ASAP7_75t_L g342 ( .A(n_203), .Y(n_342) );
OR2x2_ASAP7_75t_L g358 ( .A(n_203), .B(n_359), .Y(n_358) );
INVx3_ASAP7_75t_L g266 ( .A(n_204), .Y(n_266) );
AND2x2_ASAP7_75t_L g351 ( .A(n_204), .B(n_352), .Y(n_351) );
AO31x2_ASAP7_75t_L g245 ( .A1(n_205), .A2(n_246), .A3(n_250), .B(n_251), .Y(n_245) );
OR2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_243), .Y(n_212) );
OR2x2_ASAP7_75t_L g407 ( .A(n_213), .B(n_364), .Y(n_407) );
OR2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_230), .Y(n_213) );
AND2x2_ASAP7_75t_L g278 ( .A(n_214), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g319 ( .A(n_214), .Y(n_319) );
INVx2_ASAP7_75t_SL g327 ( .A(n_214), .Y(n_327) );
BUFx2_ASAP7_75t_L g339 ( .A(n_214), .Y(n_339) );
OR2x2_ASAP7_75t_L g427 ( .A(n_214), .B(n_245), .Y(n_427) );
OA21x2_ASAP7_75t_L g214 ( .A1(n_215), .A2(n_216), .B(n_229), .Y(n_214) );
OA21x2_ASAP7_75t_L g292 ( .A1(n_215), .A2(n_216), .B(n_229), .Y(n_292) );
OAI21x1_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_222), .B(n_228), .Y(n_216) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_220), .B(n_573), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_225), .B1(n_226), .B2(n_227), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g556 ( .A1(n_224), .A2(n_516), .B(n_557), .C(n_558), .Y(n_556) );
INVx2_ASAP7_75t_SL g224 ( .A(n_225), .Y(n_224) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_228), .A2(n_234), .B(n_238), .Y(n_233) );
AOI31xp67_ASAP7_75t_L g254 ( .A1(n_228), .A2(n_255), .A3(n_256), .B(n_259), .Y(n_254) );
INVx1_ASAP7_75t_L g563 ( .A(n_228), .Y(n_563) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_228), .A2(n_255), .A3(n_580), .B(n_583), .Y(n_579) );
AND2x2_ASAP7_75t_L g271 ( .A(n_230), .B(n_253), .Y(n_271) );
AND2x2_ASAP7_75t_L g307 ( .A(n_230), .B(n_292), .Y(n_307) );
OAI21xp5_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_233), .B(n_242), .Y(n_230) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_231), .A2(n_233), .B(n_242), .Y(n_277) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AO31x2_ASAP7_75t_L g512 ( .A1(n_232), .A2(n_513), .A3(n_519), .B(n_520), .Y(n_512) );
INVx2_ASAP7_75t_L g590 ( .A(n_237), .Y(n_590) );
INVx1_ASAP7_75t_L g345 ( .A(n_243), .Y(n_345) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_244), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g451 ( .A(n_244), .B(n_431), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_244), .B(n_274), .Y(n_475) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_253), .Y(n_244) );
INVx1_ASAP7_75t_L g279 ( .A(n_245), .Y(n_279) );
INVx2_ASAP7_75t_L g289 ( .A(n_245), .Y(n_289) );
AND2x2_ASAP7_75t_L g303 ( .A(n_245), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g318 ( .A(n_245), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_245), .B(n_292), .Y(n_332) );
OR2x2_ASAP7_75t_L g364 ( .A(n_245), .B(n_304), .Y(n_364) );
INVx1_ASAP7_75t_L g448 ( .A(n_245), .Y(n_448) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_250), .A2(n_567), .A3(n_588), .B(n_593), .Y(n_587) );
AND2x2_ASAP7_75t_L g291 ( .A(n_253), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g329 ( .A(n_253), .Y(n_329) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g305 ( .A(n_254), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_261), .Y(n_260) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_270), .B1(n_272), .B2(n_280), .Y(n_262) );
NAND2x1p5_ASAP7_75t_L g263 ( .A(n_264), .B(n_267), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx1_ASAP7_75t_L g409 ( .A(n_265), .Y(n_409) );
INVx1_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
AND2x4_ASAP7_75t_L g316 ( .A(n_266), .B(n_269), .Y(n_316) );
AND2x2_ASAP7_75t_L g425 ( .A(n_266), .B(n_296), .Y(n_425) );
AND2x2_ASAP7_75t_L g477 ( .A(n_267), .B(n_351), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_267), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g331 ( .A(n_271), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g464 ( .A(n_271), .B(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_278), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_274), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g383 ( .A(n_274), .Y(n_383) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g449 ( .A(n_275), .Y(n_449) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g336 ( .A(n_276), .Y(n_336) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g321 ( .A(n_277), .B(n_305), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_278), .B(n_320), .Y(n_436) );
AND2x2_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
INVx1_ASAP7_75t_L g468 ( .A(n_283), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_293), .B1(n_300), .B2(n_308), .C(n_313), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
AND2x2_ASAP7_75t_L g386 ( .A(n_287), .B(n_307), .Y(n_386) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_288), .B(n_307), .Y(n_355) );
OR2x2_ASAP7_75t_L g370 ( .A(n_288), .B(n_321), .Y(n_370) );
INVx2_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g335 ( .A(n_289), .B(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_L g446 ( .A(n_291), .Y(n_446) );
INVx1_ASAP7_75t_L g406 ( .A(n_292), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
AND2x2_ASAP7_75t_L g466 ( .A(n_294), .B(n_467), .Y(n_466) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
AND2x2_ASAP7_75t_L g420 ( .A(n_295), .B(n_382), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_296), .B(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g341 ( .A(n_296), .Y(n_341) );
INVx1_ASAP7_75t_L g393 ( .A(n_296), .Y(n_393) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI21xp33_ASAP7_75t_L g361 ( .A1(n_301), .A2(n_327), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_306), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g356 ( .A(n_303), .B(n_339), .Y(n_356) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_303), .Y(n_396) );
AND2x2_ASAP7_75t_L g480 ( .A(n_303), .B(n_417), .Y(n_480) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g487 ( .A(n_306), .B(n_404), .Y(n_487) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_SL g388 ( .A(n_309), .Y(n_388) );
AND2x2_ASAP7_75t_L g392 ( .A(n_309), .B(n_393), .Y(n_392) );
AND2x2_ASAP7_75t_L g452 ( .A(n_309), .B(n_312), .Y(n_452) );
AND2x2_ASAP7_75t_L g474 ( .A(n_309), .B(n_399), .Y(n_474) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g371 ( .A(n_312), .B(n_316), .Y(n_371) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g365 ( .A(n_316), .B(n_341), .Y(n_365) );
AND2x2_ASAP7_75t_L g398 ( .A(n_316), .B(n_399), .Y(n_398) );
INVx3_ASAP7_75t_L g415 ( .A(n_316), .Y(n_415) );
INVx1_ASAP7_75t_L g484 ( .A(n_317), .Y(n_484) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x4_ASAP7_75t_L g348 ( .A(n_318), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g390 ( .A(n_320), .B(n_339), .Y(n_390) );
AND2x2_ASAP7_75t_L g416 ( .A(n_320), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OR2x2_ASAP7_75t_L g426 ( .A(n_321), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_343), .Y(n_322) );
A2O1A1Ixp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B(n_333), .C(n_334), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_326), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_327), .B(n_374), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g395 ( .A(n_327), .B(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_328), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g349 ( .A(n_329), .B(n_336), .Y(n_349) );
INVx1_ASAP7_75t_L g404 ( .A(n_329), .Y(n_404) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_337), .B(n_340), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g405 ( .A(n_336), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g417 ( .A(n_339), .Y(n_417) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x4_ASAP7_75t_L g441 ( .A(n_342), .B(n_409), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_353), .Y(n_343) );
A2O1A1Ixp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_346), .B(n_348), .C(n_350), .Y(n_344) );
BUFx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g408 ( .A(n_347), .B(n_409), .Y(n_408) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI21xp5_ASAP7_75t_SL g353 ( .A1(n_354), .A2(n_356), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_359), .Y(n_368) );
OR2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g469 ( .A(n_359), .Y(n_469) );
AOI222xp33_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_365), .B1(n_366), .B2(n_369), .C1(n_371), .C2(n_372), .Y(n_360) );
NOR2x1_ASAP7_75t_L g378 ( .A(n_362), .B(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_363), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g374 ( .A(n_364), .Y(n_374) );
INVx1_ASAP7_75t_L g472 ( .A(n_364), .Y(n_472) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_367), .B(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g450 ( .A(n_367), .Y(n_450) );
AND2x4_ASAP7_75t_L g457 ( .A(n_367), .B(n_434), .Y(n_457) );
INVx2_ASAP7_75t_L g486 ( .A(n_367), .Y(n_486) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_370), .A2(n_423), .B1(n_426), .B2(n_428), .Y(n_422) );
AOI211xp5_ASAP7_75t_L g476 ( .A1(n_372), .A2(n_477), .B(n_478), .C(n_482), .Y(n_476) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR2xp67_ASAP7_75t_SL g375 ( .A(n_376), .B(n_437), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_394), .C(n_401), .D(n_421), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_383), .B(n_384), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI22xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_387), .B1(n_389), .B2(n_391), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_388), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_389), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g399 ( .A(n_393), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_400), .Y(n_397) );
INVx1_ASAP7_75t_L g424 ( .A(n_400), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_408), .B1(n_410), .B2(n_416), .C(n_418), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_407), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_403), .B(n_419), .Y(n_418) );
OR2x2_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
AND2x2_ASAP7_75t_L g456 ( .A(n_404), .B(n_431), .Y(n_456) );
INVx2_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
NAND2x1_ASAP7_75t_SL g411 ( .A(n_412), .B(n_414), .Y(n_411) );
INVx1_ASAP7_75t_L g481 ( .A(n_412), .Y(n_481) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g483 ( .A(n_420), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_429), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g465 ( .A(n_427), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_435), .B2(n_436), .Y(n_429) );
AND2x2_ASAP7_75t_L g462 ( .A(n_431), .B(n_448), .Y(n_462) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g443 ( .A(n_436), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_453), .C(n_476), .Y(n_437) );
AOI222xp33_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_443), .B1(n_444), .B2(n_450), .C1(n_451), .C2(n_452), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B(n_458), .C(n_470), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_461), .B1(n_463), .B2(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_469), .Y(n_467) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_484), .B1(n_485), .B2(n_487), .Y(n_482) );
INVx4_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_490), .Y(n_492) );
AND2x2_ASAP7_75t_L g837 ( .A(n_490), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_SL g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g821 ( .A(n_493), .Y(n_821) );
AND2x4_ASAP7_75t_L g493 ( .A(n_494), .B(n_719), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_648), .C(n_690), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_622), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_535), .B1(n_597), .B2(n_608), .Y(n_496) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_522), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_499), .A2(n_642), .B(n_644), .Y(n_641) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_499), .A2(n_715), .B(n_716), .Y(n_714) );
OR2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_511), .Y(n_499) );
INVx2_ASAP7_75t_L g634 ( .A(n_500), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_500), .B(n_512), .Y(n_664) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
OAI21xp33_ASAP7_75t_SL g541 ( .A1(n_504), .A2(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g605 ( .A(n_505), .Y(n_605) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_508), .B(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g607 ( .A(n_510), .Y(n_607) );
AND2x2_ASAP7_75t_L g704 ( .A(n_511), .B(n_552), .Y(n_704) );
INVx1_ASAP7_75t_L g737 ( .A(n_511), .Y(n_737) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g599 ( .A(n_512), .B(n_553), .Y(n_599) );
AND2x2_ASAP7_75t_L g630 ( .A(n_512), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g639 ( .A(n_512), .Y(n_639) );
OR2x2_ASAP7_75t_L g658 ( .A(n_512), .B(n_524), .Y(n_658) );
AND2x2_ASAP7_75t_L g673 ( .A(n_512), .B(n_524), .Y(n_673) );
INVx4_ASAP7_75t_L g516 ( .A(n_515), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_518), .B(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g533 ( .A(n_519), .Y(n_533) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_523), .B(n_672), .Y(n_715) );
OR2x2_ASAP7_75t_L g803 ( .A(n_523), .B(n_664), .Y(n_803) );
INVx1_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g631 ( .A(n_524), .Y(n_631) );
AND2x2_ASAP7_75t_L g640 ( .A(n_524), .B(n_603), .Y(n_640) );
AND2x2_ASAP7_75t_L g643 ( .A(n_524), .B(n_553), .Y(n_643) );
AND2x2_ASAP7_75t_L g662 ( .A(n_524), .B(n_552), .Y(n_662) );
AND2x4_ASAP7_75t_L g681 ( .A(n_524), .B(n_604), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_529), .B(n_533), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_550), .B(n_585), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_536), .B(n_676), .Y(n_779) );
CKINVDCx14_ASAP7_75t_R g536 ( .A(n_537), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_538), .B(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g612 ( .A(n_538), .Y(n_612) );
OR2x2_ASAP7_75t_L g620 ( .A(n_538), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_538), .B(n_613), .Y(n_645) );
AND2x2_ASAP7_75t_L g670 ( .A(n_538), .B(n_587), .Y(n_670) );
AND2x2_ASAP7_75t_L g688 ( .A(n_538), .B(n_618), .Y(n_688) );
INVx1_ASAP7_75t_L g727 ( .A(n_538), .Y(n_727) );
AND2x2_ASAP7_75t_L g729 ( .A(n_538), .B(n_730), .Y(n_729) );
NAND2x1p5_ASAP7_75t_SL g748 ( .A(n_538), .B(n_669), .Y(n_748) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OAI21xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_546), .B(n_549), .Y(n_540) );
OAI32xp33_ASAP7_75t_L g632 ( .A1(n_550), .A2(n_624), .A3(n_633), .B1(n_635), .B2(n_637), .Y(n_632) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_564), .Y(n_550) );
INVx1_ASAP7_75t_L g672 ( .A(n_551), .Y(n_672) );
AND2x2_ASAP7_75t_L g680 ( .A(n_551), .B(n_681), .Y(n_680) );
BUFx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g679 ( .A(n_552), .B(n_603), .Y(n_679) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g629 ( .A(n_553), .Y(n_629) );
AND2x2_ASAP7_75t_L g638 ( .A(n_553), .B(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g744 ( .A(n_553), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
OAI21x1_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_559), .B(n_562), .Y(n_555) );
INVx2_ASAP7_75t_L g614 ( .A(n_564), .Y(n_614) );
OR2x2_ASAP7_75t_L g624 ( .A(n_564), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g746 ( .A(n_564), .Y(n_746) );
OR2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_578), .Y(n_564) );
AND2x2_ASAP7_75t_L g647 ( .A(n_565), .B(n_579), .Y(n_647) );
INVx2_ASAP7_75t_L g669 ( .A(n_565), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_565), .B(n_587), .Y(n_689) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g596 ( .A(n_566), .Y(n_596) );
AOI21x1_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_568), .B(n_577), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_578), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g678 ( .A(n_578), .Y(n_678) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
BUFx2_ASAP7_75t_L g618 ( .A(n_579), .Y(n_618) );
OR2x2_ASAP7_75t_L g684 ( .A(n_579), .B(n_587), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_579), .B(n_587), .Y(n_717) );
INVx2_ASAP7_75t_L g665 ( .A(n_585), .Y(n_665) );
OR2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_595), .Y(n_585) );
OR2x2_ASAP7_75t_L g652 ( .A(n_586), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g730 ( .A(n_586), .Y(n_730) );
INVx1_ASAP7_75t_L g613 ( .A(n_587), .Y(n_613) );
INVx1_ASAP7_75t_L g621 ( .A(n_587), .Y(n_621) );
INVx1_ASAP7_75t_L g636 ( .A(n_587), .Y(n_636) );
OR2x2_ASAP7_75t_L g740 ( .A(n_595), .B(n_717), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_596), .B(n_612), .Y(n_653) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_596), .Y(n_655) );
OR2x2_ASAP7_75t_L g754 ( .A(n_596), .B(n_678), .Y(n_754) );
INVxp67_ASAP7_75t_L g778 ( .A(n_596), .Y(n_778) );
INVx2_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NAND2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_599), .B(n_640), .Y(n_707) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g656 ( .A(n_601), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g769 ( .A(n_602), .Y(n_769) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g798 ( .A(n_603), .B(n_631), .Y(n_798) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g724 ( .A(n_604), .B(n_631), .Y(n_724) );
AOI21x1_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B(n_607), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_615), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_611), .B(n_647), .Y(n_761) );
AND2x4_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx2_ASAP7_75t_L g625 ( .A(n_612), .Y(n_625) );
AND2x2_ASAP7_75t_L g675 ( .A(n_612), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_612), .B(n_669), .Y(n_718) );
OR2x2_ASAP7_75t_L g790 ( .A(n_612), .B(n_677), .Y(n_790) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g710 ( .A(n_616), .B(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx2_ASAP7_75t_L g701 ( .A(n_617), .Y(n_701) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g691 ( .A(n_620), .B(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_SL g702 ( .A(n_620), .Y(n_702) );
OR2x2_ASAP7_75t_L g753 ( .A(n_620), .B(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g808 ( .A(n_620), .Y(n_808) );
AOI211xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_632), .C(n_641), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g697 ( .A(n_625), .B(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_625), .B(n_746), .Y(n_745) );
AND2x2_ASAP7_75t_L g770 ( .A(n_625), .B(n_647), .Y(n_770) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_628), .B(n_673), .Y(n_695) );
NAND2x1p5_ASAP7_75t_L g712 ( .A(n_628), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g780 ( .A(n_628), .B(n_781), .Y(n_780) );
INVx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g723 ( .A(n_629), .Y(n_723) );
AND2x2_ASAP7_75t_L g751 ( .A(n_630), .B(n_679), .Y(n_751) );
INVx2_ASAP7_75t_L g774 ( .A(n_630), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_630), .B(n_672), .Y(n_806) );
AND2x4_ASAP7_75t_SL g760 ( .A(n_633), .B(n_638), .Y(n_760) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g713 ( .A(n_634), .B(n_639), .Y(n_713) );
OR2x2_ASAP7_75t_L g765 ( .A(n_634), .B(n_658), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_635), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_635), .B(n_647), .Y(n_801) );
BUFx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g749 ( .A(n_636), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx1_ASAP7_75t_L g732 ( .A(n_638), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_638), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g782 ( .A(n_639), .Y(n_782) );
BUFx2_ASAP7_75t_L g650 ( .A(n_640), .Y(n_650) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g768 ( .A(n_643), .B(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g692 ( .A(n_647), .Y(n_692) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_647), .Y(n_709) );
NAND3xp33_ASAP7_75t_SL g648 ( .A(n_649), .B(n_659), .C(n_674), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_651), .B1(n_654), .B2(n_656), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI222xp33_ASAP7_75t_L g762 ( .A1(n_656), .A2(n_682), .B1(n_763), .B2(n_766), .C1(n_768), .C2(n_770), .Y(n_762) );
AND2x2_ASAP7_75t_L g794 ( .A(n_657), .B(n_743), .Y(n_794) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g742 ( .A(n_658), .B(n_743), .Y(n_742) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_665), .B1(n_666), .B2(n_671), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
INVx2_ASAP7_75t_SL g738 ( .A(n_662), .Y(n_738) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
AND2x2_ASAP7_75t_L g725 ( .A(n_667), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g683 ( .A(n_668), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g677 ( .A(n_669), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g792 ( .A(n_670), .Y(n_792) );
AND2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_673), .B(n_769), .Y(n_788) );
INVx1_ASAP7_75t_L g805 ( .A(n_673), .Y(n_805) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_679), .B1(n_680), .B2(n_682), .C1(n_685), .C2(n_686), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_681), .Y(n_685) );
AND2x2_ASAP7_75t_L g703 ( .A(n_681), .B(n_704), .Y(n_703) );
INVx3_ASAP7_75t_L g734 ( .A(n_681), .Y(n_734) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g698 ( .A(n_684), .Y(n_698) );
OR2x2_ASAP7_75t_L g767 ( .A(n_684), .B(n_748), .Y(n_767) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_689), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B(n_696), .C(n_705), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_697), .A2(n_699), .B(n_703), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g783 ( .A1(n_697), .A2(n_735), .B1(n_784), .B2(n_787), .C(n_789), .Y(n_783) );
AND2x4_ASAP7_75t_L g726 ( .A(n_698), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_L g757 ( .A(n_704), .Y(n_757) );
AOI211x1_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B(n_710), .C(n_714), .Y(n_705) );
INVxp67_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g775 ( .A(n_713), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g763 ( .A(n_716), .B(n_764), .C(n_765), .Y(n_763) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g799 ( .A(n_717), .Y(n_799) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_771), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g720 ( .A(n_721), .B(n_728), .C(n_750), .D(n_762), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
AND2x2_ASAP7_75t_L g781 ( .A(n_724), .B(n_782), .Y(n_781) );
AOI221x1_ASAP7_75t_L g750 ( .A1(n_726), .A2(n_751), .B1(n_752), .B2(n_755), .C(n_758), .Y(n_750) );
AND2x2_ASAP7_75t_L g776 ( .A(n_726), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g786 ( .A(n_727), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_731), .B1(n_735), .B2(n_739), .C(n_741), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_733), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
OR2x2_ASAP7_75t_L g736 ( .A(n_737), .B(n_738), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_738), .A2(n_742), .B1(n_745), .B2(n_747), .Y(n_741) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_742), .A2(n_759), .B(n_761), .Y(n_758) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g764 ( .A(n_744), .Y(n_764) );
OR2x2_ASAP7_75t_L g747 ( .A(n_748), .B(n_749), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVxp67_ASAP7_75t_L g785 ( .A(n_754), .Y(n_785) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g804 ( .A1(n_767), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_783), .C(n_795), .Y(n_771) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_776), .B1(n_779), .B2(n_780), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
OR2x2_ASAP7_75t_L g791 ( .A(n_778), .B(n_792), .Y(n_791) );
NAND2x1_ASAP7_75t_L g807 ( .A(n_778), .B(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx2_ASAP7_75t_SL g787 ( .A(n_788), .Y(n_787) );
AOI21xp5_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_791), .B(n_793), .Y(n_789) );
INVx1_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
AOI221xp5_ASAP7_75t_L g795 ( .A1(n_796), .A2(n_799), .B1(n_800), .B2(n_802), .C(n_804), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx3_ASAP7_75t_R g802 ( .A(n_803), .Y(n_802) );
CKINVDCx16_ASAP7_75t_R g809 ( .A(n_810), .Y(n_809) );
BUFx12f_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AND2x6_ASAP7_75t_SL g811 ( .A(n_812), .B(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx3_ASAP7_75t_L g831 ( .A(n_813), .Y(n_831) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_813), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
OAI21xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_822), .B(n_828), .Y(n_818) );
INVx4_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx12f_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx4_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g829 ( .A(n_830), .Y(n_829) );
BUFx8_ASAP7_75t_SL g830 ( .A(n_831), .Y(n_830) );
INVx2_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx10_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
CKINVDCx11_ASAP7_75t_R g839 ( .A(n_840), .Y(n_839) );
endmodule