module fake_netlist_6_4924_n_2092 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2092);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2092;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_2016;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_2050;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_53),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_184),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_68),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_64),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_113),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_10),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_164),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_109),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_85),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_28),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_205),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_204),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_6),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_96),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_128),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_61),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_51),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_180),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_22),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_153),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_34),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_112),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_1),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_157),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_94),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_142),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_70),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_119),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_73),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_72),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_192),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_76),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_133),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_17),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_70),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_110),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_60),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_67),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_81),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_92),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_167),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_121),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_114),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_3),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_216),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_98),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_14),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_64),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_108),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_14),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_13),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_134),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_150),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_210),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_33),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_71),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_46),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_197),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_46),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_61),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_177),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_124),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_33),
.Y(n_293)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_52),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_189),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_132),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_154),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_179),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_95),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_123),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_17),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_139),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_54),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_50),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_146),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_141),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_44),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_116),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_59),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_111),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_182),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_58),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_2),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_29),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_115),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_209),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_49),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_48),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_158),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_208),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_87),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_79),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_68),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_84),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_178),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_88),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g330 ( 
.A(n_49),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_72),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_102),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_163),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_41),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_171),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_86),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_37),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_203),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_195),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_214),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_151),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_25),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_202),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_104),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_91),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_155),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_90),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_159),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_168),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_8),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_24),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_0),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_65),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_74),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_126),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_22),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_34),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_135),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_5),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_4),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_59),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_41),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_56),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_106),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_19),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_117),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_38),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_15),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_20),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_82),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_127),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_43),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_36),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_131),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_143),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_103),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_190),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_0),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_77),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_3),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_100),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_107),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_39),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_32),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_74),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_69),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_2),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_12),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_170),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_67),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_207),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_48),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_185),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_43),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_25),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_211),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_144),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_93),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_125),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_186),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_26),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_26),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_55),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_58),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_129),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_5),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_40),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_130),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_188),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_57),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_183),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_173),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_39),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_57),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_35),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_63),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_175),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_149),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_201),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_53),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_191),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_42),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_21),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_194),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_105),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_101),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_36),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_28),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_62),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_230),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_313),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_313),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_219),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_250),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_225),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_225),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_225),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_225),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_253),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_225),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_305),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_255),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_242),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_277),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_260),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_261),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_R g447 ( 
.A(n_292),
.B(n_78),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_277),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_327),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_277),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_277),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_283),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_263),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_277),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_347),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_254),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_304),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_304),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_304),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_270),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_273),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_304),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_304),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_275),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_402),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_257),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_258),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_283),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_265),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_284),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_402),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_266),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_267),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_330),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_283),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_218),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_236),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_303),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_310),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_240),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_246),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_252),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_314),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_232),
.B(n_7),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_256),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_290),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_315),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g491 ( 
.A(n_220),
.B(n_7),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_268),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_316),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_233),
.B(n_8),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_224),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_264),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_380),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_290),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_274),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_278),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_233),
.B(n_9),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_319),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_282),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_269),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g505 ( 
.A(n_291),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_320),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_326),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_334),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_259),
.B(n_10),
.Y(n_509)
);

INVxp67_ASAP7_75t_SL g510 ( 
.A(n_329),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_325),
.B(n_361),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_383),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_363),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_365),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_272),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_276),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_368),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_342),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_383),
.Y(n_519)
);

CKINVDCx16_ASAP7_75t_R g520 ( 
.A(n_383),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_373),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_350),
.Y(n_522)
);

NOR2xp67_ASAP7_75t_L g523 ( 
.A(n_354),
.B(n_11),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_279),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_390),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_401),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_406),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_351),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g530 ( 
.A(n_285),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_352),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_414),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_415),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_423),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_353),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_329),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_389),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_259),
.B(n_11),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_356),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_271),
.B(n_397),
.Y(n_540)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_217),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_222),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_271),
.B(n_12),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_357),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_231),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_359),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_238),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_458),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_459),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_459),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_456),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_463),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_439),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_463),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_489),
.B(n_293),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_478),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_541),
.B(n_262),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g561 ( 
.A(n_439),
.B(n_245),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_467),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_468),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_262),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_545),
.B(n_297),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_478),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_442),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_435),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_471),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_430),
.B(n_375),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_437),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_495),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_495),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_474),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_475),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_438),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_492),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_498),
.B(n_293),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_504),
.Y(n_580)
);

CKINVDCx16_ASAP7_75t_R g581 ( 
.A(n_452),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_442),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_433),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_547),
.B(n_297),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_495),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_444),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_443),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_515),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_448),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_516),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_524),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_445),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_451),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_454),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_457),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_462),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_465),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_449),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_530),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_431),
.Y(n_604)
);

OA21x2_ASAP7_75t_L g605 ( 
.A1(n_466),
.A2(n_281),
.B(n_247),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_445),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_470),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_430),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_446),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_446),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_473),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_453),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_453),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_543),
.B(n_296),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_540),
.B(n_537),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_460),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_460),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_455),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_461),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_480),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_432),
.B(n_337),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_483),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_484),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_485),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_476),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_488),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_461),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_496),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_500),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_434),
.B(n_298),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_513),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_464),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_514),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_517),
.Y(n_637)
);

CKINVDCx20_ASAP7_75t_R g638 ( 
.A(n_469),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_521),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_477),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_623),
.Y(n_641)
);

INVxp67_ASAP7_75t_SL g642 ( 
.A(n_586),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_623),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_614),
.B(n_224),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_568),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_583),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_614),
.B(n_487),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_616),
.A2(n_494),
.B1(n_509),
.B2(n_501),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_614),
.B(n_538),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_555),
.B(n_520),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_604),
.B(n_464),
.Y(n_652)
);

OR2x6_ASAP7_75t_L g653 ( 
.A(n_556),
.B(n_512),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_624),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_597),
.B(n_525),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_560),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_624),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_553),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_629),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_588),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_551),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_604),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_614),
.A2(n_301),
.B1(n_360),
.B2(n_337),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_629),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_560),
.B(n_527),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_560),
.B(n_472),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_632),
.B(n_472),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_558),
.B(n_224),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_558),
.B(n_481),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_560),
.B(n_224),
.Y(n_672)
);

INVxp67_ASAP7_75t_SL g673 ( 
.A(n_586),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_631),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_605),
.A2(n_301),
.B1(n_360),
.B2(n_491),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_561),
.B(n_224),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_579),
.B(n_481),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_551),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_551),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_568),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_574),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_556),
.B(n_348),
.Y(n_682)
);

AND3x2_ASAP7_75t_L g683 ( 
.A(n_608),
.B(n_519),
.C(n_441),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_579),
.B(n_482),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_634),
.B(n_348),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_574),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_571),
.A2(n_486),
.B1(n_490),
.B2(n_482),
.Y(n_687)
);

AND2x6_ASAP7_75t_L g688 ( 
.A(n_622),
.B(n_348),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_486),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_634),
.B(n_348),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_567),
.B(n_490),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_634),
.B(n_493),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_554),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_622),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_631),
.Y(n_695)
);

INVx8_ASAP7_75t_L g696 ( 
.A(n_609),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_633),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_634),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_634),
.B(n_493),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_605),
.A2(n_523),
.B1(n_511),
.B2(n_497),
.Y(n_700)
);

NAND2xp33_ASAP7_75t_R g701 ( 
.A(n_610),
.B(n_502),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_586),
.B(n_502),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_634),
.B(n_348),
.Y(n_703)
);

OAI22xp5_ASAP7_75t_L g704 ( 
.A1(n_608),
.A2(n_507),
.B1(n_508),
.B2(n_506),
.Y(n_704)
);

BUFx3_ASAP7_75t_L g705 ( 
.A(n_639),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_639),
.B(n_355),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_574),
.Y(n_707)
);

BUFx4f_ASAP7_75t_L g708 ( 
.A(n_639),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_582),
.B(n_507),
.C(n_506),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_581),
.B(n_508),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_605),
.A2(n_511),
.B1(n_528),
.B2(n_532),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_633),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_554),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_612),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_574),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_639),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_595),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_639),
.B(n_355),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_636),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_639),
.B(n_518),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_636),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_564),
.B(n_533),
.Y(n_723)
);

INVxp67_ASAP7_75t_L g724 ( 
.A(n_606),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_627),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_557),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_620),
.A2(n_546),
.B1(n_544),
.B2(n_539),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_613),
.A2(n_546),
.B1(n_544),
.B2(n_539),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_617),
.B(n_518),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_593),
.Y(n_730)
);

XOR2xp5_ASAP7_75t_L g731 ( 
.A(n_602),
.B(n_619),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_574),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_564),
.B(n_355),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_581),
.B(n_522),
.Y(n_734)
);

BUFx4f_ASAP7_75t_L g735 ( 
.A(n_564),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_618),
.A2(n_535),
.B1(n_531),
.B2(n_529),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_564),
.B(n_355),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_573),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_627),
.B(n_522),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_627),
.Y(n_740)
);

AND3x2_ASAP7_75t_L g741 ( 
.A(n_565),
.B(n_318),
.C(n_307),
.Y(n_741)
);

OR2x2_ASAP7_75t_L g742 ( 
.A(n_627),
.B(n_529),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_630),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_628),
.B(n_531),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_635),
.B(n_535),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_630),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_565),
.B(n_355),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_593),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_630),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_565),
.B(n_526),
.C(n_534),
.Y(n_750)
);

AND2x6_ASAP7_75t_L g751 ( 
.A(n_565),
.B(n_321),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_630),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_559),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_590),
.B(n_280),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_584),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_605),
.B(n_322),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_615),
.B(n_505),
.Y(n_757)
);

NAND2x1p5_ASAP7_75t_L g758 ( 
.A(n_584),
.B(n_345),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_570),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_638),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_570),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_590),
.B(n_399),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_572),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_584),
.B(n_447),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_559),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_SL g766 ( 
.A(n_584),
.B(n_385),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_593),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_572),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_566),
.Y(n_769)
);

BUFx4f_ASAP7_75t_L g770 ( 
.A(n_593),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_615),
.A2(n_333),
.B1(n_332),
.B2(n_328),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_577),
.Y(n_772)
);

AND2x6_ASAP7_75t_L g773 ( 
.A(n_548),
.B(n_323),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_577),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_621),
.B(n_244),
.Y(n_775)
);

INVx4_ASAP7_75t_SL g776 ( 
.A(n_573),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_573),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_585),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_621),
.B(n_324),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_585),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_625),
.B(n_287),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_625),
.B(n_289),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_573),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_590),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_640),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_587),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_566),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_590),
.B(n_548),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_587),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_637),
.B(n_367),
.C(n_362),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_573),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_573),
.Y(n_792)
);

AND2x4_ASAP7_75t_L g793 ( 
.A(n_637),
.B(n_376),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_591),
.B(n_400),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_549),
.Y(n_795)
);

INVx4_ASAP7_75t_SL g796 ( 
.A(n_611),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_591),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_596),
.B(n_223),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_735),
.B(n_396),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_755),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_735),
.B(n_396),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_669),
.B(n_294),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_657),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_755),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_704),
.B(n_563),
.C(n_562),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_756),
.A2(n_308),
.B1(n_394),
.B2(n_422),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_657),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_659),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_739),
.B(n_549),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_669),
.B(n_223),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_646),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_641),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_648),
.B(n_550),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_650),
.A2(n_649),
.B(n_664),
.C(n_671),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_643),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_671),
.B(n_226),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_692),
.B(n_552),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_757),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_680),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_680),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_693),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_781),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_655),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_658),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_660),
.Y(n_826)
);

AND3x1_ASAP7_75t_L g827 ( 
.A(n_684),
.B(n_412),
.C(n_408),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_692),
.B(n_699),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_667),
.A2(n_426),
.B1(n_425),
.B2(n_424),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_782),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_693),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_699),
.B(n_721),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_665),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_721),
.B(n_552),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_756),
.B(n_663),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_684),
.B(n_396),
.Y(n_836)
);

AND2x6_ASAP7_75t_SL g837 ( 
.A(n_653),
.B(n_421),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_675),
.B(n_598),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_677),
.B(n_396),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_674),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_666),
.B(n_598),
.Y(n_841)
);

AOI22xp5_ASAP7_75t_L g842 ( 
.A1(n_652),
.A2(n_286),
.B1(n_288),
.B2(n_295),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_775),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_695),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_708),
.A2(n_600),
.B(n_599),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_713),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_742),
.B(n_226),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_713),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_694),
.B(n_227),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_SL g850 ( 
.A(n_691),
.B(n_221),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_654),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_694),
.B(n_227),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_720),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_729),
.B(n_569),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_666),
.B(n_599),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_700),
.B(n_396),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_700),
.B(n_396),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_708),
.A2(n_673),
.B(n_642),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_666),
.B(n_600),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_654),
.Y(n_860)
);

NOR2xp33_ASAP7_75t_L g861 ( 
.A(n_689),
.B(n_228),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_664),
.A2(n_410),
.B(n_416),
.C(n_331),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_645),
.A2(n_396),
.B1(n_407),
.B2(n_387),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_725),
.B(n_396),
.Y(n_864)
);

AOI22x1_ASAP7_75t_L g865 ( 
.A1(n_740),
.A2(n_239),
.B1(n_391),
.B2(n_393),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_723),
.B(n_607),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_743),
.B(n_746),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_697),
.B(n_712),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_702),
.B(n_228),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_701),
.Y(n_870)
);

NAND2xp33_ASAP7_75t_L g871 ( 
.A(n_751),
.B(n_299),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_719),
.B(n_607),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_749),
.B(n_300),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_723),
.B(n_229),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_709),
.B(n_229),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_720),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_726),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_L g879 ( 
.A(n_736),
.B(n_576),
.C(n_575),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_759),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_761),
.Y(n_881)
);

AO221x1_ASAP7_75t_L g882 ( 
.A1(n_727),
.A2(n_724),
.B1(n_752),
.B2(n_763),
.C(n_774),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_768),
.Y(n_883)
);

A2O1A1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_711),
.A2(n_243),
.B(n_248),
.C(n_241),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_726),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_758),
.B(n_302),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_682),
.B(n_764),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_687),
.B(n_235),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_772),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_778),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_682),
.B(n_601),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_764),
.A2(n_249),
.B1(n_251),
.B2(n_239),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_758),
.B(n_306),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_780),
.B(n_601),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_744),
.B(n_578),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_651),
.B(n_580),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_711),
.B(n_795),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_786),
.B(n_601),
.Y(n_898)
);

NOR2xp67_ASAP7_75t_L g899 ( 
.A(n_728),
.B(n_589),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_789),
.B(n_601),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_797),
.B(n_611),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_795),
.B(n_309),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_656),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_753),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_754),
.B(n_311),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_762),
.B(n_312),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_670),
.B(n_611),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_656),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_766),
.A2(n_377),
.B1(n_336),
.B2(n_338),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_653),
.B(n_798),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_670),
.B(n_611),
.Y(n_911)
);

NAND2xp33_ASAP7_75t_SL g912 ( 
.A(n_717),
.B(n_701),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_653),
.B(n_592),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_765),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_645),
.B(n_611),
.Y(n_915)
);

INVx8_ASAP7_75t_L g916 ( 
.A(n_696),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_798),
.B(n_235),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_765),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_656),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_SL g920 ( 
.A(n_714),
.B(n_594),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_770),
.A2(n_343),
.B(n_370),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_784),
.B(n_317),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_770),
.A2(n_791),
.B(n_672),
.Y(n_923)
);

AND2x6_ASAP7_75t_SL g924 ( 
.A(n_745),
.B(n_221),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_672),
.B(n_723),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_788),
.B(n_335),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_731),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_794),
.B(n_339),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_794),
.B(n_340),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_769),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_787),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_794),
.B(n_341),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_710),
.B(n_734),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_696),
.Y(n_934)
);

AO221x1_ASAP7_75t_L g935 ( 
.A1(n_738),
.A2(n_792),
.B1(n_777),
.B2(n_732),
.C(n_681),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_766),
.B(n_237),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_771),
.A2(n_391),
.B1(n_237),
.B2(n_249),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_779),
.A2(n_358),
.B(n_349),
.C(n_346),
.Y(n_938)
);

BUFx8_ASAP7_75t_L g939 ( 
.A(n_793),
.Y(n_939)
);

OAI22xp33_ASAP7_75t_L g940 ( 
.A1(n_750),
.A2(n_387),
.B1(n_429),
.B2(n_428),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_793),
.Y(n_941)
);

NOR2xp67_ASAP7_75t_L g942 ( 
.A(n_790),
.B(n_603),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_793),
.B(n_344),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_698),
.B(n_364),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_705),
.B(n_366),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_644),
.Y(n_946)
);

OR2x6_ASAP7_75t_L g947 ( 
.A(n_696),
.B(n_375),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_733),
.A2(n_374),
.B(n_379),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_779),
.B(n_251),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_751),
.A2(n_676),
.B1(n_688),
.B2(n_773),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_705),
.B(n_371),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_733),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_737),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_760),
.B(n_647),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_716),
.B(n_381),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_661),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_737),
.B(n_375),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_771),
.A2(n_429),
.B1(n_428),
.B2(n_427),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_382),
.B1(n_398),
.B2(n_419),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_747),
.Y(n_960)
);

OR2x6_ASAP7_75t_L g961 ( 
.A(n_747),
.B(n_15),
.Y(n_961)
);

O2A1O1Ixp5_ASAP7_75t_L g962 ( 
.A1(n_836),
.A2(n_676),
.B(n_690),
.C(n_703),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_897),
.A2(n_706),
.B(n_718),
.Y(n_963)
);

BUFx2_ASAP7_75t_L g964 ( 
.A(n_956),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_836),
.A2(n_801),
.B(n_799),
.C(n_839),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_828),
.B(n_751),
.Y(n_966)
);

AOI22xp33_ASAP7_75t_L g967 ( 
.A1(n_802),
.A2(n_773),
.B1(n_688),
.B2(n_716),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_811),
.A2(n_773),
.B1(n_688),
.B2(n_678),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_910),
.B(n_843),
.Y(n_969)
);

O2A1O1Ixp5_ASAP7_75t_L g970 ( 
.A1(n_799),
.A2(n_685),
.B(n_690),
.C(n_703),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_897),
.A2(n_857),
.B(n_856),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_851),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_800),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_856),
.A2(n_685),
.B(n_706),
.Y(n_974)
);

AND3x2_ASAP7_75t_L g975 ( 
.A(n_888),
.B(n_785),
.C(n_683),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_910),
.B(n_393),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_SL g977 ( 
.A(n_803),
.B(n_398),
.Y(n_977)
);

CKINVDCx10_ASAP7_75t_R g978 ( 
.A(n_927),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_857),
.A2(n_718),
.B(n_776),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_823),
.B(n_234),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_808),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_835),
.A2(n_925),
.B(n_838),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_954),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_815),
.A2(n_409),
.B1(n_419),
.B2(n_418),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_803),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_917),
.B(n_668),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_817),
.B(n_405),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_830),
.B(n_847),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_815),
.A2(n_405),
.B1(n_418),
.B2(n_417),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_884),
.A2(n_678),
.B(n_679),
.C(n_681),
.Y(n_990)
);

AOI21x1_ASAP7_75t_L g991 ( 
.A1(n_867),
.A2(n_776),
.B(n_732),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_817),
.A2(n_409),
.B(n_411),
.C(n_417),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_809),
.Y(n_993)
);

OA21x2_ASAP7_75t_L g994 ( 
.A1(n_935),
.A2(n_411),
.B(n_773),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_923),
.A2(n_730),
.B(n_748),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_884),
.A2(n_679),
.B(n_777),
.C(n_738),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_814),
.B(n_792),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_858),
.A2(n_767),
.B(n_644),
.Y(n_998)
);

INVxp67_ASAP7_75t_L g999 ( 
.A(n_861),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_870),
.B(n_369),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_888),
.B(n_372),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_933),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_887),
.A2(n_767),
.B(n_686),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_847),
.B(n_644),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_835),
.A2(n_644),
.B(n_715),
.Y(n_1005)
);

INVx4_ASAP7_75t_L g1006 ( 
.A(n_916),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_810),
.B(n_686),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_819),
.B(n_378),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_812),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_820),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_849),
.B(n_234),
.Y(n_1011)
);

AO21x1_ASAP7_75t_L g1012 ( 
.A1(n_801),
.A2(n_16),
.B(n_18),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_861),
.B(n_384),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_869),
.B(n_686),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_869),
.B(n_715),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_807),
.B(n_715),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_862),
.A2(n_741),
.B(n_243),
.C(n_248),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_807),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_818),
.B(n_834),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_939),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_806),
.B(n_241),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_839),
.A2(n_783),
.B(n_662),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_804),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_813),
.B(n_816),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_867),
.A2(n_783),
.B(n_707),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_939),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_916),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_936),
.A2(n_386),
.B(n_331),
.C(n_388),
.Y(n_1028)
);

BUFx4f_ASAP7_75t_L g1029 ( 
.A(n_916),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_849),
.B(n_388),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_821),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_915),
.A2(n_898),
.B(n_894),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_900),
.A2(n_783),
.B(n_707),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_824),
.B(n_776),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_912),
.B(n_796),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_868),
.A2(n_707),
.B(n_662),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_961),
.Y(n_1037)
);

OAI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_952),
.A2(n_392),
.B1(n_395),
.B2(n_403),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_875),
.B(n_392),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_875),
.B(n_395),
.Y(n_1040)
);

AOI21x1_ASAP7_75t_L g1041 ( 
.A1(n_907),
.A2(n_796),
.B(n_707),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_953),
.A2(n_403),
.B1(n_404),
.B2(n_427),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_825),
.B(n_796),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_826),
.B(n_662),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_L g1045 ( 
.A(n_934),
.B(n_80),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_936),
.A2(n_420),
.B(n_416),
.C(n_410),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_841),
.A2(n_662),
.B(n_420),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_833),
.B(n_404),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_855),
.A2(n_407),
.B(n_89),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_852),
.B(n_16),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_911),
.A2(n_97),
.B(n_212),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_822),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_862),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_1053)
);

OAI22xp5_ASAP7_75t_L g1054 ( 
.A1(n_960),
.A2(n_99),
.B1(n_206),
.B2(n_200),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_859),
.A2(n_83),
.B(n_196),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_901),
.A2(n_215),
.B(n_187),
.Y(n_1056)
);

AOI21x1_ASAP7_75t_L g1057 ( 
.A1(n_891),
.A2(n_181),
.B(n_174),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_864),
.A2(n_169),
.B(n_166),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_L g1059 ( 
.A(n_806),
.B(n_21),
.C(n_23),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_827),
.B(n_866),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_874),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_944),
.A2(n_165),
.B(n_162),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_945),
.A2(n_160),
.B(n_156),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_852),
.B(n_896),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_829),
.A2(n_23),
.B(n_24),
.C(n_27),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_946),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_854),
.B(n_27),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_866),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_951),
.A2(n_152),
.B(n_147),
.Y(n_1069)
);

CKINVDCx8_ASAP7_75t_R g1070 ( 
.A(n_924),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_946),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_860),
.B(n_145),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_895),
.B(n_29),
.Y(n_1073)
);

NAND3xp33_ASAP7_75t_L g1074 ( 
.A(n_842),
.B(n_30),
.C(n_31),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_874),
.B(n_30),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_882),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_1076)
);

AO21x1_ASAP7_75t_L g1077 ( 
.A1(n_886),
.A2(n_38),
.B(n_42),
.Y(n_1077)
);

OAI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_930),
.A2(n_140),
.B(n_137),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_946),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_955),
.A2(n_136),
.B(n_122),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_913),
.B(n_45),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_903),
.B(n_45),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_946),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_922),
.A2(n_120),
.B(n_118),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_840),
.B(n_47),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_961),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_908),
.B(n_47),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_941),
.A2(n_50),
.B(n_52),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_926),
.A2(n_54),
.B(n_55),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_831),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_871),
.A2(n_56),
.B(n_62),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_919),
.A2(n_877),
.B1(n_890),
.B2(n_889),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_920),
.B(n_63),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_961),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_863),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_850),
.B(n_66),
.C(n_71),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_844),
.A2(n_75),
.B1(n_883),
.B2(n_881),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_949),
.A2(n_75),
.B(n_880),
.C(n_863),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_SL g1099 ( 
.A(n_928),
.B(n_932),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_949),
.B(n_872),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_846),
.B(n_876),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_848),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_853),
.Y(n_1103)
);

INVx4_ASAP7_75t_L g1104 ( 
.A(n_878),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_943),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_929),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_873),
.A2(n_905),
.B(n_906),
.Y(n_1107)
);

BUFx6f_ASAP7_75t_L g1108 ( 
.A(n_885),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_950),
.A2(n_957),
.B1(n_893),
.B2(n_886),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_873),
.A2(n_906),
.B(n_905),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_845),
.A2(n_904),
.B(n_931),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_914),
.Y(n_1112)
);

INVx2_ASAP7_75t_SL g1113 ( 
.A(n_943),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_SL g1114 ( 
.A1(n_893),
.A2(n_902),
.B(n_938),
.C(n_940),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_958),
.B(n_899),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_957),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_918),
.B(n_902),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_957),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_921),
.A2(n_948),
.B(n_892),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_959),
.A2(n_909),
.B(n_942),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_865),
.A2(n_937),
.B(n_940),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_947),
.A2(n_879),
.B(n_805),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_958),
.A2(n_837),
.B1(n_947),
.B2(n_828),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_947),
.B(n_802),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_828),
.B(n_832),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_897),
.A2(n_832),
.B(n_828),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_802),
.B(n_811),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_802),
.B(n_843),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_802),
.B(n_811),
.Y(n_1129)
);

NAND2x1p5_ASAP7_75t_L g1130 ( 
.A(n_803),
.B(n_807),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_802),
.B(n_811),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_897),
.A2(n_832),
.B(n_828),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_897),
.A2(n_832),
.B(n_828),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_897),
.A2(n_832),
.B(n_828),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_828),
.B(n_832),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_897),
.A2(n_832),
.B(n_828),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_828),
.B(n_832),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_828),
.A2(n_832),
.B1(n_815),
.B2(n_811),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_828),
.B(n_832),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_828),
.A2(n_832),
.B1(n_815),
.B2(n_811),
.Y(n_1140)
);

NAND2xp33_ASAP7_75t_L g1141 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1141)
);

A2O1A1Ixp33_ASAP7_75t_L g1142 ( 
.A1(n_1137),
.A2(n_1139),
.B(n_1129),
.C(n_1131),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_964),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1019),
.B(n_1127),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_971),
.A2(n_1132),
.B(n_1126),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_973),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_R g1148 ( 
.A(n_981),
.B(n_978),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_987),
.A2(n_1140),
.B1(n_1138),
.B2(n_1100),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_983),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1128),
.B(n_1011),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_1066),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_971),
.A2(n_1136),
.B(n_1134),
.Y(n_1153)
);

AOI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1014),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1041),
.A2(n_1005),
.B(n_1111),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_999),
.B(n_1013),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1023),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_1039),
.A2(n_1040),
.B(n_1001),
.C(n_1059),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1064),
.B(n_1106),
.Y(n_1159)
);

OAI22x1_ASAP7_75t_L g1160 ( 
.A1(n_1094),
.A2(n_1115),
.B1(n_1073),
.B2(n_1021),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1068),
.B(n_1006),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1030),
.B(n_980),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_966),
.A2(n_982),
.B(n_1007),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1005),
.A2(n_1032),
.B(n_1003),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_993),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1009),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_972),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1010),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1109),
.A2(n_1078),
.B(n_1120),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_SL g1170 ( 
.A1(n_1012),
.A2(n_1077),
.B(n_1107),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1050),
.B(n_1024),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_SL g1172 ( 
.A1(n_1098),
.A2(n_1006),
.B(n_986),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1031),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1066),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_965),
.A2(n_1099),
.B(n_997),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1052),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_1121),
.A2(n_1095),
.B(n_1053),
.C(n_1074),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1105),
.B(n_1113),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_974),
.A2(n_998),
.B(n_963),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_996),
.A2(n_990),
.B(n_970),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1066),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1033),
.A2(n_962),
.B(n_1025),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1110),
.A2(n_1119),
.B(n_1016),
.Y(n_1183)
);

AND2x4_ASAP7_75t_L g1184 ( 
.A(n_1068),
.B(n_1027),
.Y(n_1184)
);

BUFx2_ASAP7_75t_L g1185 ( 
.A(n_1002),
.Y(n_1185)
);

BUFx3_ASAP7_75t_L g1186 ( 
.A(n_972),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_972),
.B(n_1061),
.Y(n_1187)
);

OAI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1037),
.A2(n_1124),
.B1(n_1081),
.B2(n_1116),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_988),
.B(n_1092),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1121),
.A2(n_1076),
.B1(n_1096),
.B2(n_1086),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1090),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1123),
.B(n_985),
.Y(n_1192)
);

OAI22x1_ASAP7_75t_L g1193 ( 
.A1(n_1093),
.A2(n_1060),
.B1(n_1067),
.B2(n_969),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1112),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_1038),
.A2(n_1042),
.B1(n_989),
.B2(n_984),
.C(n_1046),
.Y(n_1195)
);

AO31x2_ASAP7_75t_L g1196 ( 
.A1(n_1091),
.A2(n_1119),
.A3(n_1049),
.B(n_1097),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1071),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1075),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1072),
.B(n_985),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1000),
.B(n_1008),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1071),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1072),
.B(n_1018),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1033),
.A2(n_1025),
.B(n_1022),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1117),
.A2(n_977),
.B(n_1036),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_1029),
.B(n_1079),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_1071),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1049),
.A2(n_992),
.A3(n_1089),
.B(n_1062),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_976),
.B(n_1048),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1036),
.A2(n_1130),
.B(n_1101),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_968),
.A2(n_1047),
.B(n_967),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1082),
.B(n_1085),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1086),
.A2(n_1130),
.B1(n_1104),
.B2(n_1029),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1043),
.A2(n_1034),
.B(n_1044),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1104),
.B(n_1102),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1103),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1114),
.A2(n_1047),
.B(n_1035),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1057),
.A2(n_1051),
.B(n_1055),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1087),
.B(n_1103),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1055),
.A2(n_1069),
.B(n_1063),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_1079),
.A2(n_1083),
.B1(n_1103),
.B2(n_1108),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_SL g1221 ( 
.A(n_1118),
.B(n_1079),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_1087),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_1020),
.Y(n_1223)
);

AO21x1_ASAP7_75t_L g1224 ( 
.A1(n_1062),
.A2(n_1063),
.B(n_1080),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1118),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1083),
.A2(n_1108),
.B1(n_1118),
.B2(n_1122),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_994),
.A2(n_1028),
.B(n_1069),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1108),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1045),
.B(n_1122),
.Y(n_1229)
);

AOI21x1_ASAP7_75t_SL g1230 ( 
.A1(n_994),
.A2(n_1080),
.B(n_1084),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_L g1231 ( 
.A(n_1054),
.B(n_1017),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_975),
.B(n_1083),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1026),
.B(n_1065),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1058),
.A2(n_1056),
.B(n_1088),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1056),
.Y(n_1235)
);

AO21x1_ASAP7_75t_L g1236 ( 
.A1(n_1070),
.A2(n_1140),
.B(n_1138),
.Y(n_1236)
);

INVx4_ASAP7_75t_L g1237 ( 
.A(n_1006),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1128),
.B(n_843),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1138),
.A2(n_1140),
.A3(n_1098),
.B(n_1133),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1246)
);

INVx5_ASAP7_75t_L g1247 ( 
.A(n_1066),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1252)
);

OAI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1001),
.A2(n_1129),
.B1(n_1131),
.B2(n_1127),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_1068),
.B(n_851),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1255)
);

OAI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_971),
.A2(n_1132),
.B(n_1126),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1138),
.B(n_1140),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1128),
.B(n_843),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_SL g1260 ( 
.A(n_981),
.B(n_808),
.Y(n_1260)
);

NOR2xp67_ASAP7_75t_L g1261 ( 
.A(n_1105),
.B(n_808),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_978),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_971),
.A2(n_1132),
.B(n_1126),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1000),
.Y(n_1265)
);

INVx1_ASAP7_75t_SL g1266 ( 
.A(n_964),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_971),
.A2(n_1132),
.B(n_1126),
.Y(n_1267)
);

NAND2xp33_ASAP7_75t_L g1268 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1268)
);

AO21x2_ASAP7_75t_L g1269 ( 
.A1(n_1126),
.A2(n_1133),
.B(n_1132),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1138),
.A2(n_1140),
.A3(n_1098),
.B(n_1133),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_964),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_964),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_SL g1274 ( 
.A(n_1066),
.B(n_1071),
.Y(n_1274)
);

O2A1O1Ixp5_ASAP7_75t_L g1275 ( 
.A1(n_1127),
.A2(n_1131),
.B(n_1129),
.C(n_1138),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_973),
.Y(n_1276)
);

AO21x2_ASAP7_75t_L g1277 ( 
.A1(n_1126),
.A2(n_1133),
.B(n_1132),
.Y(n_1277)
);

OAI22x1_ASAP7_75t_L g1278 ( 
.A1(n_1001),
.A2(n_1129),
.B1(n_1131),
.B2(n_1127),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1015),
.A2(n_1004),
.B(n_1014),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_1066),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_993),
.Y(n_1282)
);

BUFx12f_ASAP7_75t_L g1283 ( 
.A(n_964),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1284)
);

BUFx6f_ASAP7_75t_L g1285 ( 
.A(n_1066),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1125),
.A2(n_1137),
.B1(n_1139),
.B2(n_1135),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_973),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1125),
.B(n_1135),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_964),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1001),
.A2(n_1129),
.B1(n_1131),
.B2(n_1127),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1125),
.A2(n_832),
.B(n_828),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_991),
.A2(n_979),
.B(n_995),
.Y(n_1293)
);

O2A1O1Ixp5_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1257),
.B(n_1224),
.C(n_1149),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_SL g1295 ( 
.A1(n_1236),
.A2(n_1170),
.B(n_1229),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1161),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1151),
.B(n_1238),
.Y(n_1297)
);

AND2x4_ASAP7_75t_L g1298 ( 
.A(n_1222),
.B(n_1167),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1167),
.B(n_1186),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1158),
.B(n_1260),
.Y(n_1300)
);

INVx3_ASAP7_75t_L g1301 ( 
.A(n_1161),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1242),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1239),
.A2(n_1243),
.B(n_1241),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1147),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1195),
.A2(n_1200),
.B1(n_1190),
.B2(n_1160),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1255),
.A2(n_1272),
.B1(n_1284),
.B2(n_1259),
.Y(n_1307)
);

BUFx2_ASAP7_75t_L g1308 ( 
.A(n_1273),
.Y(n_1308)
);

OAI21xp33_ASAP7_75t_L g1309 ( 
.A1(n_1289),
.A2(n_1156),
.B(n_1159),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1157),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1286),
.A2(n_1144),
.B1(n_1190),
.B2(n_1142),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1275),
.A2(n_1208),
.B(n_1142),
.C(n_1177),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1185),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1177),
.A2(n_1171),
.B1(n_1257),
.B2(n_1243),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1283),
.B(n_1290),
.Y(n_1315)
);

INVxp67_ASAP7_75t_SL g1316 ( 
.A(n_1150),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1247),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1211),
.A2(n_1202),
.B1(n_1199),
.B2(n_1208),
.Y(n_1318)
);

INVx3_ASAP7_75t_SL g1319 ( 
.A(n_1262),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1228),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1275),
.A2(n_1141),
.B(n_1268),
.C(n_1279),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1258),
.B(n_1162),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1198),
.B(n_1265),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1244),
.A2(n_1252),
.B1(n_1292),
.B2(n_1249),
.Y(n_1324)
);

INVx2_ASAP7_75t_SL g1325 ( 
.A(n_1290),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1244),
.A2(n_1264),
.B(n_1292),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1249),
.A2(n_1252),
.B(n_1264),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1279),
.B(n_1253),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1247),
.B(n_1221),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1186),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1233),
.A2(n_1291),
.B1(n_1278),
.B2(n_1189),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1276),
.B(n_1287),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1233),
.A2(n_1192),
.B1(n_1231),
.B2(n_1193),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1271),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1165),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1192),
.A2(n_1188),
.B1(n_1254),
.B2(n_1178),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1228),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1218),
.B(n_1191),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1204),
.A2(n_1216),
.B(n_1280),
.Y(n_1339)
);

AOI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1183),
.A2(n_1179),
.B(n_1163),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1254),
.B(n_1168),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1179),
.A2(n_1163),
.B(n_1175),
.Y(n_1342)
);

AOI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1143),
.A2(n_1266),
.B(n_1214),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1184),
.B(n_1187),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_SL g1345 ( 
.A(n_1265),
.B(n_1261),
.Y(n_1345)
);

INVxp67_ASAP7_75t_SL g1346 ( 
.A(n_1274),
.Y(n_1346)
);

BUFx2_ASAP7_75t_L g1347 ( 
.A(n_1187),
.Y(n_1347)
);

AND2x4_ASAP7_75t_L g1348 ( 
.A(n_1184),
.B(n_1225),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_1223),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1173),
.B(n_1282),
.Y(n_1350)
);

AOI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1175),
.A2(n_1145),
.B(n_1256),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1166),
.B(n_1176),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_1205),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1176),
.A2(n_1194),
.B1(n_1227),
.B2(n_1210),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1153),
.A2(n_1263),
.B(n_1267),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1245),
.B(n_1270),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1245),
.B(n_1270),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1197),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1215),
.B(n_1226),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1172),
.A2(n_1216),
.B(n_1235),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1237),
.B(n_1247),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1152),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1152),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_1148),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1212),
.A2(n_1247),
.B1(n_1220),
.B2(n_1232),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1197),
.Y(n_1366)
);

OR2x2_ASAP7_75t_L g1367 ( 
.A(n_1245),
.B(n_1270),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1269),
.A2(n_1277),
.B(n_1219),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1237),
.B(n_1181),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1148),
.Y(n_1370)
);

OR2x6_ASAP7_75t_L g1371 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1197),
.A2(n_1285),
.B1(n_1206),
.B2(n_1281),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1197),
.Y(n_1373)
);

OAI21xp33_ASAP7_75t_L g1374 ( 
.A1(n_1154),
.A2(n_1234),
.B(n_1180),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1201),
.A2(n_1206),
.B1(n_1285),
.B2(n_1281),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1174),
.B(n_1285),
.Y(n_1376)
);

NAND3xp33_ASAP7_75t_L g1377 ( 
.A(n_1201),
.B(n_1281),
.C(n_1285),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1245),
.B(n_1270),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1196),
.B(n_1207),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1201),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1201),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1206),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1281),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1209),
.A2(n_1182),
.B1(n_1213),
.B2(n_1203),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1230),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1217),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1196),
.B(n_1207),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1207),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1155),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1146),
.B(n_1250),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1240),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1196),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1196),
.B(n_1246),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1288),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1164),
.B(n_1293),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_SL g1396 ( 
.A(n_1200),
.B(n_1156),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1236),
.A2(n_1001),
.B1(n_1040),
.B2(n_1039),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1148),
.Y(n_1398)
);

INVx3_ASAP7_75t_L g1399 ( 
.A(n_1161),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1159),
.B(n_983),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_L g1402 ( 
.A(n_1156),
.B(n_999),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1222),
.B(n_1167),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1290),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1185),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1147),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1147),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1147),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1147),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1158),
.A2(n_1127),
.B1(n_1131),
.B2(n_1129),
.Y(n_1414)
);

OAI21xp33_ASAP7_75t_L g1415 ( 
.A1(n_1158),
.A2(n_802),
.B(n_1001),
.Y(n_1415)
);

NAND2x1p5_ASAP7_75t_L g1416 ( 
.A(n_1247),
.B(n_1221),
.Y(n_1416)
);

OAI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1149),
.A2(n_1169),
.B(n_1158),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1242),
.A2(n_1248),
.B1(n_1255),
.B2(n_1251),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1247),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1147),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1147),
.Y(n_1421)
);

BUFx3_ASAP7_75t_L g1422 ( 
.A(n_1290),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1151),
.B(n_1128),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1290),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1151),
.B(n_1128),
.Y(n_1425)
);

OR2x2_ASAP7_75t_L g1426 ( 
.A(n_1159),
.B(n_983),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1169),
.A2(n_1241),
.B(n_1239),
.Y(n_1427)
);

INVx5_ASAP7_75t_L g1428 ( 
.A(n_1197),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1148),
.Y(n_1429)
);

BUFx4_ASAP7_75t_SL g1430 ( 
.A(n_1290),
.Y(n_1430)
);

INVxp67_ASAP7_75t_SL g1431 ( 
.A(n_1242),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1158),
.A2(n_1127),
.B(n_1131),
.C(n_1129),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1169),
.A2(n_1241),
.B(n_1239),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1242),
.A2(n_1248),
.B1(n_1255),
.B2(n_1251),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1290),
.Y(n_1436)
);

OR2x6_ASAP7_75t_L g1437 ( 
.A(n_1283),
.B(n_916),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1169),
.A2(n_1241),
.B(n_1239),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_L g1439 ( 
.A1(n_1169),
.A2(n_1241),
.B(n_1239),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1151),
.B(n_1128),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1169),
.A2(n_1241),
.B(n_1239),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1197),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1242),
.B(n_1248),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1242),
.A2(n_1248),
.B1(n_1255),
.B2(n_1251),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1296),
.B(n_1301),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1297),
.B(n_1322),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1305),
.B(n_1400),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1317),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1332),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1425),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1428),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1300),
.A2(n_1417),
.B1(n_1431),
.B2(n_1302),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1440),
.B(n_1402),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_SL g1455 ( 
.A(n_1422),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1397),
.A2(n_1415),
.B(n_1306),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_SL g1457 ( 
.A1(n_1300),
.A2(n_1417),
.B1(n_1311),
.B2(n_1434),
.Y(n_1457)
);

INVx4_ASAP7_75t_L g1458 ( 
.A(n_1428),
.Y(n_1458)
);

CKINVDCx6p67_ASAP7_75t_R g1459 ( 
.A(n_1319),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1308),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1428),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1396),
.B(n_1344),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1304),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1310),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1415),
.A2(n_1414),
.B1(n_1309),
.B2(n_1311),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1401),
.B(n_1426),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1296),
.B(n_1301),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1443),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1313),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1344),
.B(n_1404),
.Y(n_1470)
);

OAI21x1_ASAP7_75t_L g1471 ( 
.A1(n_1339),
.A2(n_1368),
.B(n_1360),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1443),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1340),
.A2(n_1342),
.B(n_1390),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1407),
.A2(n_1410),
.B1(n_1444),
.B2(n_1441),
.Y(n_1474)
);

INVx3_ASAP7_75t_SL g1475 ( 
.A(n_1437),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1409),
.B(n_1435),
.Y(n_1476)
);

OAI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1414),
.A2(n_1445),
.B1(n_1331),
.B2(n_1418),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1309),
.A2(n_1418),
.B1(n_1307),
.B2(n_1333),
.Y(n_1478)
);

BUFx8_ASAP7_75t_L g1479 ( 
.A(n_1370),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1334),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1347),
.Y(n_1481)
);

CKINVDCx11_ASAP7_75t_R g1482 ( 
.A(n_1315),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1307),
.A2(n_1314),
.B1(n_1331),
.B2(n_1318),
.Y(n_1483)
);

BUFx3_ASAP7_75t_L g1484 ( 
.A(n_1436),
.Y(n_1484)
);

OAI21xp33_ASAP7_75t_L g1485 ( 
.A1(n_1312),
.A2(n_1336),
.B(n_1432),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1317),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1408),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1385),
.A2(n_1316),
.B1(n_1338),
.B2(n_1323),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1419),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1314),
.A2(n_1328),
.B1(n_1324),
.B2(n_1351),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1411),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_L g1492 ( 
.A1(n_1324),
.A2(n_1295),
.B1(n_1427),
.B2(n_1442),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1343),
.B(n_1341),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1364),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1433),
.A2(n_1439),
.B1(n_1438),
.B2(n_1378),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1412),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1413),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1420),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1443),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1390),
.A2(n_1326),
.B(n_1327),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1421),
.Y(n_1501)
);

BUFx8_ASAP7_75t_L g1502 ( 
.A(n_1299),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1419),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1352),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1294),
.A2(n_1321),
.B(n_1354),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1350),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1299),
.B(n_1348),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1303),
.A2(n_1374),
.B(n_1387),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1374),
.A2(n_1379),
.B(n_1384),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1365),
.A2(n_1349),
.B1(n_1405),
.B2(n_1325),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1424),
.B(n_1320),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1367),
.A2(n_1392),
.B1(n_1357),
.B2(n_1356),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1430),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1345),
.A2(n_1388),
.B1(n_1359),
.B2(n_1393),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1315),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_1358),
.Y(n_1516)
);

BUFx2_ASAP7_75t_R g1517 ( 
.A(n_1398),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1393),
.A2(n_1399),
.B1(n_1353),
.B2(n_1315),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1329),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1320),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1337),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1395),
.A2(n_1375),
.B(n_1372),
.Y(n_1522)
);

BUFx8_ASAP7_75t_L g1523 ( 
.A(n_1348),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1399),
.B(n_1298),
.Y(n_1524)
);

OAI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1329),
.A2(n_1416),
.B1(n_1346),
.B2(n_1403),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1337),
.B(n_1366),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1362),
.A2(n_1363),
.B1(n_1403),
.B2(n_1298),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1371),
.A2(n_1437),
.B1(n_1380),
.B2(n_1381),
.Y(n_1528)
);

OAI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1437),
.A2(n_1429),
.B1(n_1330),
.B2(n_1371),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_L g1530 ( 
.A(n_1361),
.B(n_1369),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1416),
.A2(n_1371),
.B1(n_1377),
.B2(n_1369),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1382),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1358),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1376),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1358),
.Y(n_1535)
);

INVx4_ASAP7_75t_L g1536 ( 
.A(n_1361),
.Y(n_1536)
);

OAI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1373),
.A2(n_1383),
.B1(n_1391),
.B2(n_1389),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1391),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1389),
.B(n_1386),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1386),
.A2(n_1415),
.B1(n_1129),
.B2(n_1131),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1394),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_SL g1542 ( 
.A1(n_1300),
.A2(n_1001),
.B1(n_802),
.B2(n_1039),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1317),
.B(n_1419),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1297),
.B(n_1322),
.Y(n_1544)
);

INVx11_ASAP7_75t_L g1545 ( 
.A(n_1430),
.Y(n_1545)
);

CKINVDCx20_ASAP7_75t_R g1546 ( 
.A(n_1364),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1305),
.B(n_1400),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1428),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1364),
.Y(n_1549)
);

CKINVDCx20_ASAP7_75t_R g1550 ( 
.A(n_1364),
.Y(n_1550)
);

INVx1_ASAP7_75t_SL g1551 ( 
.A(n_1308),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1332),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1332),
.Y(n_1553)
);

CKINVDCx11_ASAP7_75t_R g1554 ( 
.A(n_1319),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1332),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1303),
.A2(n_1327),
.B(n_1326),
.Y(n_1556)
);

OAI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1300),
.A2(n_802),
.B1(n_1156),
.B2(n_1021),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1332),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1308),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1332),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1297),
.B(n_1322),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1332),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1415),
.A2(n_1129),
.B1(n_1131),
.B2(n_1127),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1305),
.B(n_1400),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_SL g1565 ( 
.A1(n_1300),
.A2(n_1001),
.B1(n_802),
.B2(n_1039),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1332),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1428),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1332),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1317),
.Y(n_1569)
);

OAI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1300),
.A2(n_802),
.B1(n_1156),
.B2(n_1021),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1332),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1332),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1332),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1297),
.B(n_1322),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1406),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1332),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1308),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1332),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1335),
.Y(n_1579)
);

NAND2x1p5_ASAP7_75t_L g1580 ( 
.A(n_1317),
.B(n_1419),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1355),
.B(n_1169),
.Y(n_1581)
);

CKINVDCx11_ASAP7_75t_R g1582 ( 
.A(n_1319),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1317),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_SL g1584 ( 
.A1(n_1300),
.A2(n_1001),
.B1(n_802),
.B2(n_1039),
.Y(n_1584)
);

OAI21xp5_ASAP7_75t_L g1585 ( 
.A1(n_1397),
.A2(n_1158),
.B(n_1129),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1332),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1317),
.B(n_1419),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1428),
.Y(n_1588)
);

AOI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1300),
.A2(n_1001),
.B1(n_802),
.B2(n_1039),
.Y(n_1589)
);

NAND2x1p5_ASAP7_75t_L g1590 ( 
.A(n_1317),
.B(n_1419),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_1364),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1364),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_1364),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1483),
.B(n_1457),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1538),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1483),
.B(n_1512),
.Y(n_1596)
);

BUFx3_ASAP7_75t_L g1597 ( 
.A(n_1502),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1463),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1504),
.Y(n_1599)
);

INVxp67_ASAP7_75t_L g1600 ( 
.A(n_1575),
.Y(n_1600)
);

HB1xp67_ASAP7_75t_L g1601 ( 
.A(n_1526),
.Y(n_1601)
);

AO21x2_ASAP7_75t_L g1602 ( 
.A1(n_1505),
.A2(n_1471),
.B(n_1500),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1509),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1512),
.B(n_1476),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1474),
.B(n_1448),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1539),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1509),
.Y(n_1607)
);

HB1xp67_ASAP7_75t_L g1608 ( 
.A(n_1470),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1446),
.B(n_1467),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1509),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1522),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1522),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1454),
.B(n_1466),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_SL g1614 ( 
.A(n_1517),
.B(n_1549),
.Y(n_1614)
);

BUFx4f_ASAP7_75t_SL g1615 ( 
.A(n_1459),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1450),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1464),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1490),
.B(n_1465),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1461),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1490),
.B(n_1465),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1547),
.B(n_1564),
.Y(n_1621)
);

BUFx3_ASAP7_75t_L g1622 ( 
.A(n_1502),
.Y(n_1622)
);

AO21x2_ASAP7_75t_L g1623 ( 
.A1(n_1477),
.A2(n_1473),
.B(n_1585),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_SL g1624 ( 
.A(n_1549),
.B(n_1591),
.Y(n_1624)
);

OA21x2_ASAP7_75t_L g1625 ( 
.A1(n_1492),
.A2(n_1495),
.B(n_1478),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1487),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1537),
.A2(n_1589),
.B(n_1456),
.Y(n_1627)
);

AO21x2_ASAP7_75t_L g1628 ( 
.A1(n_1485),
.A2(n_1570),
.B(n_1557),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1467),
.B(n_1541),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1491),
.Y(n_1630)
);

BUFx6f_ASAP7_75t_L g1631 ( 
.A(n_1461),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1496),
.Y(n_1632)
);

AO21x2_ASAP7_75t_L g1633 ( 
.A1(n_1497),
.A2(n_1498),
.B(n_1501),
.Y(n_1633)
);

AO21x1_ASAP7_75t_SL g1634 ( 
.A1(n_1478),
.A2(n_1495),
.B(n_1514),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1581),
.Y(n_1635)
);

AO21x1_ASAP7_75t_SL g1636 ( 
.A1(n_1514),
.A2(n_1518),
.B(n_1528),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1554),
.Y(n_1637)
);

OR2x6_ASAP7_75t_L g1638 ( 
.A(n_1581),
.B(n_1508),
.Y(n_1638)
);

OR2x6_ASAP7_75t_L g1639 ( 
.A(n_1581),
.B(n_1508),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1451),
.B(n_1447),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1502),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1540),
.A2(n_1563),
.B(n_1532),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1519),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1544),
.B(n_1561),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1574),
.B(n_1462),
.Y(n_1645)
);

BUFx2_ASAP7_75t_L g1646 ( 
.A(n_1556),
.Y(n_1646)
);

BUFx2_ASAP7_75t_L g1647 ( 
.A(n_1460),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1453),
.B(n_1552),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1553),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1555),
.B(n_1558),
.Y(n_1650)
);

OR2x6_ASAP7_75t_L g1651 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1651)
);

AO21x2_ASAP7_75t_L g1652 ( 
.A1(n_1520),
.A2(n_1521),
.B(n_1493),
.Y(n_1652)
);

INVx3_ASAP7_75t_L g1653 ( 
.A(n_1519),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1467),
.B(n_1534),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1560),
.B(n_1562),
.Y(n_1655)
);

OA21x2_ASAP7_75t_L g1656 ( 
.A1(n_1540),
.A2(n_1563),
.B(n_1518),
.Y(n_1656)
);

INVx2_ASAP7_75t_SL g1657 ( 
.A(n_1523),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1469),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1525),
.B(n_1536),
.Y(n_1659)
);

INVx6_ASAP7_75t_L g1660 ( 
.A(n_1523),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1484),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1566),
.B(n_1568),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1571),
.B(n_1572),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1480),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1573),
.A2(n_1576),
.B(n_1586),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1578),
.B(n_1579),
.Y(n_1666)
);

AO21x2_ASAP7_75t_L g1667 ( 
.A1(n_1529),
.A2(n_1524),
.B(n_1506),
.Y(n_1667)
);

BUFx6f_ASAP7_75t_L g1668 ( 
.A(n_1472),
.Y(n_1668)
);

OAI21x1_ASAP7_75t_L g1669 ( 
.A1(n_1528),
.A2(n_1527),
.B(n_1569),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1527),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1511),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1510),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1472),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1542),
.B(n_1565),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1449),
.Y(n_1675)
);

INVx4_ASAP7_75t_L g1676 ( 
.A(n_1472),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1577),
.Y(n_1677)
);

AO31x2_ASAP7_75t_L g1678 ( 
.A1(n_1584),
.A2(n_1468),
.A3(n_1458),
.B(n_1481),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1449),
.Y(n_1679)
);

BUFx3_ASAP7_75t_L g1680 ( 
.A(n_1484),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1486),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1551),
.Y(n_1682)
);

AO21x2_ASAP7_75t_L g1683 ( 
.A1(n_1507),
.A2(n_1486),
.B(n_1489),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1489),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1503),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1559),
.B(n_1530),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1523),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1503),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1503),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1475),
.B(n_1530),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1633),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1595),
.B(n_1475),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1615),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1678),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1617),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1625),
.B(n_1458),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1603),
.A2(n_1452),
.B(n_1567),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1605),
.B(n_1479),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1616),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1595),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1606),
.Y(n_1701)
);

BUFx2_ASAP7_75t_L g1702 ( 
.A(n_1678),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1606),
.B(n_1459),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1621),
.B(n_1479),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1635),
.B(n_1569),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1604),
.B(n_1516),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1601),
.B(n_1479),
.Y(n_1707)
);

AOI222xp33_ASAP7_75t_L g1708 ( 
.A1(n_1594),
.A2(n_1515),
.B1(n_1482),
.B2(n_1554),
.C1(n_1582),
.C2(n_1455),
.Y(n_1708)
);

BUFx3_ASAP7_75t_L g1709 ( 
.A(n_1661),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_SL g1710 ( 
.A1(n_1674),
.A2(n_1455),
.B1(n_1548),
.B2(n_1472),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1604),
.B(n_1535),
.Y(n_1711)
);

BUFx3_ASAP7_75t_L g1712 ( 
.A(n_1661),
.Y(n_1712)
);

INVx4_ASAP7_75t_R g1713 ( 
.A(n_1680),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1635),
.B(n_1638),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1630),
.B(n_1516),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1613),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1652),
.B(n_1583),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1652),
.B(n_1583),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1638),
.B(n_1516),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1678),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1671),
.B(n_1516),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1671),
.B(n_1515),
.Y(n_1722)
);

INVx4_ASAP7_75t_L g1723 ( 
.A(n_1660),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1649),
.B(n_1482),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1632),
.B(n_1452),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1645),
.B(n_1567),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1652),
.B(n_1513),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1665),
.B(n_1628),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1645),
.B(n_1499),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1598),
.B(n_1458),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1626),
.B(n_1468),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_L g1733 ( 
.A1(n_1594),
.A2(n_1582),
.B1(n_1533),
.B2(n_1494),
.Y(n_1733)
);

OAI22xp5_ASAP7_75t_L g1734 ( 
.A1(n_1672),
.A2(n_1550),
.B1(n_1494),
.B2(n_1592),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1611),
.B(n_1590),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1625),
.B(n_1468),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1648),
.B(n_1588),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1638),
.B(n_1588),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1612),
.B(n_1580),
.Y(n_1739)
);

NOR4xp25_ASAP7_75t_SL g1740 ( 
.A(n_1637),
.B(n_1545),
.C(n_1548),
.D(n_1588),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1678),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1648),
.B(n_1548),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1625),
.B(n_1580),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1625),
.B(n_1623),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1665),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1650),
.B(n_1548),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1623),
.B(n_1587),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1628),
.A2(n_1533),
.B1(n_1593),
.B2(n_1546),
.Y(n_1749)
);

INVx4_ASAP7_75t_L g1750 ( 
.A(n_1660),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1682),
.B(n_1546),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1638),
.B(n_1588),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1612),
.B(n_1543),
.Y(n_1753)
);

NAND3xp33_ASAP7_75t_L g1754 ( 
.A(n_1728),
.B(n_1672),
.C(n_1651),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1667),
.Y(n_1755)
);

OAI21xp5_ASAP7_75t_SL g1756 ( 
.A1(n_1708),
.A2(n_1596),
.B(n_1618),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1749),
.A2(n_1651),
.B1(n_1658),
.B2(n_1686),
.C(n_1600),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1706),
.B(n_1639),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1711),
.B(n_1639),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1710),
.A2(n_1651),
.B1(n_1596),
.B2(n_1660),
.Y(n_1760)
);

OAI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1698),
.A2(n_1651),
.B1(n_1659),
.B2(n_1620),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1736),
.B(n_1694),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1727),
.B(n_1629),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_R g1764 ( 
.A(n_1693),
.B(n_1637),
.Y(n_1764)
);

NAND3xp33_ASAP7_75t_SL g1765 ( 
.A(n_1740),
.B(n_1624),
.C(n_1614),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1733),
.A2(n_1660),
.B1(n_1618),
.B2(n_1620),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1727),
.B(n_1629),
.Y(n_1767)
);

OAI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1728),
.A2(n_1669),
.B(n_1663),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1734),
.A2(n_1687),
.B(n_1657),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1724),
.A2(n_1628),
.B1(n_1627),
.B2(n_1659),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1738),
.B(n_1659),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1700),
.B(n_1627),
.Y(n_1772)
);

OAI22xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1704),
.A2(n_1687),
.B1(n_1657),
.B2(n_1622),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1702),
.B(n_1603),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1701),
.B(n_1647),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1703),
.A2(n_1659),
.B1(n_1690),
.B2(n_1670),
.Y(n_1776)
);

NAND3xp33_ASAP7_75t_L g1777 ( 
.A(n_1692),
.B(n_1670),
.C(n_1664),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1722),
.A2(n_1690),
.B1(n_1662),
.B2(n_1677),
.C(n_1622),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1726),
.B(n_1677),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1700),
.B(n_1650),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1729),
.B(n_1644),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1716),
.B(n_1655),
.Y(n_1782)
);

NAND4xp25_ASAP7_75t_L g1783 ( 
.A(n_1731),
.B(n_1662),
.C(n_1655),
.D(n_1640),
.Y(n_1783)
);

OA21x2_ASAP7_75t_L g1784 ( 
.A1(n_1691),
.A2(n_1610),
.B(n_1607),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1695),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1744),
.B(n_1666),
.C(n_1688),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1725),
.B(n_1599),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1746),
.B(n_1666),
.C(n_1688),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1748),
.B(n_1689),
.C(n_1685),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1703),
.A2(n_1707),
.B1(n_1737),
.B2(n_1742),
.Y(n_1790)
);

NOR2xp33_ASAP7_75t_L g1791 ( 
.A(n_1747),
.B(n_1683),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1751),
.A2(n_1641),
.B1(n_1597),
.B2(n_1656),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1720),
.B(n_1607),
.Y(n_1793)
);

NAND3xp33_ASAP7_75t_L g1794 ( 
.A(n_1717),
.B(n_1689),
.C(n_1685),
.Y(n_1794)
);

NAND4xp25_ASAP7_75t_L g1795 ( 
.A(n_1721),
.B(n_1640),
.C(n_1597),
.D(n_1641),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1741),
.B(n_1610),
.Y(n_1796)
);

OAI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1696),
.A2(n_1718),
.B1(n_1717),
.B2(n_1753),
.C(n_1739),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1743),
.A2(n_1634),
.B1(n_1646),
.B2(n_1684),
.C(n_1679),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1718),
.B(n_1684),
.C(n_1681),
.Y(n_1799)
);

NAND3xp33_ASAP7_75t_L g1800 ( 
.A(n_1745),
.B(n_1691),
.C(n_1730),
.Y(n_1800)
);

OAI22xp5_ASAP7_75t_L g1801 ( 
.A1(n_1709),
.A2(n_1656),
.B1(n_1654),
.B2(n_1609),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1705),
.B(n_1643),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1729),
.B(n_1709),
.Y(n_1803)
);

OAI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1696),
.A2(n_1753),
.B1(n_1739),
.B2(n_1735),
.C(n_1712),
.Y(n_1804)
);

NAND3xp33_ASAP7_75t_L g1805 ( 
.A(n_1745),
.B(n_1681),
.C(n_1675),
.Y(n_1805)
);

AOI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1723),
.A2(n_1634),
.B1(n_1656),
.B2(n_1636),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1715),
.B(n_1642),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1719),
.B(n_1602),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1696),
.A2(n_1653),
.B1(n_1643),
.B2(n_1673),
.C(n_1676),
.Y(n_1809)
);

AND4x1_ASAP7_75t_L g1810 ( 
.A(n_1730),
.B(n_1732),
.C(n_1713),
.D(n_1679),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1784),
.Y(n_1811)
);

INVxp67_ASAP7_75t_L g1812 ( 
.A(n_1791),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1762),
.B(n_1714),
.Y(n_1813)
);

AND2x2_ASAP7_75t_SL g1814 ( 
.A(n_1770),
.B(n_1714),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1785),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1791),
.B(n_1755),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1784),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1774),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1793),
.Y(n_1819)
);

AND2x4_ASAP7_75t_L g1820 ( 
.A(n_1808),
.B(n_1771),
.Y(n_1820)
);

INVx3_ASAP7_75t_L g1821 ( 
.A(n_1771),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1796),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1771),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1800),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1786),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1758),
.B(n_1697),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1805),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1807),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1759),
.B(n_1697),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1768),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1794),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1801),
.B(n_1738),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1799),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

BUFx2_ASAP7_75t_SL g1835 ( 
.A(n_1810),
.Y(n_1835)
);

BUFx2_ASAP7_75t_L g1836 ( 
.A(n_1772),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1788),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1787),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1825),
.B(n_1797),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1815),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1817),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1815),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1815),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1820),
.B(n_1803),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1812),
.B(n_1775),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1812),
.B(n_1779),
.Y(n_1846)
);

OR2x2_ASAP7_75t_SL g1847 ( 
.A(n_1837),
.B(n_1765),
.Y(n_1847)
);

AND2x4_ASAP7_75t_SL g1848 ( 
.A(n_1821),
.B(n_1723),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1818),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1825),
.B(n_1763),
.Y(n_1850)
);

NAND2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1830),
.B(n_1738),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1763),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1817),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1816),
.B(n_1838),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1824),
.B(n_1767),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1818),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1820),
.B(n_1767),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1820),
.B(n_1802),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1818),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1817),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1824),
.B(n_1777),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1819),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1819),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1820),
.B(n_1802),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1823),
.B(n_1789),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1820),
.B(n_1738),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1816),
.B(n_1773),
.Y(n_1868)
);

NAND2x1_ASAP7_75t_L g1869 ( 
.A(n_1821),
.B(n_1713),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1823),
.B(n_1813),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1821),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1819),
.Y(n_1872)
);

INVxp67_ASAP7_75t_SL g1873 ( 
.A(n_1837),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1823),
.B(n_1752),
.Y(n_1874)
);

OAI21xp33_ASAP7_75t_SL g1875 ( 
.A1(n_1814),
.A2(n_1783),
.B(n_1795),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1838),
.B(n_1790),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1821),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1811),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1822),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1823),
.B(n_1752),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1838),
.B(n_1782),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1822),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1822),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1831),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1834),
.B(n_1754),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1834),
.B(n_1761),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1866),
.B(n_1870),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1888)
);

INVx2_ASAP7_75t_SL g1889 ( 
.A(n_1869),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1840),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1868),
.B(n_1831),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1840),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1876),
.B(n_1831),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1862),
.B(n_1824),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1862),
.B(n_1833),
.Y(n_1895)
);

AOI21xp33_ASAP7_75t_L g1896 ( 
.A1(n_1873),
.A2(n_1830),
.B(n_1814),
.Y(n_1896)
);

NAND3xp33_ASAP7_75t_L g1897 ( 
.A(n_1884),
.B(n_1830),
.C(n_1839),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1885),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1842),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1842),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1841),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1843),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1849),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1858),
.B(n_1821),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1841),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1849),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1859),
.B(n_1826),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1856),
.B(n_1850),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1886),
.B(n_1833),
.Y(n_1909)
);

INVx2_ASAP7_75t_SL g1910 ( 
.A(n_1869),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1859),
.B(n_1826),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1865),
.B(n_1826),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1865),
.B(n_1829),
.Y(n_1913)
);

INVx3_ASAP7_75t_L g1914 ( 
.A(n_1866),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1857),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1839),
.B(n_1833),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1853),
.Y(n_1917)
);

OR2x2_ASAP7_75t_L g1918 ( 
.A(n_1856),
.B(n_1827),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1857),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1850),
.B(n_1828),
.Y(n_1920)
);

AND2x4_ASAP7_75t_L g1921 ( 
.A(n_1870),
.B(n_1832),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1867),
.B(n_1829),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1852),
.B(n_1827),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1867),
.B(n_1851),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1853),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1852),
.B(n_1828),
.Y(n_1926)
);

OAI211xp5_ASAP7_75t_L g1927 ( 
.A1(n_1875),
.A2(n_1756),
.B(n_1827),
.C(n_1769),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1860),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1861),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1847),
.B(n_1846),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1860),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1861),
.Y(n_1932)
);

NOR3xp33_ASAP7_75t_L g1933 ( 
.A(n_1854),
.B(n_1778),
.C(n_1757),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1851),
.B(n_1829),
.Y(n_1934)
);

AND2x4_ASAP7_75t_L g1935 ( 
.A(n_1866),
.B(n_1832),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1851),
.B(n_1813),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1863),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1890),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1908),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1924),
.B(n_1855),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1890),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1898),
.B(n_1855),
.Y(n_1942)
);

AOI22xp5_ASAP7_75t_L g1943 ( 
.A1(n_1927),
.A2(n_1814),
.B1(n_1835),
.B2(n_1832),
.Y(n_1943)
);

INVx1_ASAP7_75t_SL g1944 ( 
.A(n_1908),
.Y(n_1944)
);

INVx2_ASAP7_75t_SL g1945 ( 
.A(n_1887),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1891),
.B(n_1828),
.Y(n_1946)
);

INVx1_ASAP7_75t_SL g1947 ( 
.A(n_1894),
.Y(n_1947)
);

AOI22xp33_ASAP7_75t_L g1948 ( 
.A1(n_1933),
.A2(n_1814),
.B1(n_1835),
.B2(n_1832),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1930),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1892),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1887),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1897),
.B(n_1835),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1924),
.B(n_1874),
.Y(n_1953)
);

NOR2x1_ASAP7_75t_L g1954 ( 
.A(n_1895),
.B(n_1877),
.Y(n_1954)
);

OAI22xp33_ASAP7_75t_L g1955 ( 
.A1(n_1896),
.A2(n_1832),
.B1(n_1760),
.B2(n_1804),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1895),
.B(n_1877),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1892),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1899),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1899),
.Y(n_1959)
);

HB1xp67_ASAP7_75t_L g1960 ( 
.A(n_1918),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1936),
.B(n_1874),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1900),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1900),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1887),
.Y(n_1964)
);

AOI22xp33_ASAP7_75t_L g1965 ( 
.A1(n_1909),
.A2(n_1832),
.B1(n_1792),
.B2(n_1806),
.Y(n_1965)
);

HB1xp67_ASAP7_75t_L g1966 ( 
.A(n_1918),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1902),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1916),
.B(n_1764),
.Y(n_1968)
);

OR2x2_ASAP7_75t_L g1969 ( 
.A(n_1894),
.B(n_1847),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1914),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1902),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1903),
.Y(n_1972)
);

HB1xp67_ASAP7_75t_L g1973 ( 
.A(n_1923),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1936),
.B(n_1880),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1903),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1906),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1906),
.Y(n_1977)
);

CKINVDCx16_ASAP7_75t_R g1978 ( 
.A(n_1935),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1949),
.B(n_1893),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1939),
.B(n_1923),
.Y(n_1980)
);

INVx1_ASAP7_75t_SL g1981 ( 
.A(n_1969),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1969),
.A2(n_1952),
.B(n_1968),
.C(n_1955),
.Y(n_1982)
);

OAI22xp33_ASAP7_75t_L g1983 ( 
.A1(n_1943),
.A2(n_1914),
.B1(n_1832),
.B2(n_1910),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1948),
.A2(n_1889),
.B1(n_1910),
.B2(n_1914),
.C(n_1920),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1944),
.B(n_1926),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1968),
.B(n_1550),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1960),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1942),
.B(n_1845),
.Y(n_1988)
);

OAI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1952),
.A2(n_1965),
.B1(n_1978),
.B2(n_1945),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1966),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1973),
.Y(n_1991)
);

NAND4xp75_ASAP7_75t_L g1992 ( 
.A(n_1954),
.B(n_1956),
.C(n_1945),
.D(n_1951),
.Y(n_1992)
);

HB1xp67_ASAP7_75t_L g1993 ( 
.A(n_1947),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1946),
.B(n_1881),
.Y(n_1994)
);

OAI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1952),
.A2(n_1766),
.B1(n_1832),
.B2(n_1889),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1950),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1970),
.B(n_1887),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_SL g1998 ( 
.A(n_1952),
.B(n_1723),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1951),
.A2(n_1935),
.B(n_1921),
.Y(n_1999)
);

NOR3xp33_ASAP7_75t_L g2000 ( 
.A(n_1970),
.B(n_1798),
.C(n_1935),
.Y(n_2000)
);

OR2x2_ASAP7_75t_L g2001 ( 
.A(n_1964),
.B(n_1907),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1964),
.B(n_1907),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1950),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1958),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1958),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1940),
.A2(n_1953),
.B1(n_1921),
.B2(n_1961),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1940),
.B(n_1888),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1981),
.B(n_1953),
.Y(n_2008)
);

NAND2x1_ASAP7_75t_SL g2009 ( 
.A(n_1993),
.B(n_1934),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_2001),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_2007),
.B(n_1961),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1993),
.Y(n_2012)
);

AOI22xp33_ASAP7_75t_L g2013 ( 
.A1(n_1989),
.A2(n_1971),
.B1(n_1967),
.B2(n_1941),
.Y(n_2013)
);

NOR2xp33_ASAP7_75t_L g2014 ( 
.A(n_1986),
.B(n_1592),
.Y(n_2014)
);

NOR2xp33_ASAP7_75t_L g2015 ( 
.A(n_1979),
.B(n_1593),
.Y(n_2015)
);

NOR2x1_ASAP7_75t_L g2016 ( 
.A(n_1992),
.B(n_1967),
.Y(n_2016)
);

OR2x2_ASAP7_75t_L g2017 ( 
.A(n_1980),
.B(n_1974),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1999),
.B(n_1974),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1996),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_2006),
.B(n_1888),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_2003),
.Y(n_2021)
);

NAND2x1_ASAP7_75t_SL g2022 ( 
.A(n_1987),
.B(n_1934),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2004),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_2000),
.B(n_1904),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2005),
.Y(n_2025)
);

OR2x2_ASAP7_75t_L g2026 ( 
.A(n_1985),
.B(n_1988),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1990),
.Y(n_2027)
);

AOI22xp33_ASAP7_75t_L g2028 ( 
.A1(n_1984),
.A2(n_1957),
.B1(n_1962),
.B2(n_1938),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1991),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_2002),
.Y(n_2030)
);

AND4x1_ASAP7_75t_L g2031 ( 
.A(n_2016),
.B(n_1998),
.C(n_1982),
.D(n_2000),
.Y(n_2031)
);

AOI221x1_ASAP7_75t_L g2032 ( 
.A1(n_2012),
.A2(n_1997),
.B1(n_1959),
.B2(n_1977),
.C(n_1972),
.Y(n_2032)
);

NOR2x1_ASAP7_75t_L g2033 ( 
.A(n_2015),
.B(n_1982),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_2013),
.A2(n_1995),
.B1(n_1983),
.B2(n_1959),
.C(n_1977),
.Y(n_2034)
);

NAND4xp25_ASAP7_75t_SL g2035 ( 
.A(n_2013),
.B(n_1994),
.C(n_1995),
.D(n_1904),
.Y(n_2035)
);

AOI221xp5_ASAP7_75t_L g2036 ( 
.A1(n_2028),
.A2(n_1976),
.B1(n_1975),
.B2(n_1963),
.C(n_1921),
.Y(n_2036)
);

AOI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_2024),
.A2(n_1848),
.B1(n_1919),
.B2(n_1915),
.Y(n_2037)
);

OAI21xp5_ASAP7_75t_SL g2038 ( 
.A1(n_2028),
.A2(n_1806),
.B(n_1911),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_2009),
.A2(n_2022),
.B(n_2008),
.Y(n_2039)
);

AOI221xp5_ASAP7_75t_L g2040 ( 
.A1(n_2027),
.A2(n_1915),
.B1(n_1931),
.B2(n_1919),
.C(n_1928),
.Y(n_2040)
);

NOR2xp33_ASAP7_75t_L g2041 ( 
.A(n_2015),
.B(n_1880),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_2026),
.B(n_1764),
.Y(n_2042)
);

NAND3xp33_ASAP7_75t_SL g2043 ( 
.A(n_2018),
.B(n_1912),
.C(n_1911),
.Y(n_2043)
);

NAND4xp25_ASAP7_75t_L g2044 ( 
.A(n_2029),
.B(n_1913),
.C(n_1912),
.D(n_1922),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_SL g2045 ( 
.A(n_2017),
.B(n_1913),
.C(n_1809),
.Y(n_2045)
);

NOR3x1_ASAP7_75t_L g2046 ( 
.A(n_2039),
.B(n_2030),
.C(n_2010),
.Y(n_2046)
);

NOR3xp33_ASAP7_75t_L g2047 ( 
.A(n_2033),
.B(n_2030),
.C(n_2010),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_SL g2048 ( 
.A(n_2031),
.B(n_2020),
.C(n_2019),
.Y(n_2048)
);

OA22x2_ASAP7_75t_L g2049 ( 
.A1(n_2038),
.A2(n_2020),
.B1(n_2023),
.B2(n_2021),
.Y(n_2049)
);

AOI211xp5_ASAP7_75t_L g2050 ( 
.A1(n_2035),
.A2(n_2025),
.B(n_2014),
.C(n_2011),
.Y(n_2050)
);

OR2x2_ASAP7_75t_L g2051 ( 
.A(n_2044),
.B(n_2011),
.Y(n_2051)
);

NOR2xp67_ASAP7_75t_L g2052 ( 
.A(n_2042),
.B(n_2014),
.Y(n_2052)
);

NOR3xp33_ASAP7_75t_L g2053 ( 
.A(n_2036),
.B(n_1905),
.C(n_1901),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2041),
.B(n_1922),
.Y(n_2054)
);

NOR3xp33_ASAP7_75t_L g2055 ( 
.A(n_2034),
.B(n_1905),
.C(n_1901),
.Y(n_2055)
);

XOR2xp5_ASAP7_75t_L g2056 ( 
.A(n_2037),
.B(n_1776),
.Y(n_2056)
);

INVxp67_ASAP7_75t_L g2057 ( 
.A(n_2032),
.Y(n_2057)
);

NOR2x1_ASAP7_75t_L g2058 ( 
.A(n_2048),
.B(n_2043),
.Y(n_2058)
);

NAND3xp33_ASAP7_75t_SL g2059 ( 
.A(n_2047),
.B(n_2057),
.C(n_2050),
.Y(n_2059)
);

NAND4xp75_ASAP7_75t_L g2060 ( 
.A(n_2046),
.B(n_2040),
.C(n_2045),
.D(n_1871),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2052),
.B(n_2051),
.C(n_2054),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_2049),
.A2(n_1925),
.B(n_1917),
.Y(n_2062)
);

XOR2x1_ASAP7_75t_L g2063 ( 
.A(n_2056),
.B(n_1917),
.Y(n_2063)
);

NAND4xp25_ASAP7_75t_L g2064 ( 
.A(n_2055),
.B(n_1750),
.C(n_1929),
.D(n_1925),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_2063),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2058),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2061),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2062),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_2060),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2059),
.Y(n_2070)
);

NOR3xp33_ASAP7_75t_L g2071 ( 
.A(n_2064),
.B(n_2053),
.C(n_1932),
.Y(n_2071)
);

NOR2x1_ASAP7_75t_L g2072 ( 
.A(n_2066),
.B(n_1937),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2069),
.B(n_1844),
.Y(n_2073)
);

XNOR2xp5_ASAP7_75t_L g2074 ( 
.A(n_2070),
.B(n_1848),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2065),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_2065),
.B(n_1929),
.Y(n_2076)
);

AND2x2_ASAP7_75t_L g2077 ( 
.A(n_2067),
.B(n_1844),
.Y(n_2077)
);

NOR3xp33_ASAP7_75t_L g2078 ( 
.A(n_2075),
.B(n_2068),
.C(n_2071),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2077),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2073),
.Y(n_2080)
);

AO22x2_ASAP7_75t_L g2081 ( 
.A1(n_2080),
.A2(n_2076),
.B1(n_2071),
.B2(n_2074),
.Y(n_2081)
);

NOR2x2_ASAP7_75t_L g2082 ( 
.A(n_2081),
.B(n_2078),
.Y(n_2082)
);

BUFx2_ASAP7_75t_L g2083 ( 
.A(n_2082),
.Y(n_2083)
);

OAI21xp33_ASAP7_75t_L g2084 ( 
.A1(n_2082),
.A2(n_2079),
.B(n_2072),
.Y(n_2084)
);

OAI22xp5_ASAP7_75t_L g2085 ( 
.A1(n_2083),
.A2(n_2076),
.B1(n_1932),
.B2(n_1937),
.Y(n_2085)
);

OAI21xp5_ASAP7_75t_L g2086 ( 
.A1(n_2084),
.A2(n_1931),
.B(n_1928),
.Y(n_2086)
);

OAI22xp5_ASAP7_75t_L g2087 ( 
.A1(n_2085),
.A2(n_1877),
.B1(n_1871),
.B2(n_1878),
.Y(n_2087)
);

OA21x2_ASAP7_75t_L g2088 ( 
.A1(n_2086),
.A2(n_1878),
.B(n_1864),
.Y(n_2088)
);

AO21x2_ASAP7_75t_L g2089 ( 
.A1(n_2087),
.A2(n_1864),
.B(n_1863),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_L g2090 ( 
.A1(n_2089),
.A2(n_2088),
.B1(n_1872),
.B2(n_1883),
.Y(n_2090)
);

OAI221xp5_ASAP7_75t_R g2091 ( 
.A1(n_2090),
.A2(n_1836),
.B1(n_1883),
.B2(n_1882),
.C(n_1879),
.Y(n_2091)
);

AOI211xp5_ASAP7_75t_L g2092 ( 
.A1(n_2091),
.A2(n_1668),
.B(n_1631),
.C(n_1619),
.Y(n_2092)
);


endmodule