module real_jpeg_24880_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_1),
.A2(n_39),
.B1(n_51),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_65),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_1),
.A2(n_65),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_65),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_2),
.A2(n_39),
.B1(n_51),
.B2(n_85),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_2),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_55),
.B1(n_56),
.B2(n_85),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_85),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_3),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_5),
.A2(n_39),
.B1(n_51),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_5),
.A2(n_55),
.B1(n_56),
.B2(n_62),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_62),
.Y(n_168)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_7),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_74),
.Y(n_88)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_56),
.C(n_58),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_8),
.A2(n_39),
.B1(n_43),
.B2(n_51),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_8),
.B(n_83),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_8),
.A2(n_43),
.B1(n_55),
.B2(n_56),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_26),
.C(n_91),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_8),
.A2(n_25),
.B(n_154),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_9),
.A2(n_26),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_14),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_14),
.A2(n_24),
.B1(n_167),
.B2(n_169),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_129),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_127),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_106),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_18),
.B(n_106),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_78),
.B2(n_79),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_52),
.B1(n_76),
.B2(n_77),
.Y(n_20)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_36),
.B2(n_37),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_25),
.A2(n_29),
.B1(n_73),
.B2(n_75),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_25),
.B(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_25),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_26),
.A2(n_30),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_27),
.B(n_43),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_30),
.B(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_33),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_42),
.C(n_46),
.Y(n_37)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_51),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_38),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_99)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_51),
.B1(n_58),
.B2(n_59),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_39),
.B(n_119),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g101 ( 
.A1(n_42),
.A2(n_43),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_43),
.B(n_89),
.Y(n_174)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_48),
.C(n_51),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_69),
.C(n_72),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_60),
.B(n_63),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g95 ( 
.A1(n_55),
.A2(n_56),
.B1(n_90),
.B2(n_91),
.Y(n_95)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_56),
.B(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_61),
.A2(n_66),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_64),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp33_ASAP7_75t_L g137 ( 
.A1(n_67),
.A2(n_138),
.B(n_139),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_70),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_72),
.Y(n_110)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_75),
.Y(n_176)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_97),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B(n_93),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_89),
.A2(n_93),
.B(n_135),
.Y(n_151)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_114),
.B1(n_116),
.B2(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B(n_102),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_117),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_108),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_117),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_113),
.B(n_115),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_115),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_120),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_125),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_143),
.B(n_191),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_140),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_131),
.B(n_140),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.C(n_136),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_185),
.B(n_190),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_164),
.B(n_184),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_158),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_158),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_151),
.C(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_153),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_162),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_172),
.B(n_183),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_170),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_168),
.A2(n_176),
.B(n_177),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_178),
.B(n_182),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_189),
.Y(n_190)
);


endmodule