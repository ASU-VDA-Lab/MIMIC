module fake_jpeg_18125_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g11 ( 
.A(n_6),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_9),
.B(n_1),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_24),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_11),
.B1(n_21),
.B2(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_29),
.Y(n_32)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_31),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_30),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_13),
.B1(n_2),
.B2(n_1),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_17),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_47),
.Y(n_68)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_45),
.A2(n_49),
.B1(n_58),
.B2(n_13),
.Y(n_70)
);

XOR2x2_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_18),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_50),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_20),
.B1(n_28),
.B2(n_27),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_27),
.C(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_18),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_37),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_66),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_70),
.A2(n_44),
.B1(n_55),
.B2(n_6),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_76),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_47),
.B1(n_58),
.B2(n_49),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_77),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_50),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_63),
.C(n_68),
.Y(n_83)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_45),
.B1(n_57),
.B2(n_46),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_80),
.A2(n_81),
.B1(n_65),
.B2(n_69),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_74),
.C(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_64),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_85),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_86),
.A2(n_77),
.B1(n_78),
.B2(n_80),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_88),
.B(n_86),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_90),
.C(n_82),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_74),
.C(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_92),
.Y(n_95)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_96),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_94),
.A2(n_95),
.B1(n_71),
.B2(n_7),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_73),
.C(n_71),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_97),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_4),
.B(n_5),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_98),
.A2(n_99),
.B(n_7),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_5),
.B(n_10),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_100),
.Y(n_103)
);


endmodule