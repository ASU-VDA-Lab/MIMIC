module real_jpeg_5045_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_0),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_0),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_0),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_0),
.B(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_0),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_0),
.B(n_360),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_0),
.B(n_38),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_1),
.Y(n_244)
);

INVx8_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_1),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g333 ( 
.A(n_1),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_2),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_2),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_2),
.B(n_161),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_2),
.B(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_3),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_3),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_3),
.Y(n_181)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_3),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_4),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_4),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_4),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_4),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_4),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_4),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_5),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_5),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_5),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_5),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_SL g268 ( 
.A(n_5),
.B(n_50),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_5),
.B(n_357),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_5),
.B(n_42),
.Y(n_397)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_6),
.Y(n_74)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_6),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_6),
.Y(n_124)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_6),
.Y(n_195)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_7),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_8),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_9),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_9),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_9),
.B(n_291),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_9),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_9),
.B(n_337),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_9),
.B(n_47),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_9),
.B(n_276),
.Y(n_382)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_10),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_10),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_10),
.Y(n_354)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_11),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_12),
.Y(n_256)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_14),
.B(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_14),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_14),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_14),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_14),
.B(n_331),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_14),
.B(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_15),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_15),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_15),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_15),
.B(n_294),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_15),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_15),
.B(n_218),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_15),
.B(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_15),
.B(n_340),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_16),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_16),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_16),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_16),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_16),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_16),
.B(n_384),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_17),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_17),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_17),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_17),
.B(n_254),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_17),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_17),
.B(n_294),
.Y(n_398)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_19),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_19),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_19),
.B(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_474),
.B(n_476),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_183),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_182),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_145),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_25),
.B(n_145),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_106),
.B2(n_144),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_75),
.C(n_87),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_45),
.C(n_58),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_29),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_30),
.B(n_37),
.C(n_41),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_33),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_34),
.Y(n_247)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_44),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_36),
.A2(n_37),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_36),
.B(n_110),
.C(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_40),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_41),
.B(n_90),
.C(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_41),
.A2(n_44),
.B1(n_95),
.B2(n_96),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_45),
.B(n_58),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.C(n_53),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_46),
.B(n_53),
.Y(n_165)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_48),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_48),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_49),
.B(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_51),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g337 ( 
.A(n_55),
.Y(n_337)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_56),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_56),
.Y(n_393)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_57),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_71),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_66),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_66),
.C(n_71),
.Y(n_116)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_65),
.Y(n_341)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_70),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_74),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_87),
.B1(n_88),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_79),
.C(n_86),
.Y(n_127)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_86),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.C(n_103),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_89),
.B(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_90),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_94),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_95),
.A2(n_96),
.B1(n_160),
.B2(n_203),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_156),
.C(n_160),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_103),
.A2(n_104),
.B1(n_179),
.B2(n_180),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_169),
.C(n_179),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_115),
.C(n_116),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_111),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_116),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_128),
.B2(n_143),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_127),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_125),
.Y(n_120)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_141),
.B2(n_142),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_140),
.Y(n_130)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_139),
.Y(n_200)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_139),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.C(n_151),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_146),
.B(n_149),
.CI(n_151),
.CON(n_470),
.SN(n_470)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_166),
.C(n_168),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_152),
.B(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_164),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_153),
.B(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_164),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_163),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_163),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_168),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_176),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_176),
.Y(n_190)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_175),
.Y(n_324)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AO21x1_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_468),
.B(n_472),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_279),
.B(n_467),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_228),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_186),
.B(n_228),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_223),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_187),
.B(n_224),
.C(n_226),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_204),
.C(n_206),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_188),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_201),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_189),
.B(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_191),
.A2(n_192),
.B1(n_201),
.B2(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_196),
.C(n_199),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_193),
.B(n_199),
.Y(n_442)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_196),
.B(n_442),
.Y(n_441)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_201),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_206),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.C(n_219),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.C(n_215),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_215),
.Y(n_240)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_219),
.Y(n_262)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.C(n_235),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_230),
.B(n_233),
.Y(n_462)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_235),
.B(n_462),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_260),
.C(n_263),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_237),
.B(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_248),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_238),
.A2(n_239),
.B1(n_433),
.B2(n_434),
.Y(n_432)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g420 ( 
.A1(n_241),
.A2(n_242),
.B(n_245),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_241),
.B(n_248),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJx2_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_252),
.C(n_257),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_410)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_256),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_256),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_257),
.B(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_258),
.B(n_353),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g455 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_263),
.Y(n_456)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_272),
.C(n_275),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_265),
.B(n_444),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.C(n_269),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_266),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_268),
.A2(n_269),
.B1(n_270),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_268),
.Y(n_423)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_272),
.B(n_275),
.Y(n_444)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx6_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_460),
.B(n_466),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_447),
.B(n_459),
.Y(n_280)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_429),
.B(n_446),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_403),
.B(n_428),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_377),
.B(n_402),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_345),
.B(n_376),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_326),
.B(n_344),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_307),
.B(n_325),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_301),
.B(n_306),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_297),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_290),
.B(n_293),
.Y(n_308)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_296),
.Y(n_357)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_309),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_317),
.B2(n_318),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_310),
.B(n_320),
.C(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_315),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_315),
.Y(n_334)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_343),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_327),
.B(n_343),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_335),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_334),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_329),
.B(n_334),
.C(n_347),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_332),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_335),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_336),
.B(n_365),
.C(n_366),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_339),
.Y(n_365)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_342),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_346),
.B(n_348),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_363),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_349),
.B(n_364),
.C(n_367),
.Y(n_401)
);

XOR2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_352),
.C(n_355),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.Y(n_351)
);

INVx4_ASAP7_75t_SL g353 ( 
.A(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_358),
.B1(n_359),
.B2(n_362),
.Y(n_355)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_356),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_362),
.Y(n_386)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g400 ( 
.A(n_368),
.B(n_373),
.C(n_374),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_373),
.B1(n_374),
.B2(n_375),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_371),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_373),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_401),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_401),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_388),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_387),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_380),
.B(n_387),
.C(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_383),
.Y(n_381)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_417),
.C(n_418),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_394),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_396),
.C(n_399),
.Y(n_406)
);

BUFx24_ASAP7_75t_SL g481 ( 
.A(n_389),
.Y(n_481)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_391),
.CI(n_392),
.CON(n_389),
.SN(n_389)
);

MAJx2_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_391),
.C(n_392),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_395),
.A2(n_396),
.B1(n_399),
.B2(n_400),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_397),
.B(n_398),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_400),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_426),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_426),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_415),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_407),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_406),
.B(n_407),
.C(n_415),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_409),
.B1(n_411),
.B2(n_412),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_438),
.C(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_413),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_420),
.C(n_425),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_420),
.A2(n_421),
.B1(n_424),
.B2(n_425),
.Y(n_419)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_421),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_430),
.B(n_445),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_445),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_436),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_435),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_435),
.C(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_433),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_436),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_437),
.B(n_441),
.C(n_443),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_448),
.B(n_457),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_448),
.B(n_457),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_449),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_464),
.C(n_465),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_463),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_461),
.B(n_463),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_470),
.B(n_471),
.Y(n_473)
);

BUFx24_ASAP7_75t_SL g482 ( 
.A(n_470),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx8_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx13_ASAP7_75t_L g478 ( 
.A(n_475),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_479),
.Y(n_476)
);

BUFx12f_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);


endmodule