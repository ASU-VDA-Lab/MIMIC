module real_jpeg_26832_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_213;
wire n_179;
wire n_167;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_274;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

INVx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_1),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_61),
.B1(n_62),
.B2(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_25),
.B1(n_29),
.B2(n_78),
.Y(n_192)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_48),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_4),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_7),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_99),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_99),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_25),
.B1(n_29),
.B2(n_99),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_8),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_8),
.A2(n_57),
.B(n_58),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_8),
.B(n_38),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_8),
.A2(n_38),
.B(n_42),
.C(n_203),
.D(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_8),
.B(n_72),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_8),
.A2(n_24),
.B(n_216),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g244 ( 
.A1(n_8),
.A2(n_59),
.B(n_71),
.C(n_155),
.D(n_245),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_8),
.B(n_59),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_65),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_10),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_38),
.B(n_43),
.C(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_25),
.B1(n_29),
.B2(n_45),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_12),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_12),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_12),
.A2(n_25),
.B1(n_29),
.B2(n_68),
.Y(n_218)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_14),
.A2(n_38),
.B1(n_39),
.B2(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_14),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_15),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_15),
.A2(n_25),
.B1(n_29),
.B2(n_40),
.Y(n_149)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_16),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_128),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_126),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_105),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_21),
.B(n_82),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_81),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_22),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_36),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_24),
.A2(n_34),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_24),
.A2(n_28),
.B1(n_33),
.B2(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_24),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_24),
.A2(n_33),
.B1(n_149),
.B2(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_24),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_24),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_27),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_25),
.B(n_44),
.Y(n_204)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_29),
.A2(n_39),
.A3(n_45),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_29),
.B(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_31),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_31),
.A2(n_223),
.B(n_231),
.Y(n_230)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_32),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_32),
.A2(n_94),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_32),
.B(n_217),
.Y(n_216)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_33),
.B(n_143),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_44),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g252 ( 
.A1(n_38),
.A2(n_58),
.A3(n_245),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_39),
.B(n_76),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_41),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_46),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_42),
.A2(n_46),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_42),
.B(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_42),
.A2(n_46),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_49),
.A2(n_96),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_49),
.B(n_171),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_49),
.A2(n_169),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_49),
.B(n_143),
.Y(n_229)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_69),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_52),
.B(n_69),
.C(n_81),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_63),
.B(n_66),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_54),
.B(n_67),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_54),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_56),
.A2(n_61),
.B(n_143),
.C(n_144),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_59),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_77),
.B1(n_79),
.B2(n_80),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_70),
.A2(n_152),
.B(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_72),
.B1(n_112),
.B2(n_113),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_71),
.A2(n_72),
.B1(n_153),
.B2(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_76),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_79),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_79),
.B(n_104),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_79),
.A2(n_102),
.B(n_177),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_88),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_87),
.A2(n_88),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_90),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_100),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_91),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_92),
.B(n_95),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_98),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_125),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_115),
.B1(n_116),
.B2(n_124),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_114),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_111),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B(n_122),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_122),
.B(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_120),
.B(n_143),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_158),
.B(n_274),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_156),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_130),
.B(n_156),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.C(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_131),
.B(n_134),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_135),
.A2(n_136),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.C(n_150),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_138),
.B1(n_150),
.B2(n_151),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_147),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_195),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_181),
.B(n_194),
.Y(n_160)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_161),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_178),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_162),
.B(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_165),
.C(n_166),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_166),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_175),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_168),
.B1(n_175),
.B2(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_172),
.B(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_179),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_184),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_189),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_185),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_188),
.B(n_189),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_190),
.B(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_191),
.B(n_193),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_192),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_272),
.C(n_273),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_267),
.B(n_271),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_256),
.B(n_266),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_240),
.B(n_255),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_219),
.B(n_239),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_201),
.B(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_205),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_206),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_212),
.C(n_214),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_213),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_215),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B(n_238),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_226),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_225),
.A2(n_232),
.B(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_237),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_241),
.B(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_246),
.C(n_249),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_248),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_258),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_259),
.B(n_262),
.C(n_263),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);


endmodule