module fake_jpeg_6051_n_165 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_165);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_165;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_29),
.B(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_36),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_38),
.Y(n_59)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_16),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_15),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_41),
.B(n_28),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_28),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_26),
.B(n_15),
.C(n_20),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_24),
.B(n_22),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_18),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_58),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_32),
.A2(n_18),
.B1(n_26),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_65),
.B1(n_22),
.B2(n_17),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_25),
.Y(n_61)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_1),
.Y(n_87)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_32),
.A2(n_20),
.B1(n_24),
.B2(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_21),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_12),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_31),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_71),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_72),
.A2(n_53),
.B(n_48),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_76),
.A2(n_80),
.B1(n_83),
.B2(n_89),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_22),
.B1(n_17),
.B2(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_58),
.A2(n_22),
.B1(n_17),
.B2(n_12),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_92),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_61),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_58),
.A2(n_17),
.B1(n_10),
.B2(n_6),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_43),
.A2(n_2),
.B(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_61),
.B1(n_56),
.B2(n_49),
.Y(n_105)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_71),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_82),
.B(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_78),
.B(n_44),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_105),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_104),
.C(n_84),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_65),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_85),
.B(n_94),
.Y(n_121)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_79),
.B(n_63),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_55),
.B1(n_49),
.B2(n_45),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_111),
.A2(n_51),
.B1(n_69),
.B2(n_82),
.Y(n_122)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_88),
.C(n_81),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_59),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_128),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_112),
.B(n_74),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_113),
.B(n_103),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_54),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_99),
.B(n_73),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_126),
.B(n_6),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_97),
.B(n_102),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_130),
.A2(n_132),
.B1(n_133),
.B2(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_111),
.B1(n_106),
.B2(n_100),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_109),
.B1(n_105),
.B2(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_138),
.B(n_126),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_139),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_138),
.B(n_119),
.Y(n_141)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_143),
.A2(n_146),
.B(n_147),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_148),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_129),
.A2(n_114),
.B(n_120),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_128),
.B(n_119),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_130),
.A2(n_123),
.B(n_95),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_122),
.Y(n_151)
);

BUFx4f_ASAP7_75t_SL g154 ( 
.A(n_142),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_127),
.B(n_54),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_133),
.B1(n_137),
.B2(n_140),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_90),
.B1(n_62),
.B2(n_57),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_152),
.B1(n_153),
.B2(n_131),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_159),
.A2(n_160),
.B1(n_67),
.B2(n_57),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_158),
.A3(n_131),
.B1(n_127),
.B2(n_90),
.C1(n_62),
.C2(n_67),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_163),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g165 ( 
.A1(n_164),
.A2(n_159),
.B1(n_160),
.B2(n_67),
.C(n_91),
.Y(n_165)
);


endmodule