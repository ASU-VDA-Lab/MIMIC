module fake_jpeg_27282_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx2_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_17),
.Y(n_50)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_15),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_58),
.B(n_16),
.C(n_23),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_28),
.B1(n_22),
.B2(n_15),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_18),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_35),
.A2(n_28),
.B1(n_22),
.B2(n_29),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_47),
.A2(n_34),
.B1(n_39),
.B2(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_29),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_28),
.B1(n_21),
.B2(n_17),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_41),
.B1(n_40),
.B2(n_16),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_21),
.B(n_20),
.C(n_19),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_40),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_32),
.B(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_72),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_71),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_36),
.B1(n_41),
.B2(n_34),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_56),
.B(n_49),
.C(n_54),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_37),
.C(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_79),
.Y(n_82)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_37),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_SL g89 ( 
.A(n_73),
.B(n_75),
.C(n_76),
.Y(n_89)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_36),
.C(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_39),
.B1(n_19),
.B2(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_45),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_86),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_85),
.B(n_92),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_63),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_80),
.B1(n_51),
.B2(n_60),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_42),
.B(n_32),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_99),
.Y(n_123)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_46),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_45),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_96),
.Y(n_121)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_100),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_32),
.B(n_23),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_73),
.C(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_24),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_98),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_105),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_83),
.B(n_69),
.C(n_78),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_116),
.C(n_96),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_95),
.B1(n_82),
.B2(n_89),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_75),
.B1(n_55),
.B2(n_48),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_92),
.B1(n_91),
.B2(n_94),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_55),
.B1(n_59),
.B2(n_39),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_115),
.B(n_122),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_95),
.C(n_86),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_62),
.B1(n_51),
.B2(n_74),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_113),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_120),
.A2(n_88),
.B(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_82),
.B(n_90),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_126),
.B(n_132),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_118),
.A2(n_121),
.B(n_112),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_138),
.Y(n_161)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_135),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_86),
.C(n_85),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_109),
.C(n_118),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_111),
.B1(n_103),
.B2(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_113),
.B1(n_97),
.B2(n_51),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_12),
.C(n_14),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_13),
.B1(n_24),
.B2(n_3),
.C(n_4),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_30),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_141),
.Y(n_148)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_93),
.B(n_97),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_121),
.B(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_146),
.B(n_147),
.Y(n_165)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_150),
.A2(n_46),
.B(n_2),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_154),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_1),
.C(n_2),
.Y(n_164)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_156),
.C(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_121),
.C(n_93),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_135),
.B1(n_137),
.B2(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_113),
.B1(n_60),
.B2(n_46),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_160),
.A2(n_126),
.B1(n_124),
.B2(n_137),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_162),
.B(n_170),
.C(n_175),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_166),
.B1(n_169),
.B2(n_160),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_3),
.Y(n_189)
);

OAI322xp33_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_125),
.A3(n_133),
.B1(n_131),
.B2(n_132),
.C1(n_142),
.C2(n_128),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_150),
.B(n_151),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_125),
.B1(n_136),
.B2(n_60),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_46),
.C(n_24),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_172),
.B(n_173),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_149),
.B(n_1),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_1),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_156),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_3),
.C(n_5),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_149),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_181),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_186),
.C(n_173),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_148),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_184),
.Y(n_193)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_174),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_145),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_188),
.Y(n_200)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_5),
.B(n_7),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_180),
.A2(n_171),
.B1(n_145),
.B2(n_144),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_191),
.B1(n_178),
.B2(n_8),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_179),
.A2(n_159),
.B1(n_144),
.B2(n_151),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_195),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_7),
.Y(n_204)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_170),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_177),
.B(n_181),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_175),
.C(n_8),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_9),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_204),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_202),
.Y(n_211)
);

NAND2xp33_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_8),
.Y(n_205)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_205),
.A2(n_9),
.B(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_200),
.B(n_193),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_207),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_196),
.A2(n_195),
.B(n_198),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_199),
.B1(n_10),
.B2(n_9),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_213),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_197),
.C(n_207),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_214),
.B(n_197),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

NAND2xp33_ASAP7_75t_R g221 ( 
.A(n_215),
.B(n_217),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_216),
.B(n_210),
.C(n_212),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_210),
.B(n_211),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_221),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_222),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_223),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);


endmodule