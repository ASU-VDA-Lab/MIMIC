module fake_netlist_1_8633_n_709 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_709);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_709;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g82 ( .A(n_20), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_31), .Y(n_83) );
NOR2xp67_ASAP7_75t_L g84 ( .A(n_9), .B(n_26), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_60), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_47), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_24), .Y(n_88) );
INVxp33_ASAP7_75t_SL g89 ( .A(n_43), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_59), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_6), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_51), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_42), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_5), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_0), .Y(n_96) );
INVxp33_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_2), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_12), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_25), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_22), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_35), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_11), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_54), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_19), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_61), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_53), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_12), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_27), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_5), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_24), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_4), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_55), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_9), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_44), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_21), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_30), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_69), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_38), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
INVxp67_ASAP7_75t_L g126 ( .A(n_15), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_58), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_56), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_50), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_83), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_83), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_106), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_106), .B(n_1), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_120), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_85), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_82), .B(n_1), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_102), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_101), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_117), .B(n_2), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_91), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_106), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_94), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_94), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_97), .B(n_114), .Y(n_154) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_114), .B(n_3), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
INVx4_ASAP7_75t_L g157 ( .A(n_101), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_118), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_82), .B(n_4), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_124), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_124), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_122), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_88), .B(n_7), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_101), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_122), .Y(n_165) );
AND2x6_ASAP7_75t_L g166 ( .A(n_125), .B(n_39), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_125), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_127), .B(n_7), .Y(n_168) );
HB1xp67_ASAP7_75t_L g169 ( .A(n_88), .Y(n_169) );
OR2x6_ASAP7_75t_L g170 ( .A(n_99), .B(n_40), .Y(n_170) );
CKINVDCx6p67_ASAP7_75t_R g171 ( .A(n_93), .Y(n_171) );
AND3x1_ASAP7_75t_L g172 ( .A(n_99), .B(n_8), .C(n_10), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_127), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_100), .B(n_10), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_101), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_154), .B(n_108), .Y(n_177) );
AND2x4_ASAP7_75t_SL g178 ( .A(n_171), .B(n_129), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_151), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_173), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_173), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_154), .B(n_100), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_132), .B(n_119), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_132), .B(n_128), .Y(n_185) );
HB1xp67_ASAP7_75t_L g186 ( .A(n_139), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_173), .Y(n_187) );
INVx5_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_133), .B(n_92), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_139), .A2(n_98), .B1(n_96), .B2(n_126), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_171), .B(n_95), .Y(n_191) );
AO22x2_ASAP7_75t_L g192 ( .A1(n_145), .A2(n_131), .B1(n_103), .B2(n_121), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_171), .B(n_131), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_175), .Y(n_194) );
INVx4_ASAP7_75t_SL g195 ( .A(n_166), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_133), .B(n_109), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_169), .B(n_115), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_166), .Y(n_199) );
INVx8_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_137), .A2(n_104), .B1(n_103), .B2(n_121), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_162), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_169), .B(n_104), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
INVx5_ASAP7_75t_L g205 ( .A(n_166), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_145), .B(n_116), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_137), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_141), .B(n_116), .Y(n_210) );
INVx4_ASAP7_75t_SL g211 ( .A(n_166), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_170), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_166), .B(n_123), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_170), .A2(n_172), .B1(n_158), .B2(n_147), .Y(n_214) );
AND2x6_ASAP7_75t_L g215 ( .A(n_170), .B(n_130), .Y(n_215) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_170), .B(n_89), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_151), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_151), .Y(n_219) );
AO22x2_ASAP7_75t_L g220 ( .A1(n_172), .A2(n_115), .B1(n_113), .B2(n_90), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_142), .B(n_107), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_151), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_143), .B(n_110), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_170), .B(n_130), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_162), .Y(n_225) );
INVx1_ASAP7_75t_SL g226 ( .A(n_136), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_143), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_144), .B(n_111), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_144), .Y(n_229) );
NAND2x1p5_ASAP7_75t_L g230 ( .A(n_155), .B(n_105), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_151), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_147), .B(n_101), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_148), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_138), .B(n_84), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_165), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_148), .A2(n_161), .B1(n_153), .B2(n_156), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_149), .B(n_112), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_149), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
INVxp67_ASAP7_75t_L g240 ( .A(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_152), .B(n_41), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_218), .Y(n_243) );
AND2x6_ASAP7_75t_L g244 ( .A(n_199), .B(n_153), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_213), .A2(n_158), .B(n_156), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_218), .B(n_160), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_198), .B(n_163), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_186), .B(n_174), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_215), .Y(n_250) );
AND2x2_ASAP7_75t_L g251 ( .A(n_186), .B(n_174), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_240), .B(n_160), .Y(n_252) );
OR2x6_ASAP7_75t_L g253 ( .A(n_200), .B(n_159), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_204), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_240), .B(n_161), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_214), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_208), .B(n_167), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g258 ( .A1(n_198), .A2(n_168), .B1(n_155), .B2(n_166), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_204), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_210), .Y(n_260) );
NOR2xp33_ASAP7_75t_R g261 ( .A(n_216), .B(n_200), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_209), .B(n_227), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_210), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_235), .Y(n_264) );
O2A1O1Ixp33_ASAP7_75t_L g265 ( .A1(n_184), .A2(n_138), .B(n_163), .C(n_159), .Y(n_265) );
BUFx8_ASAP7_75t_SL g266 ( .A(n_234), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_235), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_200), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_229), .B(n_166), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_221), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_223), .Y(n_273) );
INVx2_ASAP7_75t_SL g274 ( .A(n_206), .Y(n_274) );
BUFx8_ASAP7_75t_L g275 ( .A(n_193), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_192), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_206), .B(n_135), .Y(n_277) );
BUFx2_ASAP7_75t_L g278 ( .A(n_191), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_182), .B(n_165), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_178), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_233), .B(n_165), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_238), .B(n_162), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_192), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_203), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_182), .B(n_157), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_177), .B(n_157), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_192), .Y(n_287) );
AOI22xp5_ASAP7_75t_L g288 ( .A1(n_190), .A2(n_157), .B1(n_162), .B2(n_164), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_220), .B(n_157), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_178), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_234), .B(n_157), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_180), .Y(n_292) );
AOI22xp5_ASAP7_75t_L g293 ( .A1(n_215), .A2(n_162), .B1(n_164), .B2(n_140), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_177), .B(n_162), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_181), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_187), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_226), .B(n_11), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_194), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_196), .Y(n_299) );
INVxp67_ASAP7_75t_L g300 ( .A(n_189), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_234), .B(n_13), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_199), .Y(n_302) );
OR2x6_ASAP7_75t_L g303 ( .A(n_220), .B(n_164), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_207), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_236), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g306 ( .A1(n_215), .A2(n_164), .B1(n_140), .B2(n_150), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_230), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_188), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_228), .B(n_140), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_197), .B(n_140), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_212), .Y(n_311) );
NOR2xp33_ASAP7_75t_R g312 ( .A(n_213), .B(n_48), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_215), .Y(n_313) );
OR2x6_ASAP7_75t_L g314 ( .A(n_268), .B(n_212), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
INVx8_ASAP7_75t_L g316 ( .A(n_253), .Y(n_316) );
NOR2xp33_ASAP7_75t_SL g317 ( .A(n_290), .B(n_215), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_289), .A2(n_220), .B1(n_224), .B2(n_230), .Y(n_318) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_289), .A2(n_237), .B1(n_205), .B2(n_188), .Y(n_319) );
AO21x2_ASAP7_75t_L g320 ( .A1(n_312), .A2(n_241), .B(n_185), .Y(n_320) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_265), .A2(n_197), .B(n_237), .C(n_185), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_282), .Y(n_322) );
NAND2xp33_ASAP7_75t_L g323 ( .A(n_261), .B(n_224), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_260), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_263), .Y(n_326) );
INVxp67_ASAP7_75t_L g327 ( .A(n_249), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_251), .B(n_224), .Y(n_328) );
NAND3xp33_ASAP7_75t_L g329 ( .A(n_256), .B(n_201), .C(n_205), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_283), .A2(n_224), .B1(n_201), .B2(n_211), .Y(n_330) );
INVx5_ASAP7_75t_L g331 ( .A(n_268), .Y(n_331) );
NAND2x1p5_ASAP7_75t_L g332 ( .A(n_268), .B(n_205), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_299), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_270), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_253), .Y(n_335) );
A2O1A1Ixp33_ASAP7_75t_L g336 ( .A1(n_245), .A2(n_241), .B(n_205), .C(n_188), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_243), .B(n_224), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_253), .B(n_195), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_307), .B(n_195), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_275), .Y(n_341) );
BUFx2_ASAP7_75t_SL g342 ( .A(n_280), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_250), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_313), .Y(n_344) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_289), .A2(n_188), .B1(n_195), .B2(n_211), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_276), .B(n_211), .Y(n_346) );
BUFx3_ASAP7_75t_L g347 ( .A(n_244), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_274), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_258), .A2(n_134), .B(n_146), .C(n_150), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_300), .B(n_13), .Y(n_350) );
AOI33xp33_ASAP7_75t_L g351 ( .A1(n_284), .A2(n_134), .A3(n_146), .B1(n_150), .B2(n_202), .B3(n_225), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_271), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_250), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_246), .B(n_14), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g355 ( .A(n_247), .B(n_14), .Y(n_355) );
AOI21x1_ASAP7_75t_L g356 ( .A1(n_269), .A2(n_239), .B(n_225), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_269), .A2(n_202), .B(n_239), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_244), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g359 ( .A1(n_303), .A2(n_176), .B1(n_134), .B2(n_146), .Y(n_359) );
AO22x1_ASAP7_75t_L g360 ( .A1(n_280), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_303), .A2(n_176), .B1(n_231), .B2(n_222), .Y(n_361) );
AOI22xp33_ASAP7_75t_SL g362 ( .A1(n_301), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_287), .A2(n_176), .B1(n_21), .B2(n_22), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_250), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
BUFx10_ASAP7_75t_L g366 ( .A(n_301), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_246), .A2(n_176), .B1(n_23), .B2(n_25), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_275), .Y(n_368) );
AOI21xp5_ASAP7_75t_SL g369 ( .A1(n_303), .A2(n_176), .B(n_231), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g370 ( .A1(n_327), .A2(n_305), .B1(n_254), .B2(n_259), .C(n_279), .Y(n_370) );
INVx3_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
A2O1A1Ixp33_ASAP7_75t_L g372 ( .A1(n_321), .A2(n_277), .B(n_262), .C(n_252), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_318), .A2(n_278), .B1(n_291), .B2(n_272), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_342), .B(n_273), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_354), .B(n_252), .Y(n_376) );
BUFx8_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_354), .B(n_255), .Y(n_379) );
AO21x2_ASAP7_75t_L g380 ( .A1(n_349), .A2(n_294), .B(n_281), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
INVx4_ASAP7_75t_SL g382 ( .A(n_347), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_315), .B(n_262), .Y(n_383) );
BUFx12f_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_315), .B(n_257), .Y(n_385) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_362), .A2(n_288), .B1(n_297), .B2(n_248), .C(n_257), .Y(n_386) );
A2O1A1Ixp33_ASAP7_75t_L g387 ( .A1(n_355), .A2(n_351), .B(n_328), .C(n_329), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g388 ( .A1(n_369), .A2(n_330), .B(n_333), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_322), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_322), .Y(n_390) );
INVx3_ASAP7_75t_L g391 ( .A(n_343), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_350), .A2(n_291), .B1(n_266), .B2(n_285), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_325), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_337), .A2(n_286), .B(n_309), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_325), .A2(n_281), .B1(n_296), .B2(n_298), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_331), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_366), .B(n_348), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_333), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_331), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_331), .Y(n_400) );
BUFx3_ASAP7_75t_L g401 ( .A(n_331), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_350), .A2(n_304), .B1(n_264), .B2(n_267), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_335), .A2(n_244), .B1(n_311), .B2(n_309), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_324), .Y(n_404) );
AOI31xp67_ASAP7_75t_L g405 ( .A1(n_389), .A2(n_293), .A3(n_306), .B(n_310), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_383), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_370), .A2(n_334), .B1(n_352), .B2(n_326), .C(n_367), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_377), .A2(n_316), .B1(n_366), .B2(n_368), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_383), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_316), .B1(n_366), .B2(n_323), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_386), .A2(n_316), .B1(n_323), .B2(n_317), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_389), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_389), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_390), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_390), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_386), .A2(n_316), .B1(n_363), .B2(n_338), .Y(n_416) );
NOR2x1_ASAP7_75t_SL g417 ( .A(n_395), .B(n_338), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_338), .B1(n_369), .B2(n_314), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_377), .A2(n_368), .B1(n_341), .B2(n_347), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g422 ( .A1(n_392), .A2(n_338), .B1(n_314), .B2(n_358), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_373), .A2(n_314), .B1(n_358), .B2(n_339), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_376), .A2(n_314), .B1(n_344), .B2(n_359), .Y(n_425) );
OAI221xp5_ASAP7_75t_L g426 ( .A1(n_372), .A2(n_345), .B1(n_336), .B2(n_361), .C(n_357), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_384), .Y(n_427) );
AOI21xp33_ASAP7_75t_L g428 ( .A1(n_388), .A2(n_320), .B(n_319), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_374), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_377), .A2(n_360), .B1(n_320), .B2(n_250), .Y(n_430) );
BUFx12f_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_379), .A2(n_320), .B1(n_365), .B2(n_346), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_381), .B(n_346), .Y(n_433) );
OAI211xp5_ASAP7_75t_SL g434 ( .A1(n_402), .A2(n_365), .B(n_23), .C(n_26), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_410), .A2(n_379), .B1(n_397), .B2(n_388), .C(n_375), .Y(n_435) );
NAND4xp25_ASAP7_75t_L g436 ( .A(n_419), .B(n_404), .C(n_375), .D(n_387), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_431), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_416), .A2(n_404), .B1(n_395), .B2(n_403), .C(n_381), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_407), .A2(n_393), .B1(n_398), .B2(n_394), .C(n_380), .Y(n_439) );
BUFx3_ASAP7_75t_L g440 ( .A(n_412), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_409), .A2(n_398), .B1(n_393), .B2(n_377), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_434), .A2(n_401), .B1(n_399), .B2(n_396), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_409), .A2(n_400), .B1(n_401), .B2(n_399), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_431), .Y(n_444) );
OAI211xp5_ASAP7_75t_L g445 ( .A1(n_419), .A2(n_401), .B(n_399), .C(n_396), .Y(n_445) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_407), .A2(n_384), .B1(n_396), .B2(n_378), .C1(n_382), .C2(n_339), .Y(n_446) );
OAI21x1_ASAP7_75t_L g447 ( .A1(n_418), .A2(n_356), .B(n_391), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_423), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_406), .B(n_378), .Y(n_449) );
NOR2x1_ASAP7_75t_L g450 ( .A(n_434), .B(n_378), .Y(n_450) );
AOI221xp5_ASAP7_75t_L g451 ( .A1(n_406), .A2(n_380), .B1(n_391), .B2(n_371), .C(n_176), .Y(n_451) );
NOR4xp25_ASAP7_75t_L g452 ( .A(n_420), .B(n_391), .C(n_371), .D(n_20), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_416), .A2(n_391), .B1(n_371), .B2(n_365), .Y(n_453) );
AO21x2_ASAP7_75t_L g454 ( .A1(n_428), .A2(n_380), .B(n_346), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_423), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_423), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_420), .B(n_371), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_412), .Y(n_458) );
AOI22xp33_ASAP7_75t_SL g459 ( .A1(n_417), .A2(n_380), .B1(n_339), .B2(n_364), .Y(n_459) );
AOI33xp33_ASAP7_75t_L g460 ( .A1(n_408), .A2(n_176), .A3(n_29), .B1(n_32), .B2(n_33), .B3(n_34), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_421), .A2(n_382), .B1(n_244), .B2(n_353), .Y(n_461) );
AOI21xp5_ASAP7_75t_SL g462 ( .A1(n_417), .A2(n_382), .B(n_364), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_421), .B(n_382), .Y(n_463) );
INVx4_ASAP7_75t_L g464 ( .A(n_429), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_412), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_430), .B(n_242), .C(n_183), .Y(n_466) );
OAI211xp5_ASAP7_75t_L g467 ( .A1(n_408), .A2(n_343), .B(n_364), .C(n_353), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_415), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g469 ( .A1(n_430), .A2(n_343), .B(n_364), .C(n_353), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
NAND3xp33_ASAP7_75t_L g471 ( .A(n_452), .B(n_432), .C(n_428), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_449), .B(n_414), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_437), .Y(n_473) );
AOI33xp33_ASAP7_75t_L g474 ( .A1(n_452), .A2(n_422), .A3(n_432), .B1(n_424), .B2(n_411), .B3(n_414), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_448), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_448), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_455), .B(n_429), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_470), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g479 ( .A1(n_436), .A2(n_418), .B1(n_425), .B2(n_427), .C(n_426), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_446), .A2(n_425), .B1(n_433), .B2(n_431), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_460), .B(n_429), .C(n_415), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_455), .B(n_415), .Y(n_482) );
OAI21x1_ASAP7_75t_L g483 ( .A1(n_447), .A2(n_413), .B(n_433), .Y(n_483) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_436), .A2(n_433), .B1(n_426), .B2(n_413), .C(n_179), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_470), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_470), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_456), .Y(n_487) );
INVx2_ASAP7_75t_SL g488 ( .A(n_464), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_456), .Y(n_489) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_435), .A2(n_382), .B1(n_364), .B2(n_353), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_468), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_438), .A2(n_353), .B1(n_343), .B2(n_332), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_449), .B(n_28), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_458), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_441), .A2(n_332), .B1(n_405), .B2(n_302), .Y(n_495) );
NAND3xp33_ASAP7_75t_SL g496 ( .A(n_441), .B(n_332), .C(n_37), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_439), .A2(n_222), .B1(n_183), .B2(n_217), .C(n_242), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_458), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_450), .B(n_451), .C(n_442), .D(n_459), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_464), .B(n_36), .Y(n_500) );
XNOR2x2_ASAP7_75t_L g501 ( .A(n_466), .B(n_405), .Y(n_501) );
AOI221xp5_ASAP7_75t_L g502 ( .A1(n_457), .A2(n_222), .B1(n_183), .B2(n_242), .C(n_231), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_464), .B(n_45), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_440), .B(n_46), .Y(n_505) );
OAI211xp5_ASAP7_75t_SL g506 ( .A1(n_444), .A2(n_49), .B(n_52), .C(n_57), .Y(n_506) );
BUFx3_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_465), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_457), .B(n_62), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_440), .B(n_63), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_450), .B(n_65), .C(n_66), .D(n_67), .Y(n_511) );
AND2x4_ASAP7_75t_L g512 ( .A(n_447), .B(n_70), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_454), .B(n_71), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_444), .Y(n_514) );
INVx3_ASAP7_75t_L g515 ( .A(n_463), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_454), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_454), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_463), .B(n_72), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_466), .Y(n_519) );
AOI221xp5_ASAP7_75t_SL g520 ( .A1(n_453), .A2(n_183), .B1(n_217), .B2(n_242), .C(n_231), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_443), .B(n_73), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_475), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_478), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_475), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_476), .B(n_469), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_476), .B(n_467), .Y(n_526) );
NAND4xp25_ASAP7_75t_L g527 ( .A(n_480), .B(n_445), .C(n_461), .D(n_462), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_487), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_503), .B(n_462), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_478), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_473), .B(n_75), .C(n_76), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_487), .B(n_79), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_489), .B(n_80), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_485), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_491), .B(n_81), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_491), .Y(n_537) );
AND2x4_ASAP7_75t_SL g538 ( .A(n_488), .B(n_179), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_514), .Y(n_539) );
NOR2x1_ASAP7_75t_L g540 ( .A(n_481), .B(n_179), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_477), .B(n_179), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_477), .B(n_217), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_482), .B(n_217), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_482), .B(n_219), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_485), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_472), .B(n_219), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_488), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_486), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_486), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_508), .B(n_219), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_508), .B(n_219), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_474), .B(n_222), .Y(n_552) );
NOR3xp33_ASAP7_75t_SL g553 ( .A(n_479), .B(n_308), .C(n_302), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_515), .B(n_308), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_483), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_515), .B(n_308), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_494), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_511), .A2(n_484), .B1(n_499), .B2(n_471), .C(n_490), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g559 ( .A(n_515), .B(n_493), .Y(n_559) );
AOI31xp33_ASAP7_75t_SL g560 ( .A1(n_500), .A2(n_521), .A3(n_519), .B(n_509), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_498), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_516), .B(n_517), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_516), .B(n_517), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_513), .B(n_471), .Y(n_564) );
INVxp67_ASAP7_75t_L g565 ( .A(n_500), .Y(n_565) );
INVx3_ASAP7_75t_SL g566 ( .A(n_507), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_483), .B(n_504), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_504), .B(n_519), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_496), .A2(n_490), .B1(n_481), .B2(n_492), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_492), .B(n_495), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_512), .B(n_510), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_505), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_512), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_501), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_505), .B(n_510), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_518), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_512), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_501), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_512), .B(n_518), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_537), .Y(n_580) );
OAI21xp5_ASAP7_75t_L g581 ( .A1(n_531), .A2(n_506), .B(n_520), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_539), .B(n_497), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_576), .B(n_502), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_539), .B(n_558), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_522), .B(n_528), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_524), .B(n_528), .Y(n_586) );
INVx2_ASAP7_75t_SL g587 ( .A(n_566), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_524), .B(n_534), .Y(n_588) );
NOR3xp33_ASAP7_75t_L g589 ( .A(n_531), .B(n_558), .C(n_552), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
AOI22xp33_ASAP7_75t_SL g591 ( .A1(n_576), .A2(n_579), .B1(n_571), .B2(n_572), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_527), .B(n_564), .Y(n_592) );
AND2x4_ASAP7_75t_SL g593 ( .A(n_579), .B(n_571), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_566), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_527), .A2(n_559), .B1(n_564), .B2(n_565), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_565), .B(n_547), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_563), .B(n_566), .Y(n_597) );
AOI211x1_ASAP7_75t_L g598 ( .A1(n_529), .A2(n_573), .B(n_577), .C(n_525), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_529), .B(n_577), .Y(n_599) );
INVx3_ASAP7_75t_SL g600 ( .A(n_538), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_573), .B(n_567), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_526), .Y(n_602) );
NAND4xp25_ASAP7_75t_L g603 ( .A(n_569), .B(n_578), .C(n_574), .D(n_570), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_526), .Y(n_604) );
NAND4xp25_ASAP7_75t_SL g605 ( .A(n_540), .B(n_572), .C(n_575), .D(n_570), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_550), .Y(n_606) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_567), .B(n_568), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_568), .B(n_557), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_557), .B(n_561), .Y(n_609) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_540), .B(n_538), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_538), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_525), .A2(n_574), .B1(n_578), .B2(n_552), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_550), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_561), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_545), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_545), .B(n_549), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_574), .B(n_578), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_548), .B(n_549), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_523), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_523), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_551), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_548), .B(n_530), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_530), .B(n_535), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_530), .Y(n_624) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_553), .A2(n_536), .B1(n_533), .B2(n_532), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_580), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_600), .B(n_555), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_584), .B(n_536), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_593), .B(n_555), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_600), .B(n_555), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_593), .B(n_555), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_585), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_604), .B(n_532), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_594), .B(n_533), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_591), .A2(n_554), .B1(n_551), .B2(n_546), .Y(n_635) );
INVx6_ASAP7_75t_L g636 ( .A(n_622), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_587), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_611), .Y(n_638) );
AND2x4_ASAP7_75t_L g639 ( .A(n_601), .B(n_541), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
AO22x2_ASAP7_75t_L g641 ( .A1(n_598), .A2(n_560), .B1(n_556), .B2(n_544), .Y(n_641) );
INVx3_ASAP7_75t_L g642 ( .A(n_601), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_588), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_590), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_592), .B(n_542), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_584), .B(n_556), .C(n_543), .Y(n_646) );
NAND2x1_ASAP7_75t_L g647 ( .A(n_596), .B(n_544), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_599), .B(n_560), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_592), .B(n_595), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_603), .B(n_597), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_608), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_621), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_606), .B(n_613), .Y(n_653) );
INVxp67_ASAP7_75t_SL g654 ( .A(n_621), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_616), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_618), .Y(n_656) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_589), .A2(n_581), .B(n_596), .C(n_625), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_591), .A2(n_607), .B(n_612), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_589), .A2(n_605), .B1(n_607), .B2(n_599), .Y(n_659) );
O2A1O1Ixp33_ASAP7_75t_SL g660 ( .A1(n_617), .A2(n_610), .B(n_583), .C(n_582), .Y(n_660) );
OAI211xp5_ASAP7_75t_L g661 ( .A1(n_617), .A2(n_610), .B(n_615), .C(n_614), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_609), .B(n_620), .Y(n_662) );
AOI32xp33_ASAP7_75t_L g663 ( .A1(n_619), .A2(n_584), .A3(n_592), .B1(n_589), .B2(n_539), .Y(n_663) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_623), .A2(n_592), .B1(n_584), .B2(n_603), .C(n_598), .Y(n_664) );
AOI22x1_ASAP7_75t_L g665 ( .A1(n_624), .A2(n_600), .B1(n_594), .B2(n_431), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_602), .B(n_604), .Y(n_666) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_584), .A2(n_589), .B(n_592), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_601), .B(n_607), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_602), .B(n_604), .Y(n_669) );
OAI22xp5_ASAP7_75t_SL g670 ( .A1(n_600), .A2(n_584), .B1(n_594), .B2(n_592), .Y(n_670) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_584), .A2(n_592), .B(n_612), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_652), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_664), .B(n_650), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_670), .Y(n_674) );
AOI21x1_ASAP7_75t_SL g675 ( .A1(n_649), .A2(n_648), .B(n_668), .Y(n_675) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_659), .B(n_667), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_660), .A2(n_658), .B(n_657), .Y(n_677) );
BUFx8_ASAP7_75t_L g678 ( .A(n_637), .Y(n_678) );
AOI221x1_ASAP7_75t_L g679 ( .A1(n_671), .A2(n_650), .B1(n_641), .B2(n_626), .C(n_628), .Y(n_679) );
NAND3xp33_ASAP7_75t_SL g680 ( .A(n_663), .B(n_661), .C(n_627), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_641), .A2(n_628), .B1(n_635), .B2(n_654), .C(n_652), .Y(n_681) );
OAI211xp5_ASAP7_75t_L g682 ( .A1(n_665), .A2(n_647), .B(n_627), .C(n_630), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_666), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_669), .Y(n_684) );
OAI21xp5_ASAP7_75t_SL g685 ( .A1(n_648), .A2(n_630), .B(n_634), .Y(n_685) );
AO22x2_ASAP7_75t_L g686 ( .A1(n_637), .A2(n_648), .B1(n_638), .B2(n_668), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_686), .A2(n_642), .B1(n_665), .B2(n_641), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_683), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_674), .A2(n_646), .B1(n_645), .B2(n_639), .Y(n_689) );
OAI221xp5_ASAP7_75t_L g690 ( .A1(n_677), .A2(n_638), .B1(n_644), .B2(n_642), .C(n_640), .Y(n_690) );
OAI211xp5_ASAP7_75t_SL g691 ( .A1(n_681), .A2(n_634), .B(n_642), .C(n_653), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_673), .B(n_643), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_676), .B(n_636), .Y(n_693) );
NAND4xp25_ASAP7_75t_SL g694 ( .A(n_679), .B(n_631), .C(n_629), .D(n_651), .Y(n_694) );
AND4x1_ASAP7_75t_L g695 ( .A(n_678), .B(n_633), .C(n_655), .D(n_656), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_693), .A2(n_680), .B1(n_686), .B2(n_685), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_692), .B(n_684), .Y(n_697) );
INVxp67_ASAP7_75t_L g698 ( .A(n_690), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_688), .B(n_672), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_695), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_700), .B(n_689), .Y(n_701) );
NAND5xp2_ASAP7_75t_L g702 ( .A(n_696), .B(n_685), .C(n_682), .D(n_694), .E(n_675), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_698), .B(n_687), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_701), .B(n_697), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_703), .B(n_699), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_704), .Y(n_706) );
AOI222xp33_ASAP7_75t_SL g707 ( .A1(n_706), .A2(n_705), .B1(n_691), .B2(n_702), .C1(n_678), .C2(n_655), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_707), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_708), .A2(n_632), .B(n_662), .Y(n_709) );
endmodule