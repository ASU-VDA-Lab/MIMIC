module fake_netlist_1_12701_n_675 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_675);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_675;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_68), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_60), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_85), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_33), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_72), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_93), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_49), .Y(n_106) );
INVx1_ASAP7_75t_SL g107 ( .A(n_8), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_17), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_73), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_12), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_79), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_39), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
INVx2_ASAP7_75t_SL g116 ( .A(n_65), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_97), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_20), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_94), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_17), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_77), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_63), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_11), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_18), .B(n_35), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_45), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_16), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_58), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_37), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_62), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_87), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_43), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_53), .Y(n_138) );
INVxp67_ASAP7_75t_SL g139 ( .A(n_66), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_41), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_30), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_100), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_100), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_114), .B(n_0), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_105), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_126), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_105), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_101), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_114), .B(n_1), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_111), .A2(n_1), .B1(n_3), .B2(n_4), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_128), .B(n_3), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g156 ( .A(n_98), .B(n_23), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_128), .B(n_4), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_135), .B(n_5), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_116), .B(n_5), .Y(n_159) );
OR2x2_ASAP7_75t_L g160 ( .A(n_102), .B(n_6), .Y(n_160) );
OAI21xp33_ASAP7_75t_L g161 ( .A1(n_142), .A2(n_116), .B(n_135), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_158), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_158), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_151), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_142), .Y(n_165) );
AO21x2_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_127), .B(n_141), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_143), .B(n_137), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_144), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_143), .B(n_103), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_153), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_146), .B(n_99), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_148), .B(n_104), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_148), .B(n_99), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_149), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_149), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_155), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_151), .B(n_109), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_160), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_168), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_183), .B(n_151), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_165), .B(n_151), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_183), .B(n_157), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_165), .B(n_157), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_185), .B(n_157), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_171), .B(n_178), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_162), .B(n_145), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_185), .B(n_157), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_168), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_184), .B(n_145), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_164), .B(n_154), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_164), .A2(n_102), .B1(n_118), .B2(n_115), .Y(n_198) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_171), .B(n_178), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_167), .B(n_147), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_162), .B(n_113), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_179), .B(n_139), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_162), .B(n_124), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_180), .B(n_181), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_162), .B(n_110), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_180), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_181), .B(n_119), .Y(n_211) );
OAI22xp33_ASAP7_75t_L g212 ( .A1(n_163), .A2(n_152), .B1(n_150), .B2(n_122), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_163), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_163), .B(n_156), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_163), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_174), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_174), .A2(n_152), .B1(n_129), .B2(n_110), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_216), .B(n_170), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_216), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_193), .B(n_175), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_192), .A2(n_166), .B(n_177), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_203), .B(n_166), .Y(n_222) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_199), .B(n_115), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g224 ( .A1(n_192), .A2(n_177), .B(n_161), .Y(n_224) );
OAI22x1_ASAP7_75t_L g225 ( .A1(n_212), .A2(n_120), .B1(n_107), .B2(n_118), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_208), .A2(n_166), .B(n_161), .Y(n_226) );
OAI21xp33_ASAP7_75t_L g227 ( .A1(n_196), .A2(n_129), .B(n_108), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_215), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_208), .A2(n_166), .B(n_182), .Y(n_229) );
INVxp67_ASAP7_75t_L g230 ( .A(n_199), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_199), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_188), .A2(n_182), .B(n_176), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_188), .A2(n_176), .B(n_173), .Y(n_233) );
AOI21x1_ASAP7_75t_L g234 ( .A1(n_190), .A2(n_176), .B(n_173), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_217), .A2(n_138), .B1(n_130), .B2(n_119), .Y(n_235) );
NOR2xp67_ASAP7_75t_L g236 ( .A(n_217), .B(n_6), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_215), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_190), .A2(n_173), .B(n_172), .Y(n_238) );
AO22x1_ASAP7_75t_L g239 ( .A1(n_209), .A2(n_140), .B1(n_134), .B2(n_132), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_198), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_202), .A2(n_130), .B(n_141), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_202), .B(n_106), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_210), .B(n_125), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_187), .A2(n_108), .B(n_131), .C(n_125), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_209), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_189), .B(n_112), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_210), .A2(n_131), .B(n_138), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_226), .A2(n_194), .B(n_191), .Y(n_248) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_230), .A2(n_213), .B1(n_214), .B2(n_211), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_231), .B(n_204), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_219), .Y(n_251) );
AO31x2_ASAP7_75t_L g252 ( .A1(n_221), .A2(n_211), .A3(n_213), .B(n_205), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_222), .A2(n_205), .B(n_197), .C(n_206), .Y(n_253) );
OR2x6_ASAP7_75t_L g254 ( .A(n_223), .B(n_112), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_234), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_240), .B(n_186), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_218), .B(n_244), .C(n_220), .Y(n_257) );
BUFx10_ASAP7_75t_L g258 ( .A(n_245), .Y(n_258) );
OAI21x1_ASAP7_75t_L g259 ( .A1(n_229), .A2(n_207), .B(n_201), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_207), .B(n_201), .Y(n_260) );
NOR4xp25_ASAP7_75t_L g261 ( .A(n_227), .B(n_136), .C(n_123), .D(n_133), .Y(n_261) );
AO21x1_ASAP7_75t_L g262 ( .A1(n_224), .A2(n_136), .B(n_123), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_232), .A2(n_207), .B(n_201), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_230), .A2(n_200), .B1(n_195), .B2(n_186), .Y(n_264) );
OAI21xp33_ASAP7_75t_L g265 ( .A1(n_235), .A2(n_200), .B(n_195), .Y(n_265) );
INVx1_ASAP7_75t_SL g266 ( .A(n_223), .Y(n_266) );
A2O1A1Ixp33_ASAP7_75t_L g267 ( .A1(n_244), .A2(n_200), .B(n_195), .C(n_186), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_231), .B(n_7), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_225), .B(n_112), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_238), .A2(n_133), .B(n_169), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_231), .B(n_112), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_256), .A2(n_231), .B1(n_243), .B2(n_241), .Y(n_272) );
OA21x2_ASAP7_75t_L g273 ( .A1(n_255), .A2(n_262), .B(n_270), .Y(n_273) );
OAI22x1_ASAP7_75t_L g274 ( .A1(n_268), .A2(n_242), .B1(n_228), .B2(n_237), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g275 ( .A1(n_248), .A2(n_247), .B(n_246), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_270), .A2(n_121), .B(n_169), .Y(n_276) );
OA21x2_ASAP7_75t_L g277 ( .A1(n_248), .A2(n_121), .B(n_169), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_257), .B(n_237), .Y(n_280) );
A2O1A1Ixp33_ASAP7_75t_L g281 ( .A1(n_253), .A2(n_112), .B(n_121), .C(n_169), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_252), .B(n_239), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_254), .B(n_7), .Y(n_283) );
AOI21xp33_ASAP7_75t_SL g284 ( .A1(n_254), .A2(n_8), .B(n_9), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_260), .A2(n_169), .B(n_54), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_252), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_254), .A2(n_9), .B1(n_10), .B2(n_12), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_266), .A2(n_10), .B1(n_13), .B2(n_14), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_258), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_252), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_260), .A2(n_169), .B(n_59), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_252), .B(n_15), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_286), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_283), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_290), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_286), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_290), .B(n_249), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_286), .Y(n_298) );
AO21x2_ASAP7_75t_L g299 ( .A1(n_281), .A2(n_261), .B(n_263), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_278), .B(n_249), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_278), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
OA21x2_ASAP7_75t_L g304 ( .A1(n_285), .A2(n_267), .B(n_265), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_279), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_292), .B(n_249), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_283), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_292), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_280), .B(n_268), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_279), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_281), .A2(n_250), .B(n_269), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_282), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_283), .Y(n_314) );
INVxp67_ASAP7_75t_SL g315 ( .A(n_277), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_280), .A2(n_271), .B(n_264), .Y(n_316) );
BUFx4f_ASAP7_75t_SL g317 ( .A(n_289), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_273), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_293), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_314), .B(n_287), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_298), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_314), .A2(n_287), .B1(n_288), .B2(n_274), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_293), .B(n_273), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_293), .B(n_273), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_296), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_302), .B(n_273), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_318), .B(n_285), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_296), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_302), .B(n_273), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_296), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_314), .B(n_288), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_295), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_307), .A2(n_274), .B1(n_289), .B2(n_272), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_295), .B(n_274), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_318), .B(n_285), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_277), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_301), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_303), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g343 ( .A1(n_307), .A2(n_272), .B1(n_258), .B2(n_275), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_300), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_315), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
INVx2_ASAP7_75t_SL g347 ( .A(n_300), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_297), .B(n_277), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_303), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx1_ASAP7_75t_SL g351 ( .A(n_300), .Y(n_351) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_300), .B(n_284), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_308), .B(n_297), .Y(n_353) );
BUFx6f_ASAP7_75t_L g354 ( .A(n_304), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_294), .B(n_277), .Y(n_355) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_294), .A2(n_275), .B1(n_291), .B2(n_276), .Y(n_356) );
NAND2x1_ASAP7_75t_L g357 ( .A(n_303), .B(n_276), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_315), .B(n_291), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_310), .B(n_284), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_310), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_306), .B(n_276), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_335), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_361), .B(n_306), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_361), .B(n_306), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_361), .B(n_308), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_313), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_340), .B(n_313), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_360), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_360), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_320), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_320), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_340), .B(n_305), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_342), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_332), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_348), .B(n_305), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_328), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_352), .B(n_317), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_321), .B(n_317), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_328), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_348), .B(n_305), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_348), .B(n_305), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_342), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_324), .B(n_311), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_357), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_357), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_341), .B(n_309), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_353), .B(n_311), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_324), .B(n_311), .Y(n_391) );
AND2x4_ASAP7_75t_L g392 ( .A(n_347), .B(n_311), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_331), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_319), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_324), .B(n_316), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_319), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_325), .B(n_316), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_319), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_325), .B(n_316), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_326), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_349), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_325), .B(n_316), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_326), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_326), .B(n_316), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_327), .B(n_299), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_327), .B(n_299), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_327), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_330), .B(n_299), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_330), .B(n_299), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_330), .B(n_299), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_349), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_350), .Y(n_413) );
AND2x4_ASAP7_75t_L g414 ( .A(n_347), .B(n_312), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_334), .B(n_304), .Y(n_415) );
NAND2xp33_ASAP7_75t_R g416 ( .A(n_321), .B(n_15), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_353), .B(n_309), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_334), .B(n_304), .Y(n_418) );
INVx1_ASAP7_75t_SL g419 ( .A(n_322), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_322), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_350), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_350), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_352), .B(n_312), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_347), .B(n_312), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_334), .B(n_304), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_363), .B(n_338), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_362), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_368), .B(n_341), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_338), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_363), .B(n_365), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_364), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_368), .B(n_346), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_420), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_366), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_368), .B(n_346), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_369), .B(n_367), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_365), .B(n_344), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_365), .B(n_344), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_419), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_395), .B(n_322), .Y(n_442) );
INVx3_ASAP7_75t_SL g443 ( .A(n_379), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_369), .B(n_359), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_367), .B(n_345), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_366), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_370), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_395), .B(n_345), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_419), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_395), .B(n_351), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_417), .B(n_333), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_370), .Y(n_452) );
BUFx2_ASAP7_75t_L g453 ( .A(n_372), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_351), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_371), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_371), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_380), .B(n_352), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_364), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_398), .B(n_329), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_372), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_373), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_414), .B(n_424), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_364), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_417), .B(n_323), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_389), .B(n_336), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_373), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_398), .B(n_329), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_389), .B(n_337), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_400), .B(n_329), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_375), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_400), .B(n_329), .Y(n_471) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_423), .A2(n_337), .B(n_343), .C(n_355), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_390), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_378), .B(n_355), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_378), .B(n_381), .Y(n_475) );
NOR2xp33_ASAP7_75t_SL g476 ( .A(n_374), .B(n_339), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_376), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_381), .B(n_339), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_400), .B(n_329), .Y(n_479) );
INVx2_ASAP7_75t_SL g480 ( .A(n_376), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_374), .B(n_339), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_390), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_375), .Y(n_483) );
INVx2_ASAP7_75t_SL g484 ( .A(n_392), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_403), .B(n_339), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_382), .B(n_16), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_414), .B(n_358), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_393), .B(n_18), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_393), .B(n_339), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_374), .B(n_358), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_377), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_377), .Y(n_492) );
OR2x6_ASAP7_75t_L g493 ( .A(n_414), .B(n_358), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_403), .B(n_358), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_377), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_383), .Y(n_496) );
NAND4xp75_ASAP7_75t_L g497 ( .A(n_416), .B(n_276), .C(n_304), .D(n_356), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_383), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_383), .Y(n_499) );
AND3x1_ASAP7_75t_L g500 ( .A(n_403), .B(n_19), .C(n_21), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_384), .B(n_358), .Y(n_501) );
NOR2xp67_ASAP7_75t_L g502 ( .A(n_437), .B(n_387), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_464), .B(n_406), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_431), .B(n_406), .Y(n_504) );
OAI22xp5_ASAP7_75t_SL g505 ( .A1(n_443), .A2(n_387), .B1(n_388), .B2(n_424), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_475), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_473), .B(n_384), .Y(n_507) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_497), .B(n_387), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_431), .B(n_384), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_443), .B(n_387), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_445), .B(n_386), .Y(n_511) );
NOR4xp25_ASAP7_75t_SL g512 ( .A(n_453), .B(n_449), .C(n_460), .D(n_477), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_444), .B(n_407), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g514 ( .A1(n_486), .A2(n_411), .B1(n_407), .B2(n_409), .C1(n_410), .C2(n_405), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_451), .B(n_386), .Y(n_515) );
INVx2_ASAP7_75t_SL g516 ( .A(n_438), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_438), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_466), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_465), .B(n_407), .Y(n_519) );
INVxp33_ASAP7_75t_L g520 ( .A(n_486), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_482), .B(n_409), .Y(n_521) );
INVx2_ASAP7_75t_SL g522 ( .A(n_441), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_434), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_500), .A2(n_388), .B(n_424), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_488), .A2(n_388), .B1(n_392), .B2(n_414), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_491), .B(n_386), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_434), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_480), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_480), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_488), .A2(n_388), .B1(n_392), .B2(n_414), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_461), .Y(n_531) );
OAI21xp33_ASAP7_75t_L g532 ( .A1(n_476), .A2(n_424), .B(n_411), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_492), .B(n_391), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_468), .B(n_410), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_427), .Y(n_535) );
OR2x2_ASAP7_75t_L g536 ( .A(n_495), .B(n_391), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_430), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_457), .A2(n_410), .B1(n_411), .B2(n_391), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_462), .B(n_424), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_472), .A2(n_405), .B1(n_392), .B2(n_425), .C(n_418), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_461), .Y(n_541) );
INVxp33_ASAP7_75t_L g542 ( .A(n_442), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_448), .B(n_405), .Y(n_543) );
AOI21xp33_ASAP7_75t_R g544 ( .A1(n_474), .A2(n_394), .B(n_397), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_442), .Y(n_545) );
INVxp67_ASAP7_75t_SL g546 ( .A(n_432), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_426), .B(n_392), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_428), .B(n_19), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_432), .Y(n_549) );
INVx2_ASAP7_75t_SL g550 ( .A(n_426), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_448), .B(n_394), .Y(n_551) );
INVxp67_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_458), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_429), .B(n_415), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_429), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_496), .B(n_397), .Y(n_556) );
AOI222xp33_ASAP7_75t_L g557 ( .A1(n_433), .A2(n_404), .B1(n_422), .B2(n_421), .C1(n_399), .C2(n_401), .Y(n_557) );
INVx3_ASAP7_75t_L g558 ( .A(n_462), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_435), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_498), .B(n_399), .Y(n_560) );
NAND2xp33_ASAP7_75t_SL g561 ( .A(n_439), .B(n_401), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_439), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_499), .B(n_404), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_446), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_436), .B(n_408), .Y(n_565) );
OAI22xp5_ASAP7_75t_L g566 ( .A1(n_481), .A2(n_408), .B1(n_422), .B2(n_421), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_458), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_440), .B(n_413), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_447), .Y(n_569) );
OAI221xp5_ASAP7_75t_SL g570 ( .A1(n_493), .A2(n_425), .B1(n_418), .B2(n_415), .C(n_413), .Y(n_570) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_502), .A2(n_493), .B1(n_484), .B2(n_490), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_561), .A2(n_489), .B(n_493), .Y(n_572) );
AOI222xp33_ASAP7_75t_L g573 ( .A1(n_540), .A2(n_494), .B1(n_501), .B2(n_440), .C1(n_467), .C2(n_485), .Y(n_573) );
OAI21xp33_ASAP7_75t_SL g574 ( .A1(n_557), .A2(n_484), .B(n_493), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_555), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_527), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_516), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_557), .B(n_459), .Y(n_578) );
OAI221xp5_ASAP7_75t_L g579 ( .A1(n_524), .A2(n_455), .B1(n_452), .B2(n_456), .C(n_494), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_514), .B(n_459), .Y(n_580) );
AO22x2_ASAP7_75t_L g581 ( .A1(n_525), .A2(n_462), .B1(n_487), .B2(n_485), .Y(n_581) );
OA21x2_ASAP7_75t_L g582 ( .A1(n_524), .A2(n_510), .B(n_532), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_520), .A2(n_467), .B(n_479), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_514), .B(n_487), .C(n_501), .D(n_469), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_518), .Y(n_585) );
OAI322xp33_ASAP7_75t_L g586 ( .A1(n_548), .A2(n_469), .A3(n_471), .B1(n_479), .B2(n_454), .C1(n_450), .C2(n_483), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_507), .Y(n_587) );
AOI321xp33_ASAP7_75t_L g588 ( .A1(n_525), .A2(n_487), .A3(n_471), .B1(n_450), .B2(n_454), .C(n_425), .Y(n_588) );
OAI22xp33_ASAP7_75t_L g589 ( .A1(n_542), .A2(n_483), .B1(n_470), .B2(n_463), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_562), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_504), .B(n_470), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_503), .B(n_463), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_558), .B(n_418), .Y(n_593) );
AND2x4_ASAP7_75t_L g594 ( .A(n_539), .B(n_415), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_558), .B(n_412), .Y(n_595) );
OAI322xp33_ASAP7_75t_L g596 ( .A1(n_552), .A2(n_412), .A3(n_402), .B1(n_396), .B2(n_385), .C1(n_375), .C2(n_354), .Y(n_596) );
AOI31xp33_ASAP7_75t_L g597 ( .A1(n_508), .A2(n_412), .A3(n_402), .B(n_396), .Y(n_597) );
NOR2xp67_ASAP7_75t_L g598 ( .A(n_545), .B(n_21), .Y(n_598) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_539), .B(n_402), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_519), .B(n_396), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_506), .B(n_22), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_563), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_563), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_528), .B(n_385), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_509), .B(n_385), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_547), .B(n_354), .Y(n_606) );
OAI32xp33_ASAP7_75t_L g607 ( .A1(n_530), .A2(n_312), .A3(n_22), .B1(n_276), .B2(n_354), .Y(n_607) );
AOI211xp5_ASAP7_75t_L g608 ( .A1(n_570), .A2(n_354), .B(n_312), .C(n_26), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_535), .Y(n_609) );
INVxp33_ASAP7_75t_L g610 ( .A(n_505), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_538), .A2(n_354), .B1(n_304), .B2(n_27), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_541), .B(n_354), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_530), .A2(n_354), .B1(n_25), .B2(n_28), .Y(n_613) );
AOI321xp33_ASAP7_75t_L g614 ( .A1(n_566), .A2(n_24), .A3(n_29), .B1(n_31), .B2(n_32), .C(n_34), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
OAI21xp33_ASAP7_75t_SL g616 ( .A1(n_597), .A2(n_550), .B(n_522), .Y(n_616) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_574), .A2(n_512), .B(n_517), .C(n_529), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_574), .A2(n_566), .B1(n_534), .B2(n_521), .Y(n_618) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_608), .B(n_551), .C(n_531), .D(n_568), .Y(n_619) );
A2O1A1Ixp33_ASAP7_75t_L g620 ( .A1(n_610), .A2(n_511), .B(n_554), .C(n_515), .Y(n_620) );
NAND2xp33_ASAP7_75t_SL g621 ( .A(n_578), .B(n_512), .Y(n_621) );
HAxp5_ASAP7_75t_SL g622 ( .A(n_613), .B(n_544), .CON(n_622), .SN(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_598), .A2(n_546), .B(n_549), .Y(n_623) );
OAI211xp5_ASAP7_75t_L g624 ( .A1(n_573), .A2(n_523), .B(n_543), .C(n_565), .Y(n_624) );
AOI211xp5_ASAP7_75t_L g625 ( .A1(n_579), .A2(n_569), .B(n_564), .C(n_559), .Y(n_625) );
OAI21xp33_ASAP7_75t_SL g626 ( .A1(n_599), .A2(n_533), .B(n_536), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_602), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_603), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_588), .B(n_560), .C(n_556), .Y(n_629) );
INVxp67_ASAP7_75t_SL g630 ( .A(n_576), .Y(n_630) );
AOI322xp5_ASAP7_75t_L g631 ( .A1(n_580), .A2(n_513), .A3(n_553), .B1(n_567), .B2(n_526), .C1(n_44), .C2(n_46), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_586), .A2(n_36), .B1(n_38), .B2(n_40), .C(n_42), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g633 ( .A1(n_581), .A2(n_47), .B1(n_48), .B2(n_50), .C(n_51), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_577), .B(n_52), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_590), .B(n_56), .Y(n_635) );
OAI21xp33_ASAP7_75t_L g636 ( .A1(n_581), .A2(n_57), .B(n_61), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_583), .A2(n_64), .B1(n_67), .B2(n_69), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_583), .A2(n_70), .B1(n_71), .B2(n_74), .Y(n_638) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_608), .A2(n_75), .B(n_76), .C(n_78), .Y(n_639) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_584), .A2(n_582), .B1(n_572), .B2(n_571), .Y(n_640) );
OAI221xp5_ASAP7_75t_SL g641 ( .A1(n_601), .A2(n_81), .B1(n_82), .B2(n_83), .C(n_84), .Y(n_641) );
OAI211xp5_ASAP7_75t_SL g642 ( .A1(n_585), .A2(n_88), .B(n_90), .C(n_91), .Y(n_642) );
NOR2xp33_ASAP7_75t_SL g643 ( .A(n_596), .B(n_92), .Y(n_643) );
AOI31xp33_ASAP7_75t_L g644 ( .A1(n_575), .A2(n_95), .A3(n_96), .B(n_589), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_609), .A2(n_615), .B1(n_607), .B2(n_604), .C(n_592), .Y(n_645) );
AOI211xp5_ASAP7_75t_L g646 ( .A1(n_612), .A2(n_611), .B(n_594), .C(n_593), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_591), .Y(n_647) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_582), .A2(n_614), .B1(n_600), .B2(n_587), .C(n_595), .Y(n_648) );
AOI211xp5_ASAP7_75t_L g649 ( .A1(n_594), .A2(n_604), .B(n_606), .C(n_605), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_602), .Y(n_650) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_574), .A2(n_610), .B(n_598), .C(n_588), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g652 ( .A(n_633), .B(n_651), .C(n_636), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_640), .A2(n_621), .B1(n_648), .B2(n_645), .C(n_630), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g654 ( .A1(n_640), .A2(n_617), .B1(n_616), .B2(n_626), .C(n_620), .Y(n_654) );
OAI221xp5_ASAP7_75t_L g655 ( .A1(n_623), .A2(n_618), .B1(n_625), .B2(n_643), .C(n_619), .Y(n_655) );
AOI21xp33_ASAP7_75t_SL g656 ( .A1(n_644), .A2(n_623), .B(n_622), .Y(n_656) );
NAND3xp33_ASAP7_75t_SL g657 ( .A(n_632), .B(n_631), .C(n_639), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_650), .B(n_628), .Y(n_658) );
NOR3xp33_ASAP7_75t_L g659 ( .A(n_656), .B(n_641), .C(n_634), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_658), .Y(n_660) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_652), .B(n_642), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_653), .B(n_646), .C(n_649), .Y(n_662) );
NOR2x1_ASAP7_75t_L g663 ( .A(n_661), .B(n_655), .Y(n_663) );
INVx2_ASAP7_75t_L g664 ( .A(n_660), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_659), .B(n_654), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_663), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_667), .B(n_665), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_666), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_669), .Y(n_670) );
AOI22x1_ASAP7_75t_L g671 ( .A1(n_668), .A2(n_667), .B1(n_662), .B2(n_627), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_670), .A2(n_657), .B(n_637), .Y(n_672) );
AO21x2_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_671), .B(n_635), .Y(n_673) );
OR2x2_ASAP7_75t_L g674 ( .A(n_673), .B(n_647), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_674), .A2(n_624), .B1(n_629), .B2(n_638), .Y(n_675) );
endmodule