module fake_ariane_2628_n_792 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_792);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_792;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g159 ( 
.A(n_20),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_142),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_4),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_23),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_35),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_100),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_54),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_97),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_32),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_11),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_1),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_47),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_45),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_95),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_13),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_4),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_102),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_70),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_140),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_7),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_125),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_132),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_25),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_121),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_82),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_98),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_66),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_88),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_69),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_53),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_89),
.B(n_91),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_19),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_24),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_8),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_52),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_22),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_161),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_161),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_0),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_159),
.A2(n_0),
.B(n_2),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

AND2x4_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_3),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

AND2x4_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_3),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_5),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_163),
.B(n_21),
.Y(n_230)
);

BUFx8_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_163),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g235 ( 
.A1(n_167),
.A2(n_80),
.B(n_157),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

AOI22x1_ASAP7_75t_SL g239 ( 
.A1(n_174),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_173),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g243 ( 
.A1(n_176),
.A2(n_8),
.B(n_9),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_190),
.B(n_9),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_173),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

INVx5_ASAP7_75t_L g252 ( 
.A(n_173),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_212),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_177),
.B(n_10),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_192),
.B(n_194),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_195),
.B(n_12),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_224),
.Y(n_262)
);

AND3x2_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_165),
.C(n_197),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_247),
.B(n_169),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_224),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_198),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_179),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_232),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_211),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_214),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_247),
.B(n_160),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_247),
.B(n_162),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_219),
.B(n_213),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_237),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_232),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_232),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_188),
.B1(n_207),
.B2(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_254),
.B(n_166),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_218),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_248),
.Y(n_290)
);

BUFx6f_ASAP7_75t_SL g291 ( 
.A(n_223),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_168),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_255),
.B(n_210),
.C(n_201),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_248),
.Y(n_294)
);

AO21x2_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_200),
.B(n_196),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_248),
.Y(n_296)
);

AND2x2_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_170),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_225),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_216),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_248),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_251),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_178),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_251),
.Y(n_305)
);

AND3x2_ASAP7_75t_L g306 ( 
.A(n_244),
.B(n_13),
.C(n_14),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_250),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_289),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_244),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_277),
.B(n_250),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_287),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_254),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_297),
.B(n_246),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_275),
.B(n_246),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_297),
.B(n_221),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_261),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_281),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_238),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

NOR3x1_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_249),
.C(n_258),
.Y(n_326)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_265),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_245),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_303),
.B(n_218),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_238),
.Y(n_330)
);

NAND2xp33_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_230),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_218),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_L g333 ( 
.A(n_293),
.B(n_230),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_245),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_288),
.A2(n_223),
.B1(n_227),
.B2(n_253),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_265),
.B(n_245),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_298),
.B(n_253),
.Y(n_337)
);

AND2x4_ASAP7_75t_L g338 ( 
.A(n_263),
.B(n_227),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_270),
.B(n_256),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_270),
.B(n_256),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_280),
.B(n_231),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_280),
.B(n_220),
.C(n_243),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_256),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_291),
.B(n_231),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_L g347 ( 
.A1(n_298),
.A2(n_243),
.B1(n_220),
.B2(n_227),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_259),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_291),
.B(n_231),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_260),
.B(n_227),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_260),
.B(n_222),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_262),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_222),
.Y(n_353)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_262),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_234),
.Y(n_356)
);

OAI221xp5_ASAP7_75t_L g357 ( 
.A1(n_267),
.A2(n_243),
.B1(n_220),
.B2(n_234),
.C(n_236),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_267),
.Y(n_358)
);

NAND2xp33_ASAP7_75t_L g359 ( 
.A(n_268),
.B(n_230),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_295),
.B(n_216),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_295),
.Y(n_361)
);

BUFx6f_ASAP7_75t_SL g362 ( 
.A(n_295),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_268),
.B(n_236),
.Y(n_363)
);

NOR3xp33_ASAP7_75t_L g364 ( 
.A(n_269),
.B(n_239),
.C(n_235),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_269),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_273),
.B(n_217),
.Y(n_366)
);

NAND2xp33_ASAP7_75t_L g367 ( 
.A(n_273),
.B(n_230),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_305),
.B(n_217),
.Y(n_368)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_305),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_276),
.B(n_226),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_276),
.B(n_226),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_302),
.B(n_228),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_323),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_332),
.A2(n_243),
.B(n_220),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_329),
.A2(n_302),
.B(n_301),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_336),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_344),
.A2(n_230),
.B(n_300),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_314),
.B(n_180),
.Y(n_379)
);

O2A1O1Ixp33_ASAP7_75t_L g380 ( 
.A1(n_320),
.A2(n_228),
.B(n_233),
.C(n_296),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_308),
.A2(n_301),
.B(n_300),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_296),
.B(n_294),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_230),
.B1(n_233),
.B2(n_193),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_327),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_318),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_317),
.A2(n_294),
.B(n_290),
.Y(n_387)
);

BUFx4f_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_327),
.Y(n_389)
);

AO21x1_ASAP7_75t_L g390 ( 
.A1(n_347),
.A2(n_290),
.B(n_285),
.Y(n_390)
);

AOI21xp33_ASAP7_75t_L g391 ( 
.A1(n_319),
.A2(n_189),
.B(n_186),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_328),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_324),
.B(n_310),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_310),
.B(n_184),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_309),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_330),
.B(n_239),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_185),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_312),
.A2(n_285),
.B(n_284),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_337),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_340),
.Y(n_400)
);

O2A1O1Ixp33_ASAP7_75t_L g401 ( 
.A1(n_313),
.A2(n_284),
.B(n_283),
.C(n_16),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_335),
.B(n_14),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_312),
.B(n_230),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_315),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_251),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_316),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_331),
.A2(n_252),
.B(n_242),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_350),
.A2(n_252),
.B(n_242),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_322),
.B(n_242),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_346),
.B(n_18),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_344),
.A2(n_252),
.B(n_242),
.C(n_19),
.Y(n_411)
);

OAI21x1_ASAP7_75t_L g412 ( 
.A1(n_360),
.A2(n_26),
.B(n_27),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_338),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_334),
.A2(n_28),
.B(n_29),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_341),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_333),
.A2(n_252),
.B(n_242),
.Y(n_416)
);

O2A1O1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_342),
.A2(n_364),
.B(n_357),
.C(n_356),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_326),
.B(n_242),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_321),
.B(n_252),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_369),
.A2(n_252),
.B(n_31),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_351),
.A2(n_353),
.B(n_361),
.C(n_371),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_359),
.A2(n_30),
.B(n_33),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_338),
.B(n_34),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_327),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_367),
.A2(n_36),
.B(n_37),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_321),
.B(n_327),
.Y(n_427)
);

AOI21x1_ASAP7_75t_L g428 ( 
.A1(n_355),
.A2(n_38),
.B(n_39),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_321),
.B(n_158),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_327),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_343),
.B(n_349),
.Y(n_431)
);

AOI21x1_ASAP7_75t_L g432 ( 
.A1(n_358),
.A2(n_40),
.B(n_42),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_43),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_354),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_373),
.B(n_156),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_325),
.B(n_44),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

AOI21x1_ASAP7_75t_L g439 ( 
.A1(n_352),
.A2(n_46),
.B(n_48),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_49),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_362),
.B(n_50),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_368),
.A2(n_55),
.B(n_56),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_370),
.A2(n_372),
.B(n_58),
.Y(n_443)
);

OAI21x1_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_57),
.B(n_59),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g445 ( 
.A1(n_402),
.A2(n_60),
.B(n_63),
.C(n_64),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_411),
.A2(n_65),
.B(n_67),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_386),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_375),
.A2(n_73),
.B(n_74),
.Y(n_448)
);

NAND3xp33_ASAP7_75t_L g449 ( 
.A(n_397),
.B(n_76),
.C(n_78),
.Y(n_449)
);

NAND3xp33_ASAP7_75t_L g450 ( 
.A(n_391),
.B(n_79),
.C(n_81),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_410),
.A2(n_84),
.B(n_85),
.C(n_86),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_395),
.B(n_87),
.Y(n_452)
);

AND2x2_ASAP7_75t_SL g453 ( 
.A(n_396),
.B(n_90),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_427),
.A2(n_92),
.B(n_93),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_403),
.A2(n_94),
.B(n_99),
.Y(n_455)
);

AOI21xp33_ASAP7_75t_L g456 ( 
.A1(n_413),
.A2(n_101),
.B(n_103),
.Y(n_456)
);

AO31x2_ASAP7_75t_L g457 ( 
.A1(n_390),
.A2(n_441),
.A3(n_430),
.B(n_385),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_413),
.Y(n_458)
);

AOI21x1_ASAP7_75t_L g459 ( 
.A1(n_418),
.A2(n_104),
.B(n_106),
.Y(n_459)
);

AO31x2_ASAP7_75t_L g460 ( 
.A1(n_389),
.A2(n_107),
.A3(n_108),
.B(n_110),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_378),
.A2(n_111),
.B(n_112),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_395),
.A2(n_113),
.B(n_114),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_417),
.A2(n_115),
.B(n_116),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_393),
.B(n_117),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_415),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_425),
.B(n_119),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_379),
.B(n_120),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_383),
.B(n_122),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_424),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_412),
.A2(n_123),
.B(n_126),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_394),
.A2(n_128),
.B(n_129),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_434),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_381),
.A2(n_130),
.B(n_131),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_399),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

OAI21x1_ASAP7_75t_L g478 ( 
.A1(n_382),
.A2(n_133),
.B(n_135),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_407),
.A2(n_136),
.B(n_138),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_398),
.A2(n_139),
.B(n_143),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_392),
.B(n_144),
.Y(n_481)
);

AOI21x1_ASAP7_75t_L g482 ( 
.A1(n_416),
.A2(n_145),
.B(n_146),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_147),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_438),
.A2(n_423),
.B1(n_431),
.B2(n_406),
.Y(n_484)
);

O2A1O1Ixp5_ASAP7_75t_L g485 ( 
.A1(n_387),
.A2(n_148),
.B(n_150),
.C(n_151),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_376),
.A2(n_152),
.B(n_153),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_443),
.A2(n_154),
.B(n_401),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_437),
.A2(n_436),
.B(n_433),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_388),
.B(n_435),
.Y(n_489)
);

OAI21x1_ASAP7_75t_L g490 ( 
.A1(n_421),
.A2(n_439),
.B(n_420),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_438),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_380),
.A2(n_422),
.B(n_426),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_384),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_409),
.A2(n_419),
.B(n_405),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_442),
.A2(n_429),
.B(n_404),
.Y(n_495)
);

AOI21xp33_ASAP7_75t_L g496 ( 
.A1(n_414),
.A2(n_406),
.B(n_408),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_428),
.A2(n_432),
.B(n_440),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_440),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_440),
.A2(n_378),
.B(n_375),
.Y(n_499)
);

A2O1A1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_440),
.A2(n_402),
.B(n_386),
.C(n_397),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_374),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_411),
.A2(n_375),
.B(n_417),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_489),
.B(n_477),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_466),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_498),
.Y(n_505)
);

OAI21x1_ASAP7_75t_SL g506 ( 
.A1(n_464),
.A2(n_446),
.B(n_467),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_453),
.B(n_471),
.Y(n_507)
);

AO21x2_ASAP7_75t_L g508 ( 
.A1(n_497),
.A2(n_494),
.B(n_502),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_474),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_468),
.A2(n_502),
.B(n_464),
.Y(n_510)
);

OAI21x1_ASAP7_75t_L g511 ( 
.A1(n_499),
.A2(n_497),
.B(n_490),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_444),
.A2(n_461),
.B(n_488),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_471),
.Y(n_513)
);

INVx3_ASAP7_75t_SL g514 ( 
.A(n_452),
.Y(n_514)
);

NAND2x1p5_ASAP7_75t_L g515 ( 
.A(n_491),
.B(n_469),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_495),
.A2(n_500),
.B(n_470),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_495),
.A2(n_448),
.B(n_487),
.Y(n_518)
);

AO21x2_ASAP7_75t_L g519 ( 
.A1(n_448),
.A2(n_487),
.B(n_496),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_501),
.B(n_462),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_484),
.B(n_476),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_447),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g524 ( 
.A(n_481),
.Y(n_524)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_446),
.A2(n_465),
.B(n_492),
.Y(n_525)
);

OA21x2_ASAP7_75t_L g526 ( 
.A1(n_492),
.A2(n_472),
.B(n_478),
.Y(n_526)
);

AO21x2_ASAP7_75t_L g527 ( 
.A1(n_449),
.A2(n_475),
.B(n_482),
.Y(n_527)
);

INVxp33_ASAP7_75t_L g528 ( 
.A(n_493),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_483),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_479),
.A2(n_486),
.B(n_455),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g531 ( 
.A(n_447),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_457),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_456),
.Y(n_533)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_473),
.B(n_480),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_454),
.B(n_463),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_457),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_450),
.A2(n_460),
.B(n_451),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_445),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_460),
.A2(n_468),
.B(n_467),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_460),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_498),
.Y(n_542)
);

OAI21x1_ASAP7_75t_L g543 ( 
.A1(n_499),
.A2(n_497),
.B(n_490),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_499),
.A2(n_497),
.B(n_490),
.Y(n_544)
);

AO21x2_ASAP7_75t_L g545 ( 
.A1(n_497),
.A2(n_390),
.B(n_494),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_453),
.B(n_297),
.Y(n_546)
);

OAI21x1_ASAP7_75t_SL g547 ( 
.A1(n_464),
.A2(n_446),
.B(n_467),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_476),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_468),
.A2(n_467),
.B(n_502),
.Y(n_549)
);

OAI21x1_ASAP7_75t_SL g550 ( 
.A1(n_464),
.A2(n_446),
.B(n_467),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_499),
.A2(n_497),
.B(n_490),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_504),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_522),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_521),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_513),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_546),
.A2(n_531),
.B1(n_523),
.B2(n_507),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_539),
.A2(n_510),
.B1(n_525),
.B2(n_507),
.Y(n_558)
);

AO21x1_ASAP7_75t_SL g559 ( 
.A1(n_506),
.A2(n_547),
.B(n_550),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_505),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_503),
.B(n_505),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_533),
.A2(n_522),
.B1(n_524),
.B2(n_528),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_505),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_535),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_503),
.Y(n_565)
);

INVx1_ASAP7_75t_SL g566 ( 
.A(n_548),
.Y(n_566)
);

OA21x2_ASAP7_75t_L g567 ( 
.A1(n_516),
.A2(n_511),
.B(n_551),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_503),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_552),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_515),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_515),
.B(n_532),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_509),
.Y(n_573)
);

INVx6_ASAP7_75t_L g574 ( 
.A(n_505),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_509),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_542),
.Y(n_577)
);

AO21x2_ASAP7_75t_L g578 ( 
.A1(n_540),
.A2(n_549),
.B(n_519),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_537),
.B(n_508),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_542),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_509),
.B(n_533),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_537),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_542),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_529),
.Y(n_587)
);

OAI21xp33_ASAP7_75t_SL g588 ( 
.A1(n_538),
.A2(n_529),
.B(n_518),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_514),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_514),
.Y(n_590)
);

AO21x1_ASAP7_75t_SL g591 ( 
.A1(n_518),
.A2(n_519),
.B(n_536),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_508),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_536),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_511),
.A2(n_551),
.B(n_544),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_554),
.B(n_545),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_566),
.B(n_565),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_565),
.B(n_545),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_572),
.B(n_541),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_561),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_553),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_584),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_582),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_544),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_560),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_562),
.B(n_541),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_557),
.B(n_538),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_589),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_574),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_592),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_564),
.B(n_517),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_581),
.A2(n_527),
.B1(n_517),
.B2(n_526),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_590),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_568),
.B(n_543),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

OAI21xp33_ASAP7_75t_SL g616 ( 
.A1(n_558),
.A2(n_543),
.B(n_512),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_574),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_560),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_593),
.A2(n_526),
.B1(n_534),
.B2(n_517),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_556),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_574),
.A2(n_526),
.B1(n_534),
.B2(n_527),
.Y(n_622)
);

INVx3_ASAP7_75t_SL g623 ( 
.A(n_575),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_560),
.Y(n_624)
);

INVx2_ASAP7_75t_SL g625 ( 
.A(n_574),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_570),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_570),
.B(n_512),
.Y(n_627)
);

INVx2_ASAP7_75t_SL g628 ( 
.A(n_560),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g629 ( 
.A(n_588),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_585),
.Y(n_630)
);

OR2x2_ASAP7_75t_L g631 ( 
.A(n_571),
.B(n_534),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_567),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_576),
.A2(n_530),
.B1(n_580),
.B2(n_575),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_591),
.B(n_559),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_567),
.B(n_530),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_579),
.Y(n_636)
);

AO21x2_ASAP7_75t_L g637 ( 
.A1(n_578),
.A2(n_594),
.B(n_586),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_621),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_623),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_600),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_573),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_597),
.B(n_591),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_618),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_629),
.A2(n_577),
.B1(n_560),
.B2(n_563),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_621),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_626),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_597),
.B(n_567),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_626),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_611),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_595),
.B(n_573),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_623),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_610),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_595),
.B(n_578),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_603),
.B(n_578),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_629),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_608),
.B(n_579),
.Y(n_657)
);

INVx5_ASAP7_75t_SL g658 ( 
.A(n_605),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_603),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_633),
.B(n_563),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_636),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_610),
.B(n_594),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_623),
.B(n_601),
.Y(n_663)
);

BUFx2_ASAP7_75t_L g664 ( 
.A(n_634),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_614),
.B(n_559),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_615),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_614),
.B(n_579),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_605),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_615),
.Y(n_669)
);

NOR2x1p5_ASAP7_75t_L g670 ( 
.A(n_599),
.B(n_583),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_652),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_656),
.B(n_604),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_656),
.B(n_604),
.Y(n_673)
);

AND2x4_ASAP7_75t_SL g674 ( 
.A(n_668),
.B(n_605),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_647),
.B(n_637),
.Y(n_675)
);

NOR2x1p5_ASAP7_75t_L g676 ( 
.A(n_639),
.B(n_607),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_652),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_647),
.B(n_637),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_640),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_654),
.B(n_667),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_654),
.B(n_637),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_669),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_653),
.B(n_617),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_657),
.B(n_616),
.C(n_612),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_650),
.B(n_630),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_667),
.B(n_627),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_661),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_661),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_659),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_642),
.B(n_627),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_649),
.B(n_617),
.Y(n_692)
);

AND3x1_ASAP7_75t_L g693 ( 
.A(n_663),
.B(n_634),
.C(n_624),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_655),
.B(n_631),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g695 ( 
.A1(n_651),
.A2(n_664),
.B(n_602),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_641),
.B(n_619),
.Y(n_696)
);

AND2x2_ASAP7_75t_SL g697 ( 
.A(n_664),
.B(n_598),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_642),
.B(n_665),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_638),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_669),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_638),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_666),
.Y(n_702)
);

NAND2x1_ASAP7_75t_L g703 ( 
.A(n_668),
.B(n_624),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_693),
.B(n_639),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_671),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_677),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_690),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_683),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_675),
.B(n_678),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_680),
.B(n_655),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_682),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_682),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_680),
.B(n_662),
.Y(n_713)
);

NOR2x1_ASAP7_75t_L g714 ( 
.A(n_695),
.B(n_670),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_700),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_699),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_701),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_676),
.B(n_665),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_702),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_679),
.Y(n_720)
);

OR2x2_ASAP7_75t_L g721 ( 
.A(n_672),
.B(n_662),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_697),
.B(n_668),
.Y(n_722)
);

AND2x4_ASAP7_75t_SL g723 ( 
.A(n_688),
.B(n_668),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_686),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_672),
.B(n_666),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_675),
.B(n_632),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_705),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_711),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_SL g729 ( 
.A(n_714),
.B(n_697),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_723),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_724),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_706),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_716),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_714),
.B(n_703),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_710),
.B(n_709),
.Y(n_735)
);

OAI32xp33_ASAP7_75t_L g736 ( 
.A1(n_709),
.A2(n_673),
.A3(n_685),
.B1(n_696),
.B2(n_698),
.Y(n_736)
);

OR2x6_ASAP7_75t_L g737 ( 
.A(n_704),
.B(n_660),
.Y(n_737)
);

O2A1O1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_736),
.A2(n_720),
.B(n_708),
.C(n_684),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_727),
.B(n_726),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_732),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_728),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_733),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_SL g743 ( 
.A1(n_734),
.A2(n_704),
.B(n_718),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_729),
.A2(n_737),
.B1(n_735),
.B2(n_734),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_740),
.B(n_731),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_742),
.B(n_707),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_739),
.Y(n_747)
);

NAND2x1_ASAP7_75t_L g748 ( 
.A(n_743),
.B(n_737),
.Y(n_748)
);

OA22x2_ASAP7_75t_SL g749 ( 
.A1(n_744),
.A2(n_729),
.B1(n_719),
.B2(n_717),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_741),
.A2(n_737),
.B1(n_681),
.B2(n_678),
.Y(n_750)
);

AOI221xp5_ASAP7_75t_L g751 ( 
.A1(n_738),
.A2(n_726),
.B1(n_681),
.B2(n_616),
.C(n_692),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_747),
.B(n_689),
.Y(n_752)
);

OA22x2_ASAP7_75t_L g753 ( 
.A1(n_748),
.A2(n_718),
.B1(n_730),
.B2(n_722),
.Y(n_753)
);

NAND5xp2_ASAP7_75t_L g754 ( 
.A(n_751),
.B(n_745),
.C(n_746),
.D(n_749),
.E(n_750),
.Y(n_754)
);

NOR2x1_ASAP7_75t_L g755 ( 
.A(n_745),
.B(n_730),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_755),
.B(n_725),
.C(n_673),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_752),
.Y(n_757)
);

NOR2x1_ASAP7_75t_L g758 ( 
.A(n_754),
.B(n_698),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_757),
.Y(n_759)
);

NOR2x1_ASAP7_75t_L g760 ( 
.A(n_758),
.B(n_753),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_756),
.B(n_713),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_758),
.B(n_721),
.C(n_622),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_759),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_760),
.B(n_761),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_762),
.B(n_668),
.C(n_644),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_760),
.A2(n_660),
.B1(n_606),
.B2(n_694),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_759),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_763),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_764),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_691),
.Y(n_770)
);

XOR2x2_ASAP7_75t_L g771 ( 
.A(n_766),
.B(n_609),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_765),
.B(n_723),
.Y(n_772)
);

NAND4xp75_ASAP7_75t_L g773 ( 
.A(n_764),
.B(n_625),
.C(n_609),
.D(n_628),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_R g774 ( 
.A(n_768),
.B(n_772),
.Y(n_774)
);

OAI22x1_ASAP7_75t_L g775 ( 
.A1(n_769),
.A2(n_625),
.B1(n_628),
.B2(n_624),
.Y(n_775)
);

OAI22x1_ASAP7_75t_SL g776 ( 
.A1(n_773),
.A2(n_583),
.B1(n_624),
.B2(n_632),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_770),
.B(n_674),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_771),
.B(n_691),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_775),
.A2(n_777),
.B(n_776),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_774),
.A2(n_674),
.B1(n_620),
.B2(n_715),
.Y(n_780)
);

INVxp67_ASAP7_75t_SL g781 ( 
.A(n_778),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_775),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_777),
.A2(n_694),
.B1(n_658),
.B2(n_687),
.Y(n_783)
);

AOI21xp33_ASAP7_75t_L g784 ( 
.A1(n_781),
.A2(n_712),
.B(n_648),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_780),
.A2(n_687),
.B1(n_658),
.B2(n_619),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_782),
.A2(n_658),
.B1(n_635),
.B2(n_631),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_785),
.A2(n_779),
.B1(n_783),
.B2(n_563),
.Y(n_787)
);

OA21x2_ASAP7_75t_L g788 ( 
.A1(n_784),
.A2(n_646),
.B(n_645),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_788),
.B(n_786),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_789),
.B(n_787),
.Y(n_790)
);

NAND2x2_ASAP7_75t_L g791 ( 
.A(n_790),
.B(n_619),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_791),
.A2(n_563),
.B1(n_577),
.B2(n_583),
.Y(n_792)
);


endmodule