module fake_jpeg_23054_n_334 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_42),
.Y(n_49)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_22),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_44),
.A2(n_24),
.B1(n_31),
.B2(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_24),
.B1(n_31),
.B2(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_54),
.A2(n_59),
.B1(n_63),
.B2(n_21),
.Y(n_91)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_20),
.B1(n_32),
.B2(n_28),
.Y(n_59)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_17),
.B1(n_33),
.B2(n_27),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_65),
.Y(n_114)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_22),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_67),
.B(n_69),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

NOR2xp67_ASAP7_75t_R g72 ( 
.A(n_63),
.B(n_36),
.Y(n_72)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_72),
.B(n_33),
.C(n_27),
.Y(n_110)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_79),
.B1(n_82),
.B2(n_88),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_22),
.B1(n_26),
.B2(n_17),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_33),
.B1(n_27),
.B2(n_44),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_27),
.B1(n_33),
.B2(n_48),
.Y(n_103)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_85),
.B(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_61),
.A2(n_26),
.B1(n_25),
.B2(n_21),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_25),
.B(n_30),
.Y(n_123)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_41),
.B1(n_26),
.B2(n_33),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_48),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_93),
.B(n_47),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_91),
.B(n_69),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_66),
.C(n_83),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_101),
.B1(n_109),
.B2(n_113),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_41),
.B1(n_55),
.B2(n_37),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_102),
.A2(n_103),
.B1(n_107),
.B2(n_119),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_82),
.A2(n_45),
.B1(n_36),
.B2(n_40),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_81),
.B1(n_79),
.B2(n_65),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_123),
.B(n_99),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_75),
.A2(n_33),
.B1(n_20),
.B2(n_28),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_115),
.B1(n_93),
.B2(n_84),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_112),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_47),
.B1(n_30),
.B2(n_21),
.Y(n_113)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_77),
.B(n_47),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_30),
.B1(n_25),
.B2(n_32),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_74),
.B1(n_16),
.B2(n_23),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_127),
.B(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_142),
.B1(n_147),
.B2(n_149),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_131),
.A2(n_137),
.B(n_141),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_133),
.A2(n_151),
.B1(n_152),
.B2(n_96),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_97),
.B(n_106),
.Y(n_135)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_94),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_35),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_100),
.A2(n_68),
.B(n_90),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_100),
.A2(n_16),
.B1(n_23),
.B2(n_38),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_143),
.Y(n_170)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_94),
.B(n_29),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g146 ( 
.A(n_106),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_146),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_115),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_95),
.A2(n_38),
.B1(n_35),
.B2(n_42),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_101),
.A2(n_38),
.B1(n_35),
.B2(n_42),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_132),
.A2(n_102),
.B1(n_115),
.B2(n_103),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_153),
.A2(n_185),
.B1(n_183),
.B2(n_136),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_141),
.A2(n_122),
.B(n_108),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_154),
.A2(n_156),
.B(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_155),
.A2(n_160),
.B1(n_161),
.B2(n_168),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_108),
.B(n_119),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_120),
.B(n_121),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_118),
.C(n_96),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_164),
.C(n_171),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_151),
.A2(n_118),
.B1(n_105),
.B2(n_116),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_116),
.B1(n_35),
.B2(n_38),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_177),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_16),
.B(n_23),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_167),
.A2(n_182),
.B(n_2),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_133),
.A2(n_42),
.B1(n_34),
.B2(n_19),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_29),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_29),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_178),
.C(n_181),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g175 ( 
.A1(n_126),
.A2(n_29),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_175),
.B(n_0),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_127),
.B(n_71),
.C(n_34),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_19),
.C(n_1),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_129),
.A2(n_0),
.B(n_1),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_184),
.B(n_5),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_136),
.A2(n_142),
.B1(n_124),
.B2(n_125),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_173),
.Y(n_189)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_191),
.B1(n_205),
.B2(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_152),
.B1(n_137),
.B2(n_144),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_161),
.Y(n_192)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_193),
.A2(n_204),
.B1(n_216),
.B2(n_174),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_195),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_180),
.A2(n_143),
.B(n_4),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_196),
.A2(n_200),
.B(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_198),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_170),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_199),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_178),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_150),
.B1(n_4),
.B2(n_5),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_206),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_150),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_217),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_157),
.Y(n_208)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_166),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_155),
.A2(n_166),
.B1(n_180),
.B2(n_162),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_212),
.A2(n_213),
.B1(n_176),
.B2(n_181),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_214),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_15),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_7),
.C(n_8),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_218),
.A2(n_229),
.B1(n_213),
.B2(n_12),
.Y(n_259)
);

NAND3xp33_ASAP7_75t_L g219 ( 
.A(n_216),
.B(n_165),
.C(n_184),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_201),
.Y(n_257)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_208),
.B(n_163),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_236),
.B(n_196),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_172),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_231),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_156),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_168),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_211),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_182),
.B(n_167),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_239),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_240),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_187),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_246),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_231),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_209),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_212),
.B1(n_202),
.B2(n_193),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_249),
.A2(n_258),
.B1(n_261),
.B2(n_262),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_227),
.B(n_211),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_234),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_264),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_217),
.C(n_190),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_235),
.C(n_238),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_222),
.B(n_236),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_257),
.B(n_230),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_223),
.A2(n_205),
.B1(n_213),
.B2(n_8),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_263),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_213),
.B1(n_9),
.B2(n_8),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_222),
.B(n_10),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_228),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_275),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_232),
.Y(n_272)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_249),
.Y(n_276)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_276),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_233),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_279),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_280),
.B(n_281),
.C(n_263),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_218),
.C(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_237),
.Y(n_282)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_251),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_288),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_255),
.B1(n_245),
.B2(n_258),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_287),
.A2(n_281),
.B1(n_280),
.B2(n_229),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_253),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_179),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_11),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_282),
.A2(n_265),
.B(n_273),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_292),
.B(n_279),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_283),
.C(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_306),
.C(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_299),
.Y(n_311)
);

INVx11_ASAP7_75t_L g300 ( 
.A(n_290),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_301),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_295),
.A2(n_271),
.B1(n_268),
.B2(n_267),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_304),
.B1(n_307),
.B2(n_14),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_303),
.A2(n_12),
.B(n_13),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_297),
.A2(n_271),
.B1(n_267),
.B2(n_250),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_9),
.C(n_11),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_293),
.C(n_287),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g308 ( 
.A(n_283),
.B(n_9),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_308),
.A2(n_291),
.B(n_286),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_315),
.C(n_306),
.Y(n_322)
);

OAI21x1_ASAP7_75t_L g321 ( 
.A1(n_313),
.A2(n_316),
.B(n_308),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_298),
.A2(n_294),
.B(n_288),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_300),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_317),
.B(n_305),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_318),
.B(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_321),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_323),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_304),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_309),
.C(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_319),
.B(n_311),
.Y(n_329)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_329),
.A2(n_321),
.B(n_328),
.Y(n_330)
);

NAND2x1_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_327),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_313),
.B(n_13),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_13),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_14),
.Y(n_334)
);


endmodule