module fake_jpeg_17986_n_81 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_81);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_81;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_0),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_38),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_2),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_39),
.B(n_34),
.Y(n_42)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_30),
.B1(n_32),
.B2(n_29),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_31),
.B1(n_16),
.B2(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_51),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_15),
.B1(n_22),
.B2(n_6),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_57),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_3),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_4),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_41),
.Y(n_60)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_61),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_65),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_7),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_71),
.A2(n_62),
.B(n_56),
.Y(n_72)
);

AO221x1_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B1(n_71),
.B2(n_62),
.C(n_56),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_75),
.A2(n_68),
.B(n_70),
.C(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_68),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_78),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_14),
.C(n_18),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_20),
.Y(n_81)
);


endmodule