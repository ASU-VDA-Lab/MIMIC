module fake_netlist_5_1542_n_1656 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1656);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1656;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_1541;
wire n_172;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVxp67_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_40),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_45),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_58),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_149),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_109),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_50),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_62),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_53),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_18),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_110),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_82),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_4),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_94),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_30),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_86),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_25),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_57),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_78),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_3),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_60),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_26),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_95),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_1),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_41),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_51),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_1),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_104),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_66),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_69),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_87),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_119),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_26),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_142),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_90),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_48),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_15),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_115),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_51),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_120),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_63),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_6),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_39),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_97),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_49),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_10),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_9),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_113),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_108),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_3),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_28),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_132),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_99),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_70),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_89),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_47),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_34),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_13),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_39),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_42),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_68),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_126),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_10),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_48),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_107),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_30),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_52),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_20),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_93),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_32),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_117),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_92),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_14),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_123),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_150),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_103),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_154),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_116),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_130),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_5),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_105),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_54),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_5),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_20),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_138),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_121),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_9),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g269 ( 
.A(n_27),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_65),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_67),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_81),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_46),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_145),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_112),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_31),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_17),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_80),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_18),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_11),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_52),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_12),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_136),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_33),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_56),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_7),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_35),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_71),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_144),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_29),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_37),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_37),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_79),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_44),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_84),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_22),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_74),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_14),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_125),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_306),
.B(n_0),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_191),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_216),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_191),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_6),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_191),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_191),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_160),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_168),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_178),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_180),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_162),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_216),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_175),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_169),
.B(n_7),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_175),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_279),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_167),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_170),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_178),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_183),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_171),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_264),
.Y(n_334)
);

INVxp33_ASAP7_75t_SL g335 ( 
.A(n_157),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_258),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_279),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_169),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_172),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_282),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_172),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_177),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_177),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_186),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_190),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_184),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_190),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_306),
.B(n_8),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_193),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_188),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_264),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_193),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_192),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_231),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_156),
.B(n_11),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_210),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_237),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_231),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_234),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_234),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_239),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_239),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_254),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_194),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_254),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_199),
.Y(n_372)
);

INVxp33_ASAP7_75t_SL g373 ( 
.A(n_159),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_158),
.B(n_12),
.Y(n_374)
);

NOR2xp67_ASAP7_75t_L g375 ( 
.A(n_260),
.B(n_16),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_260),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_166),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_258),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_268),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_246),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_336),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_332),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_318),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_310),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_312),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_312),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_336),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_378),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_327),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_328),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_314),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_315),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_378),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_315),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_316),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_378),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_268),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_323),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_335),
.B(n_229),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_343),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_330),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_320),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_333),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_319),
.B(n_161),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_337),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_R g416 ( 
.A(n_373),
.B(n_173),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_284),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_341),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_340),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_309),
.B(n_200),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_352),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_349),
.B(n_280),
.Y(n_424)
);

AND2x6_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_258),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_351),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_355),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_358),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_361),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_325),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_369),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_374),
.B(n_203),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_362),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_377),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_371),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_354),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_345),
.B(n_218),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_354),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_372),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_345),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_311),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_325),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_416),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_257),
.Y(n_448)
);

BUFx4f_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_406),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_382),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_322),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_380),
.B(n_422),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_403),
.Y(n_454)
);

AND3x2_ASAP7_75t_L g455 ( 
.A(n_408),
.B(n_256),
.C(n_161),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g456 ( 
.A(n_435),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_431),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_414),
.B(n_375),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_422),
.B(n_204),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_414),
.B(n_256),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_403),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_406),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_386),
.Y(n_464)
);

NOR2x1p5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_324),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_414),
.B(n_293),
.Y(n_466)
);

AND2x2_ASAP7_75t_SL g467 ( 
.A(n_433),
.B(n_293),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_409),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_443),
.B(n_426),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_425),
.B(n_258),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_431),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_207),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_158),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_426),
.B(n_347),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_403),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_439),
.A2(n_262),
.B1(n_247),
.B2(n_271),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_375),
.B1(n_313),
.B2(n_324),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_417),
.B(n_258),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_402),
.B(n_163),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_431),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_419),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_425),
.B(n_209),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_419),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_403),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_382),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_339),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_SL g489 ( 
.A(n_402),
.B(n_292),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_420),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_427),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_391),
.B(n_163),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_403),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_405),
.B(n_339),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_431),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_431),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g497 ( 
.A(n_427),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_425),
.Y(n_498)
);

INVx4_ASAP7_75t_L g499 ( 
.A(n_412),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_383),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_425),
.B(n_211),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_421),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_383),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_L g505 ( 
.A(n_425),
.B(n_182),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_385),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_385),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_405),
.B(n_350),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_423),
.B(n_182),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_394),
.B(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_421),
.Y(n_513)
);

AND3x2_ASAP7_75t_L g514 ( 
.A(n_437),
.B(n_348),
.C(n_346),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_384),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_438),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_390),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_387),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

AND2x2_ASAP7_75t_SL g520 ( 
.A(n_438),
.B(n_189),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_440),
.A2(n_313),
.B1(n_290),
.B2(n_295),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_442),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_387),
.Y(n_523)
);

OAI22xp33_ASAP7_75t_L g524 ( 
.A1(n_395),
.A2(n_298),
.B1(n_360),
.B2(n_179),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_407),
.B(n_346),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_388),
.B(n_215),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_390),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_440),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_388),
.B(n_219),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_393),
.B(n_189),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_410),
.B(n_195),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_413),
.B(n_195),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_396),
.B(n_397),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_390),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_396),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g537 ( 
.A(n_398),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_412),
.A2(n_295),
.B1(n_284),
.B2(n_290),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_397),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_399),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_424),
.Y(n_541)
);

BUFx8_ASAP7_75t_SL g542 ( 
.A(n_411),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_415),
.B(n_348),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_418),
.A2(n_360),
.B1(n_251),
.B2(n_248),
.Y(n_544)
);

NAND3xp33_ASAP7_75t_L g545 ( 
.A(n_428),
.B(n_357),
.C(n_187),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_399),
.B(n_220),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_429),
.B(n_197),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_400),
.Y(n_548)
);

BUFx4f_ASAP7_75t_L g549 ( 
.A(n_400),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_444),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_432),
.B(n_197),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_398),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_436),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_441),
.B(n_225),
.Y(n_554)
);

INVx5_ASAP7_75t_L g555 ( 
.A(n_398),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_412),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_412),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_444),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_444),
.B(n_357),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_381),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_444),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_381),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_398),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_401),
.B(n_224),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_430),
.A2(n_213),
.B1(n_212),
.B2(n_217),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_381),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_404),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_401),
.B(n_226),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_404),
.B(n_185),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_404),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_401),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_401),
.B(n_359),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_389),
.B(n_225),
.Y(n_573)
);

BUFx4f_ASAP7_75t_L g574 ( 
.A(n_389),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_389),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_392),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_434),
.A2(n_238),
.B1(n_235),
.B2(n_241),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_392),
.A2(n_249),
.B1(n_250),
.B2(n_253),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_392),
.B(n_227),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_406),
.Y(n_580)
);

INVx1_ASAP7_75t_SL g581 ( 
.A(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_414),
.B(n_227),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_408),
.B(n_196),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_435),
.B(n_379),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_414),
.B(n_236),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_425),
.A2(n_303),
.B1(n_307),
.B2(n_252),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_414),
.B(n_236),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_380),
.B(n_228),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_380),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_380),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_414),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_467),
.B(n_255),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_453),
.B(n_252),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_584),
.B(n_201),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_467),
.A2(n_520),
.B1(n_473),
.B2(n_477),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_543),
.B(n_261),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_L g598 ( 
.A1(n_590),
.A2(n_259),
.B1(n_308),
.B2(n_289),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_456),
.Y(n_599)
);

INVx1_ASAP7_75t_SL g600 ( 
.A(n_581),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_590),
.B(n_202),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_458),
.B(n_259),
.Y(n_602)
);

NAND2xp33_ASAP7_75t_L g603 ( 
.A(n_473),
.B(n_267),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_500),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_458),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_592),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_464),
.B(n_459),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_591),
.B(n_270),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g609 ( 
.A1(n_591),
.A2(n_277),
.B1(n_275),
.B2(n_301),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_500),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_592),
.A2(n_263),
.B1(n_308),
.B2(n_266),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_585),
.B(n_218),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_525),
.B(n_205),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_592),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_520),
.A2(n_303),
.B1(n_307),
.B2(n_266),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_447),
.B(n_474),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_542),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_465),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_448),
.B(n_206),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_452),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_460),
.A2(n_287),
.B1(n_263),
.B2(n_272),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_459),
.B(n_272),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_447),
.B(n_273),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_459),
.B(n_273),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_208),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_473),
.B(n_281),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_473),
.B(n_281),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_503),
.Y(n_628)
);

A2O1A1Ixp33_ASAP7_75t_L g629 ( 
.A1(n_586),
.A2(n_297),
.B(n_289),
.C(n_287),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_489),
.B(n_288),
.C(n_221),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_473),
.B(n_297),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_473),
.B(n_359),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_559),
.B(n_363),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_497),
.B(n_214),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_450),
.B(n_363),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_489),
.B(n_222),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_463),
.Y(n_637)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_545),
.B(n_364),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_586),
.A2(n_291),
.B1(n_223),
.B2(n_230),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_468),
.B(n_364),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_481),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_482),
.B(n_366),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_589),
.B(n_233),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_491),
.Y(n_644)
);

NAND3xp33_ASAP7_75t_L g645 ( 
.A(n_492),
.B(n_294),
.C(n_240),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_484),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_449),
.B(n_242),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_485),
.B(n_366),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_469),
.B(n_243),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_494),
.B(n_244),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_488),
.B(n_265),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_509),
.B(n_367),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_274),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_506),
.Y(n_654)
);

BUFx4_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_586),
.A2(n_300),
.B1(n_276),
.B2(n_278),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_531),
.B(n_304),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_510),
.B(n_491),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_490),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_504),
.B(n_379),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_531),
.B(n_302),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_514),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_511),
.B(n_376),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_516),
.B(n_376),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_533),
.B(n_299),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_449),
.B(n_296),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_528),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_533),
.B(n_305),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_449),
.A2(n_286),
.B1(n_283),
.B2(n_285),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_580),
.B(n_582),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_553),
.B(n_232),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_370),
.C(n_368),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_547),
.B(n_218),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_587),
.A2(n_370),
.B1(n_368),
.B2(n_367),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_537),
.B(n_342),
.Y(n_676)
);

AND2x6_ASAP7_75t_SL g677 ( 
.A(n_519),
.B(n_342),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_532),
.B(n_326),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_518),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_551),
.A2(n_326),
.B1(n_232),
.B2(n_218),
.Y(n_681)
);

OAI22xp5_ASAP7_75t_L g682 ( 
.A1(n_498),
.A2(n_476),
.B1(n_549),
.B2(n_483),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_551),
.B(n_232),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_502),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_554),
.B(n_232),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g686 ( 
.A1(n_479),
.A2(n_17),
.B(n_19),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_513),
.B(n_19),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_540),
.B(n_61),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_548),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_518),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_553),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_523),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_523),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_544),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_451),
.B(n_21),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_499),
.B(n_64),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_498),
.A2(n_72),
.B(n_151),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_567),
.B(n_59),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_567),
.B(n_55),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_522),
.B(n_22),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_478),
.B(n_73),
.Y(n_701)
);

NOR2xp67_ASAP7_75t_L g702 ( 
.A(n_577),
.B(n_77),
.Y(n_702)
);

INVxp67_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_478),
.B(n_152),
.Y(n_704)
);

AOI22xp5_ASAP7_75t_L g705 ( 
.A1(n_479),
.A2(n_147),
.B1(n_146),
.B2(n_133),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_524),
.B(n_23),
.C(n_24),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_519),
.B(n_23),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_499),
.B(n_131),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_510),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_499),
.B(n_122),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_L g711 ( 
.A1(n_549),
.A2(n_118),
.B1(n_111),
.B2(n_106),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_510),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_507),
.B(n_101),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_507),
.B(n_100),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_505),
.A2(n_24),
.B1(n_27),
.B2(n_31),
.Y(n_715)
);

A2O1A1Ixp33_ASAP7_75t_L g716 ( 
.A1(n_461),
.A2(n_32),
.B(n_33),
.C(n_35),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_536),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_507),
.B(n_550),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_515),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_536),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_539),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_526),
.B(n_36),
.Y(n_722)
);

BUFx4_ASAP7_75t_L g723 ( 
.A(n_487),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_461),
.A2(n_98),
.B1(n_96),
.B2(n_91),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_529),
.B(n_36),
.Y(n_725)
);

INVx1_ASAP7_75t_SL g726 ( 
.A(n_487),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_588),
.B(n_88),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_583),
.B(n_38),
.C(n_41),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_539),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_507),
.B(n_50),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_556),
.B(n_38),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_546),
.B(n_42),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_557),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_558),
.B(n_561),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_534),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_560),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_578),
.B(n_43),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_572),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_560),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_583),
.B(n_43),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_508),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_508),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_466),
.B(n_44),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_588),
.B(n_45),
.Y(n_744)
);

AO221x1_ASAP7_75t_L g745 ( 
.A1(n_508),
.A2(n_49),
.B1(n_527),
.B2(n_552),
.C(n_535),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_466),
.B(n_569),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_549),
.B(n_568),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_564),
.B(n_565),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_521),
.B(n_472),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_527),
.B(n_552),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_501),
.A2(n_570),
.B1(n_576),
.B2(n_535),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_576),
.B(n_455),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_538),
.A2(n_563),
.B1(n_527),
.B2(n_535),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_530),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_552),
.B(n_576),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_530),
.A2(n_505),
.B1(n_470),
.B2(n_495),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_445),
.B(n_475),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_571),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_530),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_445),
.B(n_475),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_445),
.B(n_475),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_563),
.A2(n_574),
.B(n_470),
.Y(n_762)
);

INVx3_ASAP7_75t_L g763 ( 
.A(n_614),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_762),
.A2(n_563),
.B(n_574),
.Y(n_764)
);

AOI21x1_ASAP7_75t_L g765 ( 
.A1(n_747),
.A2(n_446),
.B(n_495),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_620),
.B(n_446),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_735),
.B(n_530),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_604),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_614),
.Y(n_769)
);

NOR3xp33_ASAP7_75t_L g770 ( 
.A(n_595),
.B(n_573),
.C(n_457),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_746),
.A2(n_755),
.B(n_607),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_596),
.A2(n_574),
.B(n_457),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_750),
.A2(n_454),
.B(n_493),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_595),
.B(n_530),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_606),
.A2(n_454),
.B(n_493),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_633),
.B(n_530),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_615),
.A2(n_596),
.B1(n_715),
.B2(n_727),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_606),
.A2(n_454),
.B(n_493),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_658),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_757),
.A2(n_496),
.B(n_471),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_615),
.B(n_471),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_610),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_760),
.A2(n_496),
.B(n_480),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_718),
.A2(n_496),
.B(n_480),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_749),
.A2(n_562),
.B(n_573),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_644),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_647),
.A2(n_562),
.B(n_486),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_600),
.B(n_462),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_691),
.Y(n_789)
);

OAI21xp5_ASAP7_75t_L g790 ( 
.A1(n_682),
.A2(n_462),
.B(n_486),
.Y(n_790)
);

O2A1O1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_593),
.A2(n_575),
.B(n_462),
.C(n_486),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_753),
.A2(n_496),
.B(n_517),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_575),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_751),
.A2(n_517),
.B(n_555),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_756),
.A2(n_575),
.B(n_579),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_593),
.A2(n_579),
.B(n_566),
.C(n_555),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_644),
.B(n_566),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_603),
.A2(n_761),
.B(n_734),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_759),
.B(n_579),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_715),
.A2(n_566),
.B1(n_555),
.B2(n_517),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_761),
.A2(n_517),
.B(n_555),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_710),
.A2(n_517),
.B(n_555),
.Y(n_802)
);

NOR2x1_ASAP7_75t_L g803 ( 
.A(n_691),
.B(n_616),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_599),
.B(n_566),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_602),
.A2(n_579),
.B(n_670),
.Y(n_805)
);

AOI22xp5_ASAP7_75t_L g806 ( 
.A1(n_748),
.A2(n_579),
.B1(n_694),
.B2(n_625),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_759),
.A2(n_579),
.B(n_622),
.Y(n_807)
);

NAND2x1p5_ASAP7_75t_L g808 ( 
.A(n_754),
.B(n_658),
.Y(n_808)
);

NAND2x1_ASAP7_75t_L g809 ( 
.A(n_736),
.B(n_739),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_628),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_686),
.A2(n_744),
.B(n_740),
.C(n_703),
.Y(n_811)
);

AOI21x1_ASAP7_75t_L g812 ( 
.A1(n_647),
.A2(n_666),
.B(n_632),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_759),
.A2(n_624),
.B(n_708),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_740),
.A2(n_744),
.B(n_737),
.C(n_716),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_613),
.B(n_738),
.Y(n_815)
);

BUFx2_ASAP7_75t_L g816 ( 
.A(n_680),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_709),
.B(n_712),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_727),
.A2(n_683),
.B1(n_674),
.B2(n_594),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_687),
.Y(n_819)
);

INVx1_ASAP7_75t_SL g820 ( 
.A(n_652),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_626),
.A2(n_631),
.B(n_627),
.Y(n_821)
);

AOI21x1_ASAP7_75t_L g822 ( 
.A1(n_666),
.A2(n_699),
.B(n_698),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_672),
.B(n_625),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_743),
.A2(n_697),
.B(n_701),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_696),
.A2(n_708),
.B(n_676),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_696),
.A2(n_704),
.B(n_742),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_741),
.A2(n_714),
.B(n_713),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_733),
.A2(n_690),
.B(n_654),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_654),
.A2(n_690),
.B(n_671),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_619),
.B(n_674),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_671),
.A2(n_720),
.B(n_693),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_637),
.B(n_641),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_619),
.B(n_623),
.Y(n_833)
);

O2A1O1Ixp33_ASAP7_75t_L g834 ( 
.A1(n_621),
.A2(n_598),
.B(n_725),
.C(n_732),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_677),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_646),
.B(n_659),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_683),
.A2(n_653),
.B1(n_722),
.B2(n_725),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_667),
.B(n_689),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_722),
.A2(n_732),
.B(n_629),
.C(n_731),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_679),
.A2(n_693),
.B(n_717),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_612),
.B(n_649),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_679),
.A2(n_717),
.B(n_720),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_605),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_643),
.A2(n_748),
.B(n_653),
.C(n_636),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_649),
.B(n_601),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_688),
.A2(n_758),
.B(n_692),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_726),
.B(n_601),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_721),
.A2(n_729),
.B(n_608),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_739),
.A2(n_754),
.B(n_597),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_700),
.B(n_651),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_707),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_730),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_752),
.A2(n_702),
.B1(n_630),
.B2(n_618),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_678),
.Y(n_854)
);

NAND3xp33_ASAP7_75t_L g855 ( 
.A(n_645),
.B(n_639),
.C(n_656),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_634),
.A2(n_642),
.B(n_663),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_635),
.A2(n_660),
.B(n_664),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_662),
.Y(n_858)
);

AO21x1_ASAP7_75t_L g859 ( 
.A1(n_711),
.A2(n_728),
.B(n_668),
.Y(n_859)
);

AOI21x1_ASAP7_75t_L g860 ( 
.A1(n_640),
.A2(n_648),
.B(n_638),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_745),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_673),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_695),
.Y(n_863)
);

INVxp67_ASAP7_75t_L g864 ( 
.A(n_719),
.Y(n_864)
);

INVxp67_ASAP7_75t_L g865 ( 
.A(n_650),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_681),
.A2(n_611),
.B1(n_705),
.B2(n_724),
.Y(n_866)
);

O2A1O1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_657),
.A2(n_661),
.B(n_665),
.C(n_685),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_752),
.A2(n_675),
.B(n_609),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_669),
.B(n_617),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_723),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_706),
.A2(n_449),
.B(n_762),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_655),
.B(n_456),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_599),
.Y(n_873)
);

INVx4_ASAP7_75t_L g874 ( 
.A(n_614),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_684),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_644),
.Y(n_877)
);

AO32x1_ASAP7_75t_L g878 ( 
.A1(n_621),
.A2(n_711),
.A3(n_682),
.B1(n_721),
.B2(n_692),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_595),
.A2(n_683),
.B(n_674),
.C(n_653),
.Y(n_879)
);

AND2x2_ASAP7_75t_SL g880 ( 
.A(n_615),
.B(n_451),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_644),
.B(n_658),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_735),
.B(n_453),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_613),
.A2(n_584),
.B(n_625),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_735),
.B(n_453),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_735),
.B(n_453),
.Y(n_887)
);

AOI21xp33_ASAP7_75t_L g888 ( 
.A1(n_595),
.A2(n_467),
.B(n_596),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_889)
);

INVx4_ASAP7_75t_L g890 ( 
.A(n_614),
.Y(n_890)
);

O2A1O1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_593),
.A2(n_686),
.B(n_744),
.C(n_740),
.Y(n_891)
);

BUFx6f_ASAP7_75t_L g892 ( 
.A(n_644),
.Y(n_892)
);

NAND2x1_ASAP7_75t_L g893 ( 
.A(n_606),
.B(n_592),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_735),
.B(n_453),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_604),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_615),
.A2(n_596),
.B1(n_715),
.B2(n_477),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_735),
.B(n_453),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_644),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_604),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_SL g902 ( 
.A1(n_701),
.A2(n_704),
.B(n_697),
.C(n_696),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_735),
.B(n_453),
.Y(n_903)
);

CKINVDCx10_ASAP7_75t_R g904 ( 
.A(n_655),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_595),
.A2(n_607),
.B1(n_748),
.B2(n_596),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_615),
.A2(n_596),
.B1(n_715),
.B2(n_477),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_620),
.B(n_585),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_735),
.B(n_453),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_735),
.B(n_453),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_607),
.B(n_456),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_644),
.B(n_658),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_644),
.B(n_658),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_735),
.B(n_453),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_604),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_607),
.B(n_456),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_595),
.B(n_456),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_735),
.B(n_453),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_620),
.B(n_585),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_919)
);

BUFx2_ASAP7_75t_L g920 ( 
.A(n_599),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_595),
.A2(n_607),
.B1(n_748),
.B2(n_596),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_595),
.B(n_456),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_600),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_615),
.A2(n_596),
.B1(n_715),
.B2(n_477),
.Y(n_924)
);

NAND2xp33_ASAP7_75t_L g925 ( 
.A(n_596),
.B(n_615),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_607),
.B(n_456),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_735),
.B(n_453),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_930)
);

BUFx2_ASAP7_75t_L g931 ( 
.A(n_599),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_684),
.Y(n_932)
);

A2O1A1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_595),
.A2(n_683),
.B(n_674),
.C(n_653),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_735),
.B(n_453),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_735),
.B(n_453),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_762),
.A2(n_449),
.B(n_747),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_595),
.A2(n_607),
.B1(n_748),
.B2(n_596),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_595),
.B(n_456),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_599),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_596),
.A2(n_749),
.B(n_467),
.Y(n_941)
);

OAI21xp5_ASAP7_75t_L g942 ( 
.A1(n_596),
.A2(n_749),
.B(n_467),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_735),
.B(n_453),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_786),
.Y(n_944)
);

INVxp67_ASAP7_75t_L g945 ( 
.A(n_873),
.Y(n_945)
);

NOR2x1_ASAP7_75t_SL g946 ( 
.A(n_777),
.B(n_897),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_875),
.A2(n_884),
.B(n_882),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_889),
.A2(n_899),
.B(n_895),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_780),
.A2(n_783),
.B(n_765),
.Y(n_950)
);

AO21x1_ASAP7_75t_L g951 ( 
.A1(n_837),
.A2(n_818),
.B(n_777),
.Y(n_951)
);

OR2x6_ASAP7_75t_L g952 ( 
.A(n_870),
.B(n_932),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_825),
.A2(n_771),
.B(n_919),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_883),
.B(n_886),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_879),
.A2(n_933),
.B(n_885),
.C(n_833),
.Y(n_955)
);

O2A1O1Ixp5_ASAP7_75t_L g956 ( 
.A1(n_837),
.A2(n_830),
.B(n_845),
.C(n_818),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_773),
.A2(n_842),
.B(n_827),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_887),
.B(n_894),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_768),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_926),
.A2(n_930),
.B(n_928),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_842),
.A2(n_784),
.B(n_935),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_923),
.Y(n_962)
);

AOI21x1_ASAP7_75t_L g963 ( 
.A1(n_937),
.A2(n_798),
.B(n_812),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_881),
.B(n_911),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_941),
.A2(n_942),
.B(n_888),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_829),
.A2(n_840),
.B(n_831),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_898),
.B(n_903),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_888),
.A2(n_906),
.B(n_897),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_782),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_941),
.A2(n_942),
.B(n_921),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_916),
.B(n_922),
.Y(n_971)
);

BUFx4f_ASAP7_75t_SL g972 ( 
.A(n_923),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_939),
.B(n_907),
.Y(n_973)
);

OAI21x1_ASAP7_75t_SL g974 ( 
.A1(n_859),
.A2(n_906),
.B(n_924),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_908),
.B(n_909),
.Y(n_975)
);

OAI21x1_ASAP7_75t_L g976 ( 
.A1(n_795),
.A2(n_826),
.B(n_792),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_813),
.A2(n_902),
.B(n_774),
.Y(n_977)
);

NOR2x1_ASAP7_75t_SL g978 ( 
.A(n_924),
.B(n_800),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_821),
.A2(n_824),
.B(n_776),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_820),
.Y(n_980)
);

AO31x2_ASAP7_75t_L g981 ( 
.A1(n_866),
.A2(n_871),
.A3(n_861),
.B(n_805),
.Y(n_981)
);

AO31x2_ASAP7_75t_L g982 ( 
.A1(n_866),
.A2(n_793),
.A3(n_800),
.B(n_846),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_905),
.A2(n_938),
.B(n_891),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_795),
.A2(n_790),
.B(n_828),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_918),
.B(n_820),
.Y(n_985)
);

NAND2x1p5_ASAP7_75t_L g986 ( 
.A(n_789),
.B(n_893),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_821),
.A2(n_824),
.B(n_772),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_913),
.A2(n_936),
.B1(n_917),
.B2(n_934),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_790),
.A2(n_778),
.B(n_775),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_929),
.B(n_943),
.Y(n_990)
);

OR2x6_ASAP7_75t_L g991 ( 
.A(n_870),
.B(n_920),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_841),
.A2(n_925),
.B1(n_823),
.B2(n_806),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_815),
.B(n_854),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_870),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_772),
.A2(n_799),
.B(n_857),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_931),
.B(n_940),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_847),
.B(n_819),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_880),
.A2(n_850),
.B1(n_915),
.B2(n_910),
.Y(n_998)
);

OAI21xp5_ASAP7_75t_L g999 ( 
.A1(n_814),
.A2(n_811),
.B(n_781),
.Y(n_999)
);

AOI221x1_ASAP7_75t_L g1000 ( 
.A1(n_770),
.A2(n_868),
.B1(n_852),
.B2(n_856),
.C(n_855),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_767),
.A2(n_807),
.B(n_849),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_834),
.A2(n_844),
.B(n_839),
.C(n_867),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_781),
.A2(n_796),
.B(n_797),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_797),
.A2(n_791),
.B(n_848),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_L g1005 ( 
.A1(n_802),
.A2(n_822),
.B(n_794),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_816),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_852),
.B(n_862),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_851),
.B(n_927),
.Y(n_1008)
);

OAI22x1_ASAP7_75t_L g1009 ( 
.A1(n_853),
.A2(n_869),
.B1(n_865),
.B2(n_863),
.Y(n_1009)
);

INVx11_ASAP7_75t_L g1010 ( 
.A(n_904),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_SL g1011 ( 
.A1(n_860),
.A2(n_838),
.B(n_836),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_786),
.Y(n_1012)
);

INVx6_ASAP7_75t_L g1013 ( 
.A(n_858),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_858),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_864),
.B(n_789),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_809),
.A2(n_801),
.B(n_914),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_788),
.B(n_863),
.Y(n_1017)
);

AO31x2_ASAP7_75t_L g1018 ( 
.A1(n_878),
.A2(n_810),
.A3(n_901),
.B(n_896),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_786),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_763),
.A2(n_769),
.B(n_804),
.Y(n_1020)
);

OAI21x1_ASAP7_75t_L g1021 ( 
.A1(n_843),
.A2(n_808),
.B(n_769),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_808),
.A2(n_763),
.B(n_779),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_858),
.B(n_877),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_881),
.A2(n_912),
.B(n_911),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_912),
.A2(n_779),
.B(n_878),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_832),
.B(n_766),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_803),
.B(n_832),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_835),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_878),
.A2(n_874),
.B(n_890),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_817),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_817),
.A2(n_874),
.B(n_890),
.Y(n_1031)
);

NAND2xp33_ASAP7_75t_L g1032 ( 
.A(n_877),
.B(n_892),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_877),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_892),
.B(n_900),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_892),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_900),
.A2(n_785),
.B(n_764),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_900),
.A2(n_785),
.B(n_764),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_872),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_837),
.A2(n_879),
.A3(n_933),
.B(n_818),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_L g1040 ( 
.A(n_885),
.B(n_933),
.C(n_879),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_SL g1041 ( 
.A(n_777),
.B(n_897),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_825),
.A2(n_771),
.B(n_875),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_825),
.A2(n_771),
.B(n_875),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_879),
.A2(n_933),
.B(n_941),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_876),
.Y(n_1046)
);

INVx1_ASAP7_75t_SL g1047 ( 
.A(n_923),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_875),
.A2(n_449),
.B(n_762),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_881),
.B(n_911),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_786),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_SL g1053 ( 
.A1(n_777),
.A2(n_906),
.B(n_897),
.Y(n_1053)
);

OAI21x1_ASAP7_75t_L g1054 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_916),
.B(n_922),
.Y(n_1055)
);

BUFx5_ASAP7_75t_L g1056 ( 
.A(n_768),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1057)
);

AOI21x1_ASAP7_75t_SL g1058 ( 
.A1(n_774),
.A2(n_845),
.B(n_767),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_881),
.B(n_911),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_916),
.B(n_456),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_879),
.A2(n_933),
.B(n_941),
.Y(n_1061)
);

OAI21x1_ASAP7_75t_L g1062 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_L g1063 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_768),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_883),
.B(n_886),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_825),
.A2(n_771),
.B(n_875),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_787),
.A2(n_765),
.B(n_875),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_879),
.A2(n_933),
.B(n_885),
.C(n_833),
.Y(n_1069)
);

OR2x2_ASAP7_75t_L g1070 ( 
.A(n_820),
.B(n_456),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_875),
.A2(n_449),
.B(n_762),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_916),
.B(n_922),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_879),
.A2(n_933),
.B(n_885),
.C(n_833),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_825),
.A2(n_771),
.B(n_875),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_916),
.B(n_456),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_883),
.B(n_886),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_785),
.A2(n_764),
.B(n_787),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_883),
.B(n_886),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_SL g1080 ( 
.A1(n_777),
.A2(n_906),
.B(n_897),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_883),
.B(n_886),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_879),
.A2(n_933),
.B(n_885),
.C(n_833),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_944),
.Y(n_1083)
);

AOI21xp33_ASAP7_75t_SL g1084 ( 
.A1(n_1055),
.A2(n_1072),
.B(n_1009),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_954),
.B(n_958),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1070),
.B(n_996),
.Y(n_1086)
);

NAND2xp33_ASAP7_75t_L g1087 ( 
.A(n_1040),
.B(n_955),
.Y(n_1087)
);

AOI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_971),
.A2(n_1060),
.B1(n_1076),
.B2(n_973),
.Y(n_1088)
);

OR2x2_ASAP7_75t_L g1089 ( 
.A(n_954),
.B(n_958),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_972),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1013),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_967),
.B(n_975),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_959),
.Y(n_1093)
);

HB1xp67_ASAP7_75t_L g1094 ( 
.A(n_1047),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_962),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_967),
.B(n_975),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_998),
.A2(n_988),
.B1(n_1017),
.B2(n_997),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1010),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_985),
.B(n_1008),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_969),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1047),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_L g1102 ( 
.A(n_1069),
.B(n_1074),
.C(n_1082),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_990),
.A2(n_1077),
.B1(n_1065),
.B2(n_1081),
.Y(n_1103)
);

INVx5_ASAP7_75t_L g1104 ( 
.A(n_944),
.Y(n_1104)
);

AOI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_951),
.A2(n_968),
.B1(n_983),
.B2(n_974),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1064),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_964),
.B(n_1050),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_990),
.A2(n_1081),
.B1(n_1065),
.B2(n_1079),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_980),
.Y(n_1109)
);

INVx3_ASAP7_75t_SL g1110 ( 
.A(n_994),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1042),
.A2(n_1067),
.B(n_1075),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1077),
.B(n_1079),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_964),
.B(n_1050),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_980),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1075),
.A2(n_995),
.B(n_977),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_946),
.A2(n_1041),
.B1(n_978),
.B2(n_983),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_988),
.B(n_993),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_993),
.B(n_1006),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_L g1119 ( 
.A1(n_1044),
.A2(n_1061),
.B(n_956),
.C(n_949),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_948),
.A2(n_960),
.B(n_1048),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1026),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_991),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1026),
.B(n_945),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1059),
.B(n_1038),
.Y(n_1124)
);

OR2x6_ASAP7_75t_L g1125 ( 
.A(n_991),
.B(n_952),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_1059),
.B(n_1030),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_992),
.A2(n_1044),
.B1(n_1061),
.B2(n_1080),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_1013),
.Y(n_1128)
);

NAND2x1p5_ASAP7_75t_L g1129 ( 
.A(n_944),
.B(n_1012),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1033),
.B(n_1046),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1007),
.B(n_999),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1007),
.B(n_999),
.Y(n_1132)
);

OR2x2_ASAP7_75t_SL g1133 ( 
.A(n_1034),
.B(n_1035),
.Y(n_1133)
);

NOR2xp67_ASAP7_75t_SL g1134 ( 
.A(n_1053),
.B(n_1028),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_1071),
.A2(n_987),
.B(n_979),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1012),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1023),
.B(n_1015),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1024),
.B(n_970),
.Y(n_1138)
);

INVx3_ASAP7_75t_SL g1139 ( 
.A(n_952),
.Y(n_1139)
);

NOR2xp67_ASAP7_75t_L g1140 ( 
.A(n_1014),
.B(n_1031),
.Y(n_1140)
);

AOI222xp33_ASAP7_75t_L g1141 ( 
.A1(n_970),
.A2(n_965),
.B1(n_1002),
.B2(n_1027),
.C1(n_1032),
.C2(n_1011),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1039),
.B(n_965),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1039),
.B(n_979),
.Y(n_1143)
);

INVx1_ASAP7_75t_SL g1144 ( 
.A(n_952),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1012),
.B(n_1019),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1001),
.A2(n_1000),
.B(n_1004),
.Y(n_1146)
);

NOR2x1_ASAP7_75t_L g1147 ( 
.A(n_1019),
.B(n_1052),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_1019),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_1052),
.B(n_1022),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_1052),
.Y(n_1150)
);

CKINVDCx6p67_ASAP7_75t_R g1151 ( 
.A(n_1056),
.Y(n_1151)
);

INVx3_ASAP7_75t_L g1152 ( 
.A(n_986),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1039),
.B(n_981),
.Y(n_1153)
);

NAND2xp33_ASAP7_75t_L g1154 ( 
.A(n_986),
.B(n_1020),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1021),
.B(n_981),
.Y(n_1155)
);

CKINVDCx8_ASAP7_75t_R g1156 ( 
.A(n_1058),
.Y(n_1156)
);

HB1xp67_ASAP7_75t_L g1157 ( 
.A(n_981),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1025),
.B(n_982),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1003),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1018),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_982),
.B(n_984),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1018),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1036),
.B(n_1037),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_982),
.B(n_1029),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_976),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_1016),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_961),
.B(n_1005),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_963),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1068),
.B(n_957),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_950),
.Y(n_1170)
);

AOI21x1_ASAP7_75t_L g1171 ( 
.A1(n_947),
.A2(n_1057),
.B(n_1073),
.Y(n_1171)
);

INVx4_ASAP7_75t_L g1172 ( 
.A(n_1045),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1049),
.B(n_1062),
.Y(n_1173)
);

NOR2xp33_ASAP7_75t_L g1174 ( 
.A(n_989),
.B(n_966),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1051),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1054),
.A2(n_1063),
.B(n_1066),
.C(n_1078),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_964),
.B(n_1050),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1010),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_953),
.A2(n_1043),
.B(n_1042),
.Y(n_1179)
);

OR2x2_ASAP7_75t_L g1180 ( 
.A(n_1070),
.B(n_456),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1055),
.A2(n_879),
.B1(n_933),
.B2(n_1072),
.Y(n_1181)
);

AO22x1_ASAP7_75t_L g1182 ( 
.A1(n_1055),
.A2(n_1072),
.B1(n_916),
.B2(n_939),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_972),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_944),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1055),
.B(n_1072),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_955),
.A2(n_777),
.B(n_906),
.C(n_897),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_964),
.B(n_1050),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_944),
.Y(n_1188)
);

INVx2_ASAP7_75t_SL g1189 ( 
.A(n_972),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_959),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_954),
.Y(n_1191)
);

NAND2x1p5_ASAP7_75t_L g1192 ( 
.A(n_944),
.B(n_789),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_972),
.Y(n_1193)
);

CKINVDCx11_ASAP7_75t_R g1194 ( 
.A(n_994),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1055),
.B(n_1072),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1060),
.B(n_1076),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_953),
.A2(n_1043),
.B(n_1042),
.Y(n_1197)
);

INVx5_ASAP7_75t_L g1198 ( 
.A(n_944),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1010),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_951),
.A2(n_777),
.B1(n_837),
.B2(n_1040),
.Y(n_1200)
);

A2O1A1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1040),
.A2(n_595),
.B(n_837),
.C(n_1044),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1055),
.A2(n_879),
.B1(n_933),
.B2(n_1072),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1055),
.B(n_1072),
.Y(n_1203)
);

AND2x4_ASAP7_75t_SL g1204 ( 
.A(n_991),
.B(n_952),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1055),
.B(n_1072),
.Y(n_1205)
);

BUFx6f_ASAP7_75t_L g1206 ( 
.A(n_944),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_1055),
.B(n_1072),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1207),
.A2(n_1202),
.B1(n_1181),
.B2(n_1087),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1104),
.Y(n_1209)
);

NAND3xp33_ASAP7_75t_SL g1210 ( 
.A(n_1207),
.B(n_1084),
.C(n_1185),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1087),
.A2(n_1102),
.B1(n_1127),
.B2(n_1200),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1093),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1102),
.A2(n_1200),
.B1(n_1203),
.B2(n_1195),
.Y(n_1213)
);

AOI21xp33_ASAP7_75t_L g1214 ( 
.A1(n_1201),
.A2(n_1159),
.B(n_1205),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1085),
.A2(n_1096),
.B1(n_1092),
.B2(n_1089),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1182),
.A2(n_1191),
.B1(n_1112),
.B2(n_1108),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1100),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1094),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1107),
.B(n_1113),
.Y(n_1219)
);

BUFx6f_ASAP7_75t_SL g1220 ( 
.A(n_1095),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1106),
.Y(n_1221)
);

NAND2x1p5_ASAP7_75t_L g1222 ( 
.A(n_1104),
.B(n_1198),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1120),
.Y(n_1223)
);

OAI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1191),
.A2(n_1117),
.B1(n_1103),
.B2(n_1097),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1137),
.A2(n_1196),
.B1(n_1099),
.B2(n_1204),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1121),
.B(n_1105),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1190),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1176),
.A2(n_1120),
.B(n_1115),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1198),
.B(n_1152),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1134),
.A2(n_1116),
.B1(n_1105),
.B2(n_1088),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1142),
.B(n_1143),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1198),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1146),
.A2(n_1115),
.B(n_1179),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1151),
.Y(n_1234)
);

OAI21xp33_ASAP7_75t_L g1235 ( 
.A1(n_1186),
.A2(n_1180),
.B(n_1116),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1138),
.A2(n_1124),
.B1(n_1141),
.B2(n_1095),
.Y(n_1236)
);

OAI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1110),
.A2(n_1086),
.B1(n_1118),
.B2(n_1121),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1123),
.B(n_1131),
.Y(n_1238)
);

BUFx3_ASAP7_75t_L g1239 ( 
.A(n_1090),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1107),
.A2(n_1177),
.B1(n_1113),
.B2(n_1187),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1132),
.B(n_1094),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1122),
.A2(n_1101),
.B1(n_1125),
.B2(n_1109),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1126),
.A2(n_1177),
.B1(n_1187),
.B2(n_1101),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1170),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_SL g1246 ( 
.A1(n_1125),
.A2(n_1144),
.B1(n_1201),
.B2(n_1114),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1110),
.A2(n_1125),
.B1(n_1139),
.B2(n_1193),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1186),
.B(n_1158),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1133),
.A2(n_1156),
.B1(n_1139),
.B2(n_1168),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1155),
.A2(n_1194),
.B1(n_1153),
.B2(n_1165),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1155),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1194),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1111),
.A2(n_1197),
.B(n_1135),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1140),
.A2(n_1130),
.B1(n_1164),
.B2(n_1157),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1136),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_R g1256 ( 
.A(n_1098),
.B(n_1199),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1157),
.B(n_1149),
.Y(n_1257)
);

OAI21xp5_ASAP7_75t_SL g1258 ( 
.A1(n_1183),
.A2(n_1189),
.B(n_1192),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1091),
.B(n_1128),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1119),
.B(n_1162),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1178),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1154),
.A2(n_1145),
.B1(n_1192),
.B2(n_1150),
.Y(n_1262)
);

OAI21xp5_ASAP7_75t_L g1263 ( 
.A1(n_1119),
.A2(n_1169),
.B(n_1174),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1161),
.A2(n_1169),
.B1(n_1174),
.B2(n_1167),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1129),
.Y(n_1265)
);

BUFx10_ASAP7_75t_L g1266 ( 
.A(n_1145),
.Y(n_1266)
);

AO21x2_ASAP7_75t_L g1267 ( 
.A1(n_1175),
.A2(n_1173),
.B(n_1163),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1160),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1083),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1163),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1147),
.B(n_1083),
.Y(n_1271)
);

OR2x2_ASAP7_75t_L g1272 ( 
.A(n_1172),
.B(n_1166),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1148),
.B(n_1083),
.Y(n_1273)
);

OAI22xp5_ASAP7_75t_L g1274 ( 
.A1(n_1184),
.A2(n_1206),
.B1(n_1188),
.B2(n_1166),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1188),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_1206),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1207),
.B(n_1055),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1151),
.Y(n_1278)
);

AO21x1_ASAP7_75t_SL g1279 ( 
.A1(n_1200),
.A2(n_1061),
.B(n_1044),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_1194),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1207),
.A2(n_1055),
.B1(n_1072),
.B2(n_885),
.Y(n_1281)
);

HB1xp67_ASAP7_75t_L g1282 ( 
.A(n_1094),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1207),
.A2(n_1055),
.B1(n_1072),
.B2(n_777),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1207),
.A2(n_1055),
.B1(n_1072),
.B2(n_885),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1181),
.A2(n_837),
.B(n_1202),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_SL g1286 ( 
.A1(n_1207),
.A2(n_1055),
.B1(n_1072),
.B2(n_777),
.Y(n_1286)
);

BUFx2_ASAP7_75t_L g1287 ( 
.A(n_1094),
.Y(n_1287)
);

BUFx2_ASAP7_75t_R g1288 ( 
.A(n_1110),
.Y(n_1288)
);

INVx1_ASAP7_75t_SL g1289 ( 
.A(n_1086),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1093),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1086),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1151),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_1094),
.Y(n_1293)
);

INVx6_ASAP7_75t_L g1294 ( 
.A(n_1104),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1094),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1207),
.A2(n_1055),
.B1(n_1072),
.B2(n_777),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_SL g1297 ( 
.A1(n_1117),
.A2(n_951),
.B(n_978),
.Y(n_1297)
);

INVx3_ASAP7_75t_L g1298 ( 
.A(n_1151),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1171),
.A2(n_1176),
.B(n_1005),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1151),
.Y(n_1300)
);

BUFx2_ASAP7_75t_R g1301 ( 
.A(n_1110),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1268),
.Y(n_1302)
);

OAI21xp33_ASAP7_75t_L g1303 ( 
.A1(n_1283),
.A2(n_1296),
.B(n_1286),
.Y(n_1303)
);

HB1xp67_ASAP7_75t_L g1304 ( 
.A(n_1267),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1260),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1267),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1231),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1231),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_1267),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1270),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1257),
.Y(n_1311)
);

NOR2xp33_ASAP7_75t_L g1312 ( 
.A(n_1210),
.B(n_1277),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1248),
.B(n_1279),
.Y(n_1313)
);

OAI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1208),
.A2(n_1284),
.B(n_1281),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1279),
.B(n_1263),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1251),
.B(n_1264),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1251),
.B(n_1226),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1218),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1253),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1218),
.Y(n_1320)
);

HB1xp67_ASAP7_75t_L g1321 ( 
.A(n_1287),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1223),
.A2(n_1299),
.B(n_1228),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1226),
.B(n_1285),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1287),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1285),
.B(n_1233),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1272),
.Y(n_1326)
);

OAI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1214),
.A2(n_1211),
.B(n_1224),
.Y(n_1327)
);

INVxp67_ASAP7_75t_SL g1328 ( 
.A(n_1282),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1223),
.Y(n_1329)
);

OR2x2_ASAP7_75t_L g1330 ( 
.A(n_1241),
.B(n_1293),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1295),
.Y(n_1331)
);

AOI222xp33_ASAP7_75t_L g1332 ( 
.A1(n_1213),
.A2(n_1235),
.B1(n_1215),
.B2(n_1230),
.C1(n_1291),
.C2(n_1289),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1297),
.A2(n_1274),
.B(n_1237),
.Y(n_1333)
);

NAND2xp33_ASAP7_75t_R g1334 ( 
.A(n_1244),
.B(n_1234),
.Y(n_1334)
);

AO21x2_ASAP7_75t_L g1335 ( 
.A1(n_1297),
.A2(n_1217),
.B(n_1227),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1238),
.B(n_1216),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1254),
.A2(n_1250),
.B(n_1236),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1249),
.B(n_1225),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1247),
.A2(n_1246),
.B1(n_1243),
.B2(n_1212),
.Y(n_1339)
);

NOR2xp33_ASAP7_75t_L g1340 ( 
.A(n_1258),
.B(n_1245),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1255),
.B(n_1239),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1266),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1221),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1290),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1262),
.B(n_1242),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1266),
.Y(n_1346)
);

INVx1_ASAP7_75t_SL g1347 ( 
.A(n_1266),
.Y(n_1347)
);

INVx11_ASAP7_75t_L g1348 ( 
.A(n_1269),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1294),
.Y(n_1349)
);

INVxp67_ASAP7_75t_L g1350 ( 
.A(n_1220),
.Y(n_1350)
);

AO21x2_ASAP7_75t_L g1351 ( 
.A1(n_1271),
.A2(n_1240),
.B(n_1273),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1352)
);

INVxp67_ASAP7_75t_SL g1353 ( 
.A(n_1318),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1315),
.B(n_1265),
.Y(n_1354)
);

INVx3_ASAP7_75t_L g1355 ( 
.A(n_1306),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1319),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1304),
.Y(n_1357)
);

INVx5_ASAP7_75t_SL g1358 ( 
.A(n_1333),
.Y(n_1358)
);

OR2x2_ASAP7_75t_L g1359 ( 
.A(n_1325),
.B(n_1278),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1315),
.B(n_1265),
.Y(n_1360)
);

HB1xp67_ASAP7_75t_L g1361 ( 
.A(n_1335),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1310),
.B(n_1292),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1315),
.B(n_1219),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1318),
.Y(n_1364)
);

OAI31xp33_ASAP7_75t_L g1365 ( 
.A1(n_1303),
.A2(n_1252),
.A3(n_1219),
.B(n_1229),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1325),
.B(n_1219),
.Y(n_1366)
);

INVxp67_ASAP7_75t_L g1367 ( 
.A(n_1320),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1302),
.Y(n_1368)
);

OR2x2_ASAP7_75t_L g1369 ( 
.A(n_1325),
.B(n_1300),
.Y(n_1369)
);

AOI222xp33_ASAP7_75t_L g1370 ( 
.A1(n_1314),
.A2(n_1280),
.B1(n_1220),
.B2(n_1256),
.C1(n_1259),
.C2(n_1301),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1308),
.B(n_1298),
.Y(n_1371)
);

NAND2x1_ASAP7_75t_L g1372 ( 
.A(n_1306),
.B(n_1298),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_1306),
.B(n_1305),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1313),
.B(n_1292),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1308),
.B(n_1278),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1320),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1314),
.A2(n_1220),
.B1(n_1280),
.B2(n_1275),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1312),
.B(n_1288),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1323),
.B(n_1276),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1323),
.B(n_1229),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1343),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1335),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1303),
.A2(n_1269),
.B1(n_1275),
.B2(n_1294),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_SL g1384 ( 
.A(n_1334),
.B(n_1261),
.C(n_1222),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1330),
.B(n_1209),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1330),
.B(n_1232),
.Y(n_1386)
);

OAI221xp5_ASAP7_75t_L g1387 ( 
.A1(n_1377),
.A2(n_1312),
.B1(n_1370),
.B2(n_1365),
.C(n_1338),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1378),
.B(n_1350),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1353),
.B(n_1330),
.Y(n_1389)
);

OR2x2_ASAP7_75t_SL g1390 ( 
.A(n_1359),
.B(n_1337),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1366),
.B(n_1311),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1385),
.B(n_1328),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1373),
.B(n_1311),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1366),
.B(n_1317),
.Y(n_1394)
);

NAND3xp33_ASAP7_75t_L g1395 ( 
.A(n_1370),
.B(n_1332),
.C(n_1327),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1353),
.B(n_1321),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1377),
.B(n_1332),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1366),
.B(n_1317),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1364),
.B(n_1321),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1354),
.B(n_1317),
.Y(n_1400)
);

NAND3xp33_ASAP7_75t_L g1401 ( 
.A(n_1365),
.B(n_1327),
.C(n_1336),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1354),
.B(n_1360),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1385),
.B(n_1386),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1361),
.A2(n_1322),
.B(n_1329),
.Y(n_1404)
);

AOI221xp5_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1336),
.B1(n_1340),
.B2(n_1338),
.C(n_1341),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1383),
.B(n_1339),
.C(n_1345),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1386),
.B(n_1352),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1374),
.A2(n_1337),
.B1(n_1345),
.B2(n_1351),
.Y(n_1408)
);

NAND2xp33_ASAP7_75t_SL g1409 ( 
.A(n_1384),
.B(n_1334),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1364),
.B(n_1324),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_1324),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1367),
.B(n_1328),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1363),
.B(n_1350),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1374),
.A2(n_1337),
.B1(n_1351),
.B2(n_1339),
.Y(n_1414)
);

NAND2xp33_ASAP7_75t_SL g1415 ( 
.A(n_1384),
.B(n_1349),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_SL g1416 ( 
.A(n_1379),
.B(n_1349),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1381),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1359),
.B(n_1326),
.Y(n_1418)
);

AOI211xp5_ASAP7_75t_L g1419 ( 
.A1(n_1379),
.A2(n_1340),
.B(n_1341),
.C(n_1342),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1371),
.B(n_1331),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1376),
.B(n_1368),
.Y(n_1421)
);

OA21x2_ASAP7_75t_L g1422 ( 
.A1(n_1361),
.A2(n_1322),
.B(n_1329),
.Y(n_1422)
);

AOI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1375),
.A2(n_1347),
.B1(n_1346),
.B2(n_1342),
.C(n_1344),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1381),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1369),
.B(n_1309),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1379),
.A2(n_1316),
.B(n_1347),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1369),
.B(n_1309),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1419),
.B(n_1362),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1425),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_SL g1430 ( 
.A(n_1419),
.B(n_1362),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1402),
.B(n_1358),
.Y(n_1431)
);

AND2x4_ASAP7_75t_L g1432 ( 
.A(n_1427),
.B(n_1355),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1417),
.Y(n_1433)
);

OR2x2_ASAP7_75t_L g1434 ( 
.A(n_1390),
.B(n_1373),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1407),
.B(n_1403),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1417),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1389),
.B(n_1357),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1424),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1402),
.B(n_1358),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1404),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1421),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1390),
.B(n_1373),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1393),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1393),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1396),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1396),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1399),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1389),
.B(n_1358),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1394),
.B(n_1358),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1394),
.B(n_1358),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1399),
.B(n_1358),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1410),
.B(n_1357),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1404),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1416),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1398),
.B(n_1356),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1398),
.B(n_1400),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1422),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1400),
.B(n_1356),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1411),
.B(n_1382),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1440),
.Y(n_1462)
);

INVxp67_ASAP7_75t_L g1463 ( 
.A(n_1452),
.Y(n_1463)
);

AOI211xp5_ASAP7_75t_L g1464 ( 
.A1(n_1428),
.A2(n_1395),
.B(n_1387),
.C(n_1397),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1436),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1454),
.B(n_1418),
.Y(n_1466)
);

AOI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1428),
.A2(n_1395),
.B1(n_1401),
.B2(n_1406),
.Y(n_1467)
);

NAND4xp25_ASAP7_75t_L g1468 ( 
.A(n_1430),
.B(n_1401),
.C(n_1406),
.D(n_1405),
.Y(n_1468)
);

INVx1_ASAP7_75t_SL g1469 ( 
.A(n_1454),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1433),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1432),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1418),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1433),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1438),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1438),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1441),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1458),
.B(n_1391),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1445),
.B(n_1412),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1458),
.B(n_1391),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1446),
.B(n_1392),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1443),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1459),
.B(n_1420),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1443),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1469),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1468),
.B(n_1388),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1463),
.B(n_1459),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1461),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1459),
.Y(n_1490)
);

INVxp67_ASAP7_75t_L g1491 ( 
.A(n_1467),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1461),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1467),
.B(n_1464),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1469),
.B(n_1434),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1470),
.Y(n_1495)
);

INVxp67_ASAP7_75t_SL g1496 ( 
.A(n_1473),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1470),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1468),
.B(n_1426),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.B(n_1456),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1474),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1474),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1464),
.A2(n_1414),
.B1(n_1408),
.B2(n_1430),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1471),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1475),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1466),
.B(n_1456),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1472),
.B(n_1456),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1481),
.B(n_1435),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1483),
.B(n_1460),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1472),
.B(n_1455),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1482),
.B(n_1460),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1481),
.B(n_1435),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1471),
.B(n_1455),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1475),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1476),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1482),
.B(n_1434),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1476),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1473),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1434),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1479),
.B(n_1446),
.Y(n_1520)
);

OAI211xp5_ASAP7_75t_L g1521 ( 
.A1(n_1479),
.A2(n_1426),
.B(n_1423),
.C(n_1448),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1461),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1484),
.B(n_1442),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1442),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1471),
.B(n_1442),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1485),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1462),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1486),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1500),
.B(n_1506),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1500),
.B(n_1477),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1491),
.B(n_1477),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1486),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1488),
.B(n_1452),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1504),
.Y(n_1535)
);

NOR2xp33_ASAP7_75t_L g1536 ( 
.A(n_1493),
.B(n_1261),
.Y(n_1536)
);

NAND2x1p5_ASAP7_75t_L g1537 ( 
.A(n_1494),
.B(n_1372),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1494),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1494),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1497),
.Y(n_1540)
);

OR2x2_ASAP7_75t_L g1541 ( 
.A(n_1488),
.B(n_1437),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1501),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1490),
.B(n_1437),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1503),
.A2(n_1451),
.B1(n_1448),
.B2(n_1337),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1525),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1502),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1504),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1498),
.B(n_1409),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1525),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1514),
.Y(n_1551)
);

NOR2x1_ASAP7_75t_L g1552 ( 
.A(n_1487),
.B(n_1465),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1504),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1506),
.B(n_1478),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1515),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1508),
.A2(n_1415),
.B1(n_1337),
.B2(n_1448),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1518),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1525),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1517),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1490),
.B(n_1447),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1512),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1507),
.B(n_1478),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1539),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1561),
.B(n_1496),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1555),
.Y(n_1565)
);

INVx2_ASAP7_75t_SL g1566 ( 
.A(n_1528),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1558),
.B(n_1507),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1528),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1557),
.A2(n_1509),
.B1(n_1499),
.B2(n_1451),
.Y(n_1569)
);

OAI22xp5_ASAP7_75t_L g1570 ( 
.A1(n_1552),
.A2(n_1521),
.B1(n_1510),
.B2(n_1451),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1558),
.B(n_1510),
.Y(n_1571)
);

OAI332xp33_ASAP7_75t_L g1572 ( 
.A1(n_1532),
.A2(n_1523),
.A3(n_1516),
.B1(n_1524),
.B2(n_1519),
.B3(n_1499),
.C1(n_1509),
.C2(n_1526),
.Y(n_1572)
);

OAI33xp33_ASAP7_75t_L g1573 ( 
.A1(n_1532),
.A2(n_1511),
.A3(n_1524),
.B1(n_1523),
.B2(n_1516),
.B3(n_1519),
.Y(n_1573)
);

INVxp67_ASAP7_75t_SL g1574 ( 
.A(n_1528),
.Y(n_1574)
);

OAI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1549),
.A2(n_1520),
.B(n_1511),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1557),
.B(n_1489),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1533),
.A2(n_1513),
.B(n_1522),
.C(n_1527),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1533),
.A2(n_1513),
.B(n_1413),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1552),
.B(n_1492),
.C(n_1489),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1545),
.Y(n_1580)
);

AOI322xp5_ASAP7_75t_L g1581 ( 
.A1(n_1556),
.A2(n_1439),
.A3(n_1431),
.B1(n_1457),
.B2(n_1453),
.C1(n_1449),
.C2(n_1450),
.Y(n_1581)
);

NOR2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1533),
.B(n_1348),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1544),
.A2(n_1536),
.B1(n_1538),
.B2(n_1550),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_L g1584 ( 
.A1(n_1544),
.A2(n_1538),
.B(n_1550),
.Y(n_1584)
);

OAI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1545),
.A2(n_1369),
.B1(n_1380),
.B2(n_1429),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1545),
.B(n_1480),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1574),
.B(n_1538),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1571),
.B(n_1545),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1563),
.B(n_1534),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1529),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1570),
.B(n_1550),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1566),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1568),
.B(n_1529),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1566),
.B(n_1554),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1567),
.B(n_1554),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1580),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1565),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1567),
.B(n_1530),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1580),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1587),
.B(n_1530),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1576),
.B(n_1534),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1587),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1586),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1564),
.B(n_1562),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1576),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1592),
.A2(n_1572),
.B(n_1575),
.Y(n_1608)
);

OAI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1607),
.A2(n_1579),
.B1(n_1584),
.B2(n_1569),
.Y(n_1609)
);

NAND3xp33_ASAP7_75t_L g1610 ( 
.A(n_1593),
.B(n_1583),
.C(n_1577),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1606),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1594),
.A2(n_1605),
.B(n_1588),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1599),
.B(n_1582),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1595),
.B(n_1573),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1606),
.Y(n_1616)
);

AOI22xp5_ASAP7_75t_SL g1617 ( 
.A1(n_1589),
.A2(n_1597),
.B1(n_1603),
.B2(n_1591),
.Y(n_1617)
);

AOI321xp33_ASAP7_75t_L g1618 ( 
.A1(n_1591),
.A2(n_1540),
.A3(n_1551),
.B1(n_1542),
.B2(n_1546),
.C(n_1559),
.Y(n_1618)
);

OAI211xp5_ASAP7_75t_L g1619 ( 
.A1(n_1608),
.A2(n_1604),
.B(n_1598),
.C(n_1590),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1617),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1609),
.B(n_1598),
.C(n_1603),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1615),
.B(n_1596),
.C(n_1590),
.D(n_1589),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1612),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1614),
.Y(n_1624)
);

INVxp33_ASAP7_75t_L g1625 ( 
.A(n_1611),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1613),
.B(n_1602),
.Y(n_1626)
);

INVx2_ASAP7_75t_SL g1627 ( 
.A(n_1616),
.Y(n_1627)
);

AOI221xp5_ASAP7_75t_L g1628 ( 
.A1(n_1621),
.A2(n_1609),
.B1(n_1610),
.B2(n_1597),
.C(n_1601),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_L g1629 ( 
.A(n_1625),
.B(n_1602),
.Y(n_1629)
);

NOR3xp33_ASAP7_75t_L g1630 ( 
.A(n_1626),
.B(n_1600),
.C(n_1601),
.Y(n_1630)
);

AOI211xp5_ASAP7_75t_L g1631 ( 
.A1(n_1619),
.A2(n_1600),
.B(n_1553),
.C(n_1618),
.Y(n_1631)
);

O2A1O1Ixp33_ASAP7_75t_L g1632 ( 
.A1(n_1620),
.A2(n_1627),
.B(n_1622),
.C(n_1624),
.Y(n_1632)
);

NOR2x1_ASAP7_75t_L g1633 ( 
.A(n_1629),
.B(n_1623),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1630),
.B(n_1553),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1632),
.B(n_1535),
.Y(n_1635)
);

NOR3xp33_ASAP7_75t_L g1636 ( 
.A(n_1628),
.B(n_1535),
.C(n_1547),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1631),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1632),
.Y(n_1638)
);

OAI211xp5_ASAP7_75t_L g1639 ( 
.A1(n_1636),
.A2(n_1581),
.B(n_1547),
.C(n_1531),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1638),
.B(n_1531),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1634),
.Y(n_1641)
);

OAI211xp5_ASAP7_75t_L g1642 ( 
.A1(n_1635),
.A2(n_1633),
.B(n_1637),
.C(n_1547),
.Y(n_1642)
);

NAND4xp75_ASAP7_75t_L g1643 ( 
.A(n_1635),
.B(n_1559),
.C(n_1540),
.D(n_1548),
.Y(n_1643)
);

NAND2x1_ASAP7_75t_L g1644 ( 
.A(n_1640),
.B(n_1542),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1641),
.B(n_1546),
.Y(n_1645)
);

XNOR2xp5_ASAP7_75t_L g1646 ( 
.A(n_1643),
.B(n_1548),
.Y(n_1646)
);

NAND4xp25_ASAP7_75t_L g1647 ( 
.A(n_1645),
.B(n_1642),
.C(n_1639),
.D(n_1551),
.Y(n_1647)
);

AOI211xp5_ASAP7_75t_L g1648 ( 
.A1(n_1647),
.A2(n_1646),
.B(n_1644),
.C(n_1585),
.Y(n_1648)
);

OAI21xp5_ASAP7_75t_L g1649 ( 
.A1(n_1648),
.A2(n_1537),
.B(n_1541),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1649),
.B(n_1541),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1650),
.A2(n_1522),
.B(n_1492),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1651),
.A2(n_1560),
.B(n_1543),
.Y(n_1652)
);

BUFx4_ASAP7_75t_R g1653 ( 
.A(n_1652),
.Y(n_1653)
);

XNOR2xp5_ASAP7_75t_L g1654 ( 
.A(n_1652),
.B(n_1348),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1537),
.B1(n_1543),
.B2(n_1560),
.C(n_1527),
.Y(n_1655)
);

AOI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1653),
.B(n_1348),
.C(n_1462),
.Y(n_1656)
);


endmodule