module fake_jpeg_20374_n_215 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_215);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_215;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_14),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_42),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_54),
.B1(n_36),
.B2(n_1),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_30),
.B1(n_17),
.B2(n_33),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_50),
.B1(n_58),
.B2(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_20),
.B1(n_31),
.B2(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_29),
.B1(n_32),
.B2(n_23),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_14),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_61),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_69),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_68),
.Y(n_77)
);

AO22x2_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_25),
.B1(n_28),
.B2(n_2),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_36),
.B(n_1),
.C(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_13),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_89),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_82),
.B(n_86),
.Y(n_110)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_76),
.A2(n_92),
.B1(n_84),
.B2(n_72),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_77),
.B(n_78),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_0),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_1),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_68),
.A2(n_67),
.B1(n_62),
.B2(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

OAI21xp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_2),
.B(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_4),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_4),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_91),
.A2(n_65),
.B1(n_46),
.B2(n_55),
.Y(n_102)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_96),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_49),
.B(n_5),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_57),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_93),
.B1(n_71),
.B2(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_47),
.B(n_8),
.Y(n_95)
);

OAI32xp33_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_99),
.A3(n_94),
.B1(n_98),
.B2(n_72),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_11),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_50),
.B(n_58),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_77),
.A2(n_52),
.B(n_67),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_73),
.B(n_85),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_104),
.B(n_120),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_57),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_106),
.B(n_112),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_99),
.A2(n_46),
.B1(n_82),
.B2(n_90),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_111),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_71),
.B1(n_91),
.B2(n_93),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_87),
.C(n_88),
.Y(n_112)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_113),
.A2(n_70),
.B1(n_81),
.B2(n_80),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_75),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_74),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_83),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_107),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_127),
.A2(n_139),
.B(n_123),
.Y(n_161)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_132),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_131),
.Y(n_157)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_145),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_75),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_107),
.C(n_109),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_96),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_138),
.B(n_144),
.Y(n_162)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_118),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_142),
.Y(n_156)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_101),
.C(n_110),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_112),
.C(n_124),
.Y(n_159)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_116),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_131),
.A2(n_110),
.B(n_104),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_149),
.B(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_135),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_104),
.B(n_106),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_128),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_158),
.Y(n_170)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

OAI211xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_115),
.B(n_113),
.C(n_102),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_155),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_101),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_139),
.C(n_130),
.Y(n_176)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_111),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_163),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

HAxp5_ASAP7_75t_SL g168 ( 
.A(n_147),
.B(n_139),
.CON(n_168),
.SN(n_168)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_150),
.B1(n_126),
.B2(n_144),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_171),
.A2(n_176),
.B1(n_153),
.B2(n_142),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_143),
.C(n_125),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_174),
.B(n_177),
.C(n_148),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_164),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_126),
.C(n_137),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_152),
.C(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_187),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_161),
.B1(n_146),
.B2(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_169),
.A2(n_146),
.B1(n_150),
.B2(n_162),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_182),
.A2(n_170),
.B1(n_167),
.B2(n_172),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_156),
.C(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_188),
.B(n_182),
.Y(n_191)
);

HAxp5_ASAP7_75t_SL g190 ( 
.A(n_183),
.B(n_165),
.CON(n_190),
.SN(n_190)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_170),
.B(n_167),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_180),
.B1(n_185),
.B2(n_178),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_165),
.B1(n_166),
.B2(n_173),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_196),
.B(n_181),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_200),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_184),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_193),
.B(n_194),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_192),
.B(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_202),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_206),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_189),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_195),
.C(n_186),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_205),
.A2(n_193),
.B1(n_198),
.B2(n_132),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_208),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_210),
.B(n_203),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_213),
.B(n_209),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_211),
.Y(n_215)
);


endmodule