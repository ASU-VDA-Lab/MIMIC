module fake_jpeg_30536_n_54 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_18),
.B(n_9),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_0),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

FAx1_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_0),
.CI(n_1),
.CON(n_28),
.SN(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_20),
.B(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_25),
.B1(n_22),
.B2(n_21),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_17),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_42),
.B(n_45),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_28),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_5),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_44),
.A2(n_36),
.B1(n_6),
.B2(n_7),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

AOI31xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_8),
.A3(n_13),
.B(n_14),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_51),
.A2(n_49),
.B(n_16),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_15),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_50),
.B(n_48),
.Y(n_54)
);


endmodule