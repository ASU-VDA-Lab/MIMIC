module fake_ibex_418_n_1330 (n_151, n_147, n_85, n_251, n_167, n_128, n_253, n_208, n_234, n_84, n_64, n_244, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_205, n_204, n_139, n_247, n_274, n_55, n_130, n_275, n_63, n_98, n_129, n_161, n_237, n_29, n_143, n_106, n_177, n_203, n_148, n_2, n_76, n_233, n_267, n_268, n_8, n_118, n_224, n_273, n_183, n_245, n_67, n_229, n_9, n_209, n_164, n_38, n_198, n_264, n_124, n_37, n_256, n_110, n_193, n_47, n_169, n_108, n_217, n_10, n_82, n_21, n_263, n_27, n_165, n_242, n_278, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_255, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_262, n_162, n_13, n_180, n_194, n_122, n_223, n_116, n_240, n_61, n_201, n_249, n_282, n_14, n_0, n_239, n_94, n_134, n_12, n_266, n_42, n_77, n_112, n_257, n_150, n_88, n_133, n_44, n_142, n_51, n_226, n_46, n_258, n_80, n_172, n_215, n_250, n_279, n_49, n_40, n_66, n_17, n_74, n_90, n_235, n_176, n_58, n_192, n_43, n_140, n_216, n_22, n_136, n_261, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_206, n_221, n_166, n_195, n_163, n_212, n_26, n_188, n_200, n_114, n_199, n_236, n_281, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_260, n_99, n_280, n_269, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_252, n_141, n_18, n_89, n_83, n_32, n_53, n_222, n_107, n_115, n_149, n_186, n_227, n_50, n_11, n_248, n_92, n_144, n_170, n_213, n_254, n_101, n_190, n_113, n_138, n_270, n_230, n_96, n_185, n_271, n_241, n_68, n_117, n_214, n_238, n_79, n_81, n_265, n_35, n_159, n_202, n_231, n_158, n_211, n_218, n_259, n_132, n_174, n_276, n_277, n_210, n_157, n_219, n_160, n_220, n_225, n_184, n_272, n_246, n_31, n_56, n_23, n_146, n_232, n_91, n_207, n_54, n_243, n_19, n_228, n_1330);

input n_151;
input n_147;
input n_85;
input n_251;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_84;
input n_64;
input n_244;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_205;
input n_204;
input n_139;
input n_247;
input n_274;
input n_55;
input n_130;
input n_275;
input n_63;
input n_98;
input n_129;
input n_161;
input n_237;
input n_29;
input n_143;
input n_106;
input n_177;
input n_203;
input n_148;
input n_2;
input n_76;
input n_233;
input n_267;
input n_268;
input n_8;
input n_118;
input n_224;
input n_273;
input n_183;
input n_245;
input n_67;
input n_229;
input n_9;
input n_209;
input n_164;
input n_38;
input n_198;
input n_264;
input n_124;
input n_37;
input n_256;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_217;
input n_10;
input n_82;
input n_21;
input n_263;
input n_27;
input n_165;
input n_242;
input n_278;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_255;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_262;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_223;
input n_116;
input n_240;
input n_61;
input n_201;
input n_249;
input n_282;
input n_14;
input n_0;
input n_239;
input n_94;
input n_134;
input n_12;
input n_266;
input n_42;
input n_77;
input n_112;
input n_257;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_226;
input n_46;
input n_258;
input n_80;
input n_172;
input n_215;
input n_250;
input n_279;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_235;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_216;
input n_22;
input n_136;
input n_261;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_206;
input n_221;
input n_166;
input n_195;
input n_163;
input n_212;
input n_26;
input n_188;
input n_200;
input n_114;
input n_199;
input n_236;
input n_281;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_260;
input n_99;
input n_280;
input n_269;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_252;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_222;
input n_107;
input n_115;
input n_149;
input n_186;
input n_227;
input n_50;
input n_11;
input n_248;
input n_92;
input n_144;
input n_170;
input n_213;
input n_254;
input n_101;
input n_190;
input n_113;
input n_138;
input n_270;
input n_230;
input n_96;
input n_185;
input n_271;
input n_241;
input n_68;
input n_117;
input n_214;
input n_238;
input n_79;
input n_81;
input n_265;
input n_35;
input n_159;
input n_202;
input n_231;
input n_158;
input n_211;
input n_218;
input n_259;
input n_132;
input n_174;
input n_276;
input n_277;
input n_210;
input n_157;
input n_219;
input n_160;
input n_220;
input n_225;
input n_184;
input n_272;
input n_246;
input n_31;
input n_56;
input n_23;
input n_146;
input n_232;
input n_91;
input n_207;
input n_54;
input n_243;
input n_19;
input n_228;

output n_1330;

wire n_1084;
wire n_1295;
wire n_507;
wire n_992;
wire n_766;
wire n_1110;
wire n_309;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_773;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_957;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_312;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_457;
wire n_494;
wire n_930;
wire n_1044;
wire n_1134;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_829;
wire n_825;
wire n_939;
wire n_655;
wire n_306;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_496;
wire n_434;
wire n_1258;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_518;
wire n_852;
wire n_1133;
wire n_904;
wire n_355;
wire n_646;
wire n_448;
wire n_466;
wire n_1030;
wire n_1094;
wire n_715;
wire n_530;
wire n_1214;
wire n_1274;
wire n_420;
wire n_769;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1071;
wire n_793;
wire n_937;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1215;
wire n_629;
wire n_573;
wire n_359;
wire n_433;
wire n_439;
wire n_1007;
wire n_643;
wire n_1276;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_369;
wire n_1301;
wire n_869;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_307;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_564;
wire n_562;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_308;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_397;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_451;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_314;
wire n_563;
wire n_881;
wire n_734;
wire n_1073;
wire n_1108;
wire n_382;
wire n_1239;
wire n_1209;
wire n_288;
wire n_379;
wire n_551;
wire n_729;
wire n_603;
wire n_422;
wire n_324;
wire n_391;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_544;
wire n_1281;
wire n_695;
wire n_639;
wire n_482;
wire n_870;
wire n_1298;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1154;
wire n_345;
wire n_455;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_462;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_823;
wire n_657;
wire n_1156;
wire n_1293;
wire n_749;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_583;
wire n_1015;
wire n_663;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1318;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_340;
wire n_1255;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_840;
wire n_1203;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1053;
wire n_1207;
wire n_310;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1210;
wire n_591;
wire n_1201;
wire n_1246;
wire n_732;
wire n_1236;
wire n_832;
wire n_316;
wire n_590;
wire n_325;
wire n_1184;
wire n_1013;
wire n_929;
wire n_315;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_944;
wire n_623;
wire n_585;
wire n_483;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_295;
wire n_1120;
wire n_576;
wire n_388;
wire n_1279;
wire n_290;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_429;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_413;
wire n_1069;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_696;
wire n_837;
wire n_640;
wire n_954;
wire n_363;
wire n_725;
wire n_596;
wire n_351;
wire n_456;
wire n_998;
wire n_1115;
wire n_801;
wire n_1046;
wire n_882;
wire n_942;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_444;
wire n_986;
wire n_495;
wire n_411;
wire n_927;
wire n_615;
wire n_803;
wire n_1087;
wire n_757;
wire n_712;
wire n_650;
wire n_409;
wire n_332;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_780;
wire n_502;
wire n_633;
wire n_532;
wire n_726;
wire n_863;
wire n_597;
wire n_285;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_291;
wire n_318;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_997;
wire n_891;
wire n_303;
wire n_717;
wire n_668;
wire n_871;
wire n_485;
wire n_1315;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1048;
wire n_774;
wire n_588;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1263;
wire n_443;
wire n_1185;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1163;
wire n_677;
wire n_964;
wire n_916;
wire n_503;
wire n_292;
wire n_895;
wire n_687;
wire n_1035;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1104;
wire n_1011;
wire n_529;
wire n_626;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_991;
wire n_961;
wire n_1223;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_423;
wire n_357;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_542;
wire n_1294;
wire n_900;
wire n_377;
wire n_647;
wire n_1291;
wire n_317;
wire n_326;
wire n_339;
wire n_348;
wire n_674;
wire n_287;
wire n_552;
wire n_1112;
wire n_1267;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_508;
wire n_453;
wire n_400;
wire n_1055;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_296;
wire n_690;
wire n_1225;
wire n_982;
wire n_785;
wire n_604;
wire n_977;
wire n_719;
wire n_370;
wire n_289;
wire n_716;
wire n_923;
wire n_642;
wire n_286;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1021;
wire n_746;
wire n_1188;
wire n_742;
wire n_1191;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1224;
wire n_356;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_922;
wire n_851;
wire n_993;
wire n_300;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_826;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_935;
wire n_925;
wire n_1054;
wire n_722;
wire n_804;
wire n_484;
wire n_480;
wire n_1057;
wire n_354;
wire n_516;
wire n_329;
wire n_1149;
wire n_1176;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1139;
wire n_1018;
wire n_858;
wire n_385;
wire n_1324;
wire n_782;
wire n_616;
wire n_833;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1221;
wire n_284;
wire n_1047;
wire n_792;
wire n_1314;
wire n_575;
wire n_313;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_513;
wire n_877;
wire n_311;
wire n_1088;
wire n_896;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_302;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_912;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_298;
wire n_1256;
wire n_587;
wire n_1303;
wire n_764;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_756;
wire n_1257;
wire n_387;
wire n_688;
wire n_946;
wire n_707;
wire n_1097;
wire n_293;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_586;
wire n_638;
wire n_304;
wire n_593;
wire n_1212;
wire n_1199;
wire n_478;
wire n_336;
wire n_861;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_828;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1098;
wire n_584;
wire n_1187;
wire n_698;
wire n_1061;
wire n_682;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1068;
wire n_617;
wire n_301;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1192;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1166;
wire n_758;
wire n_710;
wire n_720;
wire n_1023;
wire n_568;
wire n_813;
wire n_1211;
wire n_1284;
wire n_1116;
wire n_791;
wire n_543;
wire n_580;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1074;
wire n_759;
wire n_953;
wire n_1180;
wire n_536;
wire n_1220;
wire n_467;
wire n_427;
wire n_1262;
wire n_442;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_335;
wire n_966;
wire n_299;
wire n_949;
wire n_704;
wire n_924;
wire n_477;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_735;
wire n_305;
wire n_566;
wire n_581;
wire n_416;
wire n_1089;
wire n_392;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_658;
wire n_1216;
wire n_1026;
wire n_283;
wire n_366;
wire n_1033;
wire n_627;
wire n_990;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1002;
wire n_1111;
wire n_405;
wire n_1310;
wire n_612;
wire n_955;
wire n_440;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1145;
wire n_537;
wire n_1113;
wire n_913;
wire n_509;
wire n_1164;
wire n_1277;
wire n_1016;
wire n_680;
wire n_809;
wire n_856;
wire n_779;
wire n_294;
wire n_1280;
wire n_493;
wire n_519;
wire n_408;
wire n_361;
wire n_319;
wire n_1091;
wire n_1287;
wire n_860;
wire n_661;
wire n_848;
wire n_683;
wire n_1150;
wire n_1194;
wire n_620;
wire n_450;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_297;
wire n_921;
wire n_489;
wire n_908;
wire n_565;
wire n_1123;
wire n_1272;
wire n_984;
wire n_394;
wire n_364;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_265),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_264),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_120),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_213),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_258),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_208),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_274),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_18),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_75),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_234),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_211),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_110),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_135),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_129),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_100),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_192),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_140),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_245),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_187),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_88),
.Y(n_306)
);

BUFx2_ASAP7_75t_SL g307 ( 
.A(n_183),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_130),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_230),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_95),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_2),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_11),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_209),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_176),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_215),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_255),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_128),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_204),
.Y(n_318)
);

BUFx10_ASAP7_75t_L g319 ( 
.A(n_184),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_122),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_117),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_247),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_52),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_280),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_243),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_257),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_266),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_106),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_224),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_181),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_261),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_46),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_227),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_246),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_276),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_194),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_111),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_24),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_193),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_236),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_149),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_86),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_188),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_216),
.Y(n_345)
);

INVx2_ASAP7_75t_SL g346 ( 
.A(n_59),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_150),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_263),
.Y(n_348)
);

BUFx2_ASAP7_75t_SL g349 ( 
.A(n_101),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_207),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_152),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_219),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_268),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_32),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_269),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_199),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_254),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_38),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_157),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_271),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_242),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_267),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_186),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_190),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_50),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_9),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_37),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_218),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_93),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_248),
.Y(n_371)
);

BUFx10_ASAP7_75t_L g372 ( 
.A(n_273),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_49),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_156),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_175),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_136),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_231),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_191),
.Y(n_378)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_103),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_85),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_0),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_212),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_82),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_214),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_95),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_44),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_166),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_272),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_232),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_144),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_222),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_173),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_237),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_278),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_124),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_201),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_148),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_49),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_88),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_198),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_85),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_200),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_113),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_195),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_249),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_260),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_84),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_57),
.Y(n_408)
);

BUFx2_ASAP7_75t_L g409 ( 
.A(n_91),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_1),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_189),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_155),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_250),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_18),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_238),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_145),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_180),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_240),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_177),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_277),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_244),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_270),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_223),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_67),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_141),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_196),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_134),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_252),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_65),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_185),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_146),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_159),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_259),
.Y(n_433)
);

BUFx10_ASAP7_75t_L g434 ( 
.A(n_154),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_27),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_282),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_142),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_171),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_114),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_217),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_253),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_76),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_139),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_235),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_226),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_126),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_133),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_78),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_220),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_233),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_71),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_48),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_279),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_14),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_8),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_275),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_251),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_69),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_205),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_33),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_43),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_228),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_105),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_239),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_178),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_170),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_225),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_14),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_123),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_87),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_202),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_23),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_77),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_84),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_162),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_29),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_76),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_20),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_54),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_44),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_127),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_28),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_41),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_241),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_197),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_262),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_158),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_74),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_62),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_182),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_65),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_99),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_151),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_312),
.B(n_2),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_306),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_290),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_377),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_310),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_310),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_469),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_303),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_383),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_316),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_435),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_469),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_409),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_429),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_291),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_321),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_474),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_361),
.B(n_3),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_346),
.B(n_3),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_291),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_330),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_285),
.B(n_4),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_329),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_330),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_359),
.Y(n_520)
);

NOR2xp67_ASAP7_75t_L g521 ( 
.A(n_407),
.B(n_4),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_332),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_398),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_337),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_398),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_339),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_386),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_343),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_354),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_386),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_410),
.Y(n_532)
);

INVxp33_ASAP7_75t_SL g533 ( 
.A(n_293),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_374),
.Y(n_534)
);

INVxp33_ASAP7_75t_L g535 ( 
.A(n_399),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_410),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_370),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_283),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_414),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_382),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_443),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_288),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_309),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_475),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_460),
.Y(n_546)
);

INVxp67_ASAP7_75t_SL g547 ( 
.A(n_479),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_467),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_327),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_391),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_318),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_484),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_288),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_490),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_295),
.Y(n_555)
);

NOR2xp67_ASAP7_75t_L g556 ( 
.A(n_289),
.B(n_5),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_411),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_295),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_319),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_485),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_292),
.B(n_5),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_L g562 ( 
.A(n_296),
.B(n_6),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_394),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_319),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_394),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_502),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_499),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_504),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_500),
.B(n_501),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_527),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_507),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_551),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_551),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_505),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_564),
.B(n_292),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_533),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_538),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_551),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_526),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_510),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_511),
.Y(n_582)
);

CKINVDCx9p33_ASAP7_75t_R g583 ( 
.A(n_495),
.Y(n_583)
);

CKINVDCx8_ASAP7_75t_R g584 ( 
.A(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_529),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_538),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_549),
.B(n_395),
.Y(n_587)
);

INVx5_ASAP7_75t_L g588 ( 
.A(n_564),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_518),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_508),
.B(n_333),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_522),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_524),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_515),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_539),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_541),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_543),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_564),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_545),
.B(n_297),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_552),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_554),
.B(n_297),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_519),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_559),
.B(n_318),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_534),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_520),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_540),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_523),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_525),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_561),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_497),
.B(n_328),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_547),
.Y(n_613)
);

HB1xp67_ASAP7_75t_L g614 ( 
.A(n_544),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_556),
.B(n_395),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_513),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_514),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_498),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_535),
.B(n_311),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_546),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_562),
.B(n_328),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_521),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_SL g623 ( 
.A(n_550),
.B(n_406),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_548),
.Y(n_624)
);

BUFx6f_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_535),
.Y(n_626)
);

INVx6_ASAP7_75t_L g627 ( 
.A(n_509),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_560),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_563),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_506),
.B(n_301),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_512),
.B(n_319),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_503),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_503),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_565),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_542),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_542),
.B(n_307),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_553),
.Y(n_637)
);

AND2x2_ASAP7_75t_SL g638 ( 
.A(n_553),
.B(n_304),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_555),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_555),
.B(n_301),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_558),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_558),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_537),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_528),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_531),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_532),
.Y(n_646)
);

BUFx2_ASAP7_75t_L g647 ( 
.A(n_536),
.Y(n_647)
);

INVxp33_ASAP7_75t_SL g648 ( 
.A(n_527),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_502),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_502),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_499),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_564),
.B(n_372),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_499),
.B(n_347),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_499),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_R g655 ( 
.A(n_549),
.B(n_406),
.Y(n_655)
);

BUFx2_ASAP7_75t_L g656 ( 
.A(n_527),
.Y(n_656)
);

NOR2xp67_ASAP7_75t_L g657 ( 
.A(n_564),
.B(n_325),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_564),
.B(n_384),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_544),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_502),
.Y(n_661)
);

HB1xp67_ASAP7_75t_L g662 ( 
.A(n_527),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_499),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_551),
.Y(n_664)
);

CKINVDCx20_ASAP7_75t_R g665 ( 
.A(n_538),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_564),
.B(n_384),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_499),
.B(n_347),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_551),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_551),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_551),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_499),
.B(n_418),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_527),
.Y(n_672)
);

BUFx3_ASAP7_75t_L g673 ( 
.A(n_551),
.Y(n_673)
);

OAI21x1_ASAP7_75t_L g674 ( 
.A1(n_564),
.A2(n_465),
.B(n_418),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_505),
.B(n_333),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_499),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_323),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_538),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_499),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_499),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_502),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_538),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_499),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_419),
.Y(n_684)
);

INVx1_ASAP7_75t_SL g685 ( 
.A(n_527),
.Y(n_685)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_538),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_505),
.B(n_453),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_610),
.B(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_674),
.Y(n_689)
);

BUFx4f_ASAP7_75t_L g690 ( 
.A(n_625),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_594),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_616),
.B(n_372),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_567),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_598),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_685),
.B(n_367),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_572),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_619),
.B(n_284),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_572),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_575),
.B(n_453),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_673),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_581),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_599),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_588),
.Y(n_703)
);

BUFx8_ASAP7_75t_SL g704 ( 
.A(n_645),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_613),
.B(n_286),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_577),
.B(n_453),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_616),
.B(n_372),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_608),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_603),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_588),
.Y(n_710)
);

BUFx2_ASAP7_75t_L g711 ( 
.A(n_656),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_606),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_627),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_572),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_609),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_403),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_616),
.B(n_403),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_651),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_612),
.B(n_403),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_654),
.Y(n_721)
);

AND2x6_ASAP7_75t_L g722 ( 
.A(n_658),
.B(n_419),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_660),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_663),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_618),
.A2(n_416),
.B1(n_482),
.B2(n_422),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_658),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_612),
.B(n_434),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_584),
.Y(n_728)
);

INVx1_ASAP7_75t_SL g729 ( 
.A(n_577),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_666),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_676),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_611),
.B(n_416),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_643),
.Y(n_733)
);

OR2x6_ASAP7_75t_L g734 ( 
.A(n_636),
.B(n_349),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_612),
.B(n_434),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_664),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_677),
.B(n_287),
.Y(n_737)
);

BUFx4f_ASAP7_75t_L g738 ( 
.A(n_625),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_679),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_640),
.A2(n_482),
.B1(n_487),
.B2(n_422),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_611),
.B(n_487),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_666),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_580),
.A2(n_326),
.B1(n_345),
.B2(n_335),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_585),
.B(n_294),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_680),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_683),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_589),
.B(n_298),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_668),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_569),
.Y(n_749)
);

INVx1_ASAP7_75t_SL g750 ( 
.A(n_648),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_662),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_669),
.Y(n_752)
);

AND3x4_ASAP7_75t_L g753 ( 
.A(n_633),
.B(n_450),
.C(n_439),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_625),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_569),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_604),
.B(n_299),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_672),
.B(n_300),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_617),
.B(n_379),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_587),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_657),
.B(n_366),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_595),
.B(n_302),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_684),
.B(n_439),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_627),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_675),
.A2(n_373),
.B1(n_380),
.B2(n_368),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_576),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_576),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_653),
.Y(n_768)
);

INVx4_ASAP7_75t_L g769 ( 
.A(n_684),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_653),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_604),
.B(n_305),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_687),
.B(n_308),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_621),
.Y(n_773)
);

INVx6_ASAP7_75t_L g774 ( 
.A(n_659),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_640),
.B(n_614),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_566),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_596),
.B(n_313),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_622),
.B(n_621),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_628),
.B(n_381),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_591),
.B(n_385),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_667),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_597),
.A2(n_358),
.B1(n_363),
.B2(n_362),
.Y(n_782)
);

INVx5_ASAP7_75t_L g783 ( 
.A(n_573),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_667),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_601),
.A2(n_365),
.B1(n_388),
.B2(n_369),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_631),
.B(n_401),
.Y(n_786)
);

OR2x6_ASAP7_75t_L g787 ( 
.A(n_636),
.B(n_389),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_638),
.B(n_408),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_655),
.B(n_424),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_573),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_568),
.Y(n_791)
);

BUFx6f_ASAP7_75t_SL g792 ( 
.A(n_636),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_600),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_630),
.B(n_449),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_671),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_600),
.B(n_455),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_632),
.B(n_456),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_615),
.B(n_314),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_582),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_SL g800 ( 
.A(n_615),
.B(n_459),
.Y(n_800)
);

INVx5_ASAP7_75t_L g801 ( 
.A(n_574),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_579),
.Y(n_802)
);

OR2x2_ASAP7_75t_L g803 ( 
.A(n_644),
.B(n_461),
.Y(n_803)
);

AO21x2_ASAP7_75t_L g804 ( 
.A1(n_602),
.A2(n_396),
.B(n_390),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_642),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_579),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_634),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_583),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_641),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_637),
.B(n_466),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_639),
.B(n_315),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_623),
.B(n_320),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_629),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_590),
.B(n_462),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_641),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_592),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_593),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_641),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_639),
.Y(n_819)
);

AND2x4_ASAP7_75t_SL g820 ( 
.A(n_634),
.B(n_402),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_605),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_607),
.Y(n_822)
);

AND2x2_ASAP7_75t_SL g823 ( 
.A(n_647),
.B(n_417),
.Y(n_823)
);

INVxp67_ASAP7_75t_SL g824 ( 
.A(n_578),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_620),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_624),
.B(n_322),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_649),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_646),
.B(n_324),
.Y(n_828)
);

AND2x2_ASAP7_75t_SL g829 ( 
.A(n_650),
.B(n_420),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_661),
.Y(n_830)
);

OAI22xp33_ASAP7_75t_L g831 ( 
.A1(n_681),
.A2(n_477),
.B1(n_478),
.B2(n_471),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_635),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_586),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_665),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_678),
.B(n_331),
.Y(n_835)
);

NAND2x1p5_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_450),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_686),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_610),
.A2(n_421),
.B1(n_426),
.B2(n_425),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_626),
.Y(n_839)
);

AND2x4_ASAP7_75t_L g840 ( 
.A(n_626),
.B(n_480),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_610),
.B(n_334),
.Y(n_841)
);

AND2x2_ASAP7_75t_SL g842 ( 
.A(n_659),
.B(n_428),
.Y(n_842)
);

BUFx4f_ASAP7_75t_L g843 ( 
.A(n_625),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_674),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_685),
.B(n_481),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_626),
.B(n_483),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_570),
.Y(n_847)
);

INVx3_ASAP7_75t_L g848 ( 
.A(n_594),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_626),
.B(n_489),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_674),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_674),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_610),
.B(n_336),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_SL g853 ( 
.A1(n_645),
.A2(n_438),
.B1(n_445),
.B2(n_437),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_674),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_626),
.B(n_338),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_674),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_610),
.B(n_340),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_674),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_610),
.B(n_341),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_674),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_610),
.B(n_342),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_674),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_610),
.B(n_344),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_674),
.Y(n_864)
);

INVx2_ASAP7_75t_SL g865 ( 
.A(n_626),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

AND2x2_ASAP7_75t_SL g867 ( 
.A(n_659),
.B(n_446),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_844),
.A2(n_448),
.B(n_447),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_768),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_793),
.B(n_348),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_694),
.Y(n_871)
);

OAI22xp5_ASAP7_75t_L g872 ( 
.A1(n_766),
.A2(n_494),
.B1(n_457),
.B2(n_464),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_688),
.A2(n_451),
.B1(n_470),
.B2(n_468),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_751),
.B(n_729),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_770),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_749),
.A2(n_755),
.B1(n_767),
.B2(n_766),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_770),
.B(n_350),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_775),
.B(n_351),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_781),
.B(n_352),
.Y(n_879)
);

INVx2_ASAP7_75t_SL g880 ( 
.A(n_847),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_781),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_794),
.B(n_353),
.Y(n_882)
);

CKINVDCx20_ASAP7_75t_R g883 ( 
.A(n_704),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_784),
.B(n_355),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_794),
.B(n_356),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_784),
.A2(n_488),
.B1(n_491),
.B2(n_476),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_749),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_SL g888 ( 
.A(n_755),
.B(n_493),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_774),
.Y(n_889)
);

NOR3xp33_ASAP7_75t_L g890 ( 
.A(n_750),
.B(n_360),
.C(n_357),
.Y(n_890)
);

NAND2x1p5_ASAP7_75t_L g891 ( 
.A(n_711),
.B(n_6),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_734),
.B(n_7),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_800),
.B(n_364),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_774),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_795),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_695),
.B(n_7),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_796),
.B(n_865),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_839),
.A2(n_375),
.B1(n_376),
.B2(n_371),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_846),
.B(n_378),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_693),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_845),
.B(n_387),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_849),
.B(n_392),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_693),
.B(n_393),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_840),
.B(n_486),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_724),
.B(n_397),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_724),
.A2(n_10),
.B(n_8),
.C(n_9),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_746),
.B(n_400),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_709),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_746),
.B(n_404),
.Y(n_909)
);

BUFx3_ASAP7_75t_L g910 ( 
.A(n_764),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_852),
.B(n_859),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_712),
.B(n_715),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_717),
.B(n_405),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_734),
.B(n_10),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_841),
.B(n_412),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_732),
.B(n_12),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_719),
.B(n_413),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_721),
.A2(n_317),
.B1(n_423),
.B2(n_415),
.Y(n_918)
);

NAND4xp25_ASAP7_75t_SL g919 ( 
.A(n_725),
.B(n_827),
.C(n_788),
.D(n_706),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_701),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_723),
.B(n_427),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_740),
.A2(n_472),
.B1(n_431),
.B2(n_432),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_809),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_786),
.B(n_430),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_730),
.A2(n_317),
.B1(n_436),
.B2(n_433),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_857),
.B(n_861),
.Y(n_926)
);

BUFx8_ASAP7_75t_L g927 ( 
.A(n_792),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_731),
.B(n_440),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_863),
.B(n_463),
.Y(n_929)
);

NOR2x1_ASAP7_75t_R g930 ( 
.A(n_728),
.B(n_441),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_733),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_787),
.B(n_13),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_786),
.B(n_442),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_730),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_699),
.B(n_444),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_690),
.B(n_15),
.Y(n_936)
);

OR2x2_ASAP7_75t_L g937 ( 
.A(n_741),
.B(n_15),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_739),
.B(n_454),
.Y(n_938)
);

NAND3xp33_ASAP7_75t_L g939 ( 
.A(n_757),
.B(n_458),
.C(n_317),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_702),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_745),
.A2(n_317),
.B1(n_19),
.B2(n_16),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_737),
.B(n_17),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_838),
.B(n_17),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_708),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_787),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_780),
.B(n_21),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_753),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_947)
);

NOR2x1p5_ASAP7_75t_L g948 ( 
.A(n_776),
.B(n_25),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_691),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_822),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_713),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_726),
.B(n_25),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_726),
.B(n_26),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_765),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_691),
.Y(n_955)
);

INVxp67_ASAP7_75t_SL g956 ( 
.A(n_791),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_742),
.Y(n_957)
);

INVx8_ASAP7_75t_L g958 ( 
.A(n_792),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_742),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_779),
.B(n_29),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_772),
.B(n_30),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_769),
.B(n_31),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_848),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_33),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_773),
.B(n_34),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_689),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_773),
.B(n_34),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_797),
.B(n_35),
.Y(n_968)
);

AOI22xp5_ASAP7_75t_L g969 ( 
.A1(n_804),
.A2(n_37),
.B1(n_35),
.B2(n_36),
.Y(n_969)
);

INVx2_ASAP7_75t_SL g970 ( 
.A(n_818),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_799),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_722),
.B(n_36),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_803),
.B(n_39),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_763),
.B(n_40),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_705),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_815),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_763),
.B(n_697),
.Y(n_977)
);

NOR2xp67_ASAP7_75t_SL g978 ( 
.A(n_821),
.B(n_40),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_819),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_710),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_710),
.Y(n_981)
);

NOR2x1p5_ASAP7_75t_L g982 ( 
.A(n_816),
.B(n_42),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_850),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_761),
.B(n_42),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_761),
.B(n_43),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_805),
.B(n_45),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_754),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_756),
.B(n_45),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_771),
.B(n_46),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_744),
.B(n_47),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_851),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_853),
.A2(n_51),
.B1(n_47),
.B2(n_50),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_862),
.B(n_102),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_808),
.B(n_51),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_829),
.B(n_52),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_851),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_747),
.B(n_53),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_789),
.B(n_832),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_762),
.B(n_54),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_738),
.B(n_55),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_743),
.B(n_55),
.Y(n_1001)
);

AND2x6_ASAP7_75t_L g1002 ( 
.A(n_854),
.B(n_104),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_782),
.B(n_56),
.Y(n_1003)
);

AOI22x1_ASAP7_75t_L g1004 ( 
.A1(n_868),
.A2(n_856),
.B1(n_858),
.B2(n_854),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_876),
.A2(n_823),
.B1(n_867),
.B2(n_842),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_887),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_876),
.Y(n_1007)
);

NAND2x2_ASAP7_75t_L g1008 ( 
.A(n_948),
.B(n_817),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_919),
.A2(n_947),
.B1(n_998),
.B2(n_932),
.Y(n_1009)
);

AND2x4_ASAP7_75t_L g1010 ( 
.A(n_895),
.B(n_821),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_932),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_889),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_880),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_869),
.B(n_785),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_R g1015 ( 
.A(n_883),
.B(n_760),
.Y(n_1015)
);

OR2x4_ASAP7_75t_L g1016 ( 
.A(n_937),
.B(n_833),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_923),
.Y(n_1017)
);

INVxp67_ASAP7_75t_L g1018 ( 
.A(n_874),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_875),
.B(n_814),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_881),
.A2(n_813),
.B1(n_830),
.B2(n_825),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_894),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_912),
.Y(n_1022)
);

BUFx4f_ASAP7_75t_L g1023 ( 
.A(n_932),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_897),
.B(n_716),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_892),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_966),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_975),
.B(n_810),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_900),
.B(n_856),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_892),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_896),
.B(n_758),
.Y(n_1030)
);

AND3x1_ASAP7_75t_SL g1031 ( 
.A(n_982),
.B(n_834),
.C(n_824),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_950),
.B(n_837),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_873),
.B(n_855),
.Y(n_1033)
);

AND2x6_ASAP7_75t_L g1034 ( 
.A(n_914),
.B(n_858),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

INVx5_ASAP7_75t_L g1036 ( 
.A(n_892),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_908),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_920),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_940),
.Y(n_1039)
);

INVx2_ASAP7_75t_SL g1040 ( 
.A(n_958),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_924),
.B(n_933),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_983),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_956),
.B(n_818),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_R g1044 ( 
.A(n_931),
.B(n_843),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_991),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_916),
.B(n_818),
.Y(n_1046)
);

CKINVDCx6p67_ASAP7_75t_R g1047 ( 
.A(n_958),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_996),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_873),
.B(n_807),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_926),
.A2(n_864),
.B(n_860),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_944),
.Y(n_1051)
);

NOR3xp33_ASAP7_75t_SL g1052 ( 
.A(n_945),
.B(n_831),
.C(n_835),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_934),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_995),
.A2(n_820),
.B1(n_798),
.B2(n_828),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_911),
.B(n_692),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_979),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_971),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_949),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_955),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_968),
.B(n_707),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_878),
.B(n_718),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_952),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_973),
.B(n_720),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_891),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_946),
.B(n_811),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_976),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_930),
.Y(n_1067)
);

OR2x6_ASAP7_75t_L g1068 ( 
.A(n_958),
.B(n_836),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_953),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_927),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_957),
.B(n_703),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_872),
.B(n_727),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_959),
.B(n_703),
.Y(n_1073)
);

BUFx2_ASAP7_75t_L g1074 ( 
.A(n_930),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_962),
.Y(n_1075)
);

BUFx4_ASAP7_75t_SL g1076 ( 
.A(n_987),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_886),
.B(n_960),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_994),
.B(n_735),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_984),
.B(n_812),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_985),
.B(n_777),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_943),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1001),
.Y(n_1082)
);

NAND2xp33_ASAP7_75t_SL g1083 ( 
.A(n_978),
.B(n_826),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_SL g1084 ( 
.A(n_994),
.B(n_862),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_972),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_877),
.B(n_866),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_961),
.B(n_700),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_1003),
.Y(n_1088)
);

OR2x2_ASAP7_75t_SL g1089 ( 
.A(n_951),
.B(n_57),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_882),
.B(n_58),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_936),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_964),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_922),
.B(n_862),
.Y(n_1093)
);

INVx2_ASAP7_75t_SL g1094 ( 
.A(n_970),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_871),
.Y(n_1095)
);

BUFx5_ASAP7_75t_L g1096 ( 
.A(n_1002),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_992),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_899),
.B(n_58),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_965),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_967),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_941),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_988),
.B(n_866),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_992),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_974),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_954),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_1002),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_885),
.A2(n_748),
.B1(n_752),
.B2(n_736),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_870),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_879),
.B(n_759),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1086),
.A2(n_1065),
.B(n_1028),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1004),
.A2(n_1050),
.B(n_1086),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1028),
.A2(n_977),
.B(n_993),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_1005),
.B(n_941),
.C(n_890),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_1009),
.A2(n_906),
.B(n_942),
.C(n_989),
.Y(n_1114)
);

AOI21xp33_ASAP7_75t_L g1115 ( 
.A1(n_1041),
.A2(n_997),
.B(n_990),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1022),
.B(n_935),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1101),
.B(n_1009),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1005),
.B(n_986),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1026),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1105),
.B(n_1097),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1006),
.Y(n_1121)
);

AND2x2_ASAP7_75t_L g1122 ( 
.A(n_1023),
.B(n_902),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1007),
.B(n_904),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1027),
.A2(n_999),
.B(n_905),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_1036),
.B(n_980),
.Y(n_1125)
);

AO21x1_ASAP7_75t_L g1126 ( 
.A1(n_1093),
.A2(n_969),
.B(n_1000),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1102),
.A2(n_939),
.B(n_907),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_1042),
.A2(n_981),
.A3(n_903),
.B(n_909),
.Y(n_1128)
);

OAI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1033),
.A2(n_918),
.B(n_917),
.Y(n_1129)
);

OAI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1024),
.A2(n_918),
.B(n_913),
.Y(n_1130)
);

AND2x4_ASAP7_75t_L g1131 ( 
.A(n_1036),
.B(n_884),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1045),
.Y(n_1132)
);

BUFx3_ASAP7_75t_L g1133 ( 
.A(n_1047),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1103),
.A2(n_1049),
.B1(n_1077),
.B2(n_1011),
.Y(n_1134)
);

OR2x6_ASAP7_75t_L g1135 ( 
.A(n_1068),
.B(n_1070),
.Y(n_1135)
);

NAND3x1_ASAP7_75t_L g1136 ( 
.A(n_1089),
.B(n_1002),
.C(n_928),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_1076),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1055),
.A2(n_938),
.B(n_921),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1048),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1034),
.A2(n_901),
.B1(n_898),
.B2(n_888),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1099),
.A2(n_929),
.B(n_915),
.C(n_925),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1019),
.B(n_893),
.Y(n_1142)
);

BUFx2_ASAP7_75t_R g1143 ( 
.A(n_1008),
.Y(n_1143)
);

OAI21xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1062),
.A2(n_1002),
.B(n_963),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_1012),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1037),
.Y(n_1146)
);

AOI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1061),
.A2(n_1060),
.B(n_1063),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1066),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1014),
.B(n_60),
.Y(n_1149)
);

INVx4_ASAP7_75t_SL g1150 ( 
.A(n_1034),
.Y(n_1150)
);

NAND2x1p5_ASAP7_75t_L g1151 ( 
.A(n_1040),
.B(n_783),
.Y(n_1151)
);

AO31x2_ASAP7_75t_L g1152 ( 
.A1(n_1081),
.A2(n_698),
.A3(n_714),
.B(n_696),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_1034),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1052),
.B(n_61),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1063),
.A2(n_1079),
.B(n_1109),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1025),
.A2(n_801),
.B1(n_802),
.B2(n_790),
.Y(n_1156)
);

AO22x2_ASAP7_75t_L g1157 ( 
.A1(n_1091),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1056),
.Y(n_1158)
);

AND2x4_ASAP7_75t_L g1159 ( 
.A(n_1010),
.B(n_1034),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1030),
.A2(n_802),
.B(n_790),
.Y(n_1160)
);

AOI22x1_ASAP7_75t_L g1161 ( 
.A1(n_1082),
.A2(n_806),
.B1(n_108),
.B2(n_109),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_1106),
.B(n_1029),
.Y(n_1162)
);

OA21x2_ASAP7_75t_L g1163 ( 
.A1(n_1088),
.A2(n_112),
.B(n_107),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_1044),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_SL g1165 ( 
.A1(n_1096),
.A2(n_64),
.B(n_66),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1016),
.B(n_66),
.Y(n_1166)
);

INVx1_ASAP7_75t_SL g1167 ( 
.A(n_1145),
.Y(n_1167)
);

BUFx3_ASAP7_75t_L g1168 ( 
.A(n_1133),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1121),
.Y(n_1169)
);

BUFx4f_ASAP7_75t_L g1170 ( 
.A(n_1135),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1148),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1146),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1111),
.A2(n_1075),
.B(n_1069),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1126),
.A2(n_1100),
.A3(n_1092),
.B(n_1109),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_1147),
.A2(n_1032),
.B1(n_1020),
.B2(n_1108),
.C(n_1090),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1146),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_SL g1177 ( 
.A1(n_1134),
.A2(n_1096),
.B1(n_1106),
.B2(n_1064),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1155),
.A2(n_1084),
.B(n_1083),
.C(n_1039),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_1112),
.A2(n_1110),
.B(n_1117),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1158),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1150),
.B(n_1017),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1113),
.B(n_1118),
.Y(n_1182)
);

NAND2x1p5_ASAP7_75t_L g1183 ( 
.A(n_1153),
.B(n_1074),
.Y(n_1183)
);

OR2x2_ASAP7_75t_L g1184 ( 
.A(n_1119),
.B(n_1057),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1127),
.A2(n_1087),
.B(n_1085),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1137),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_1164),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1114),
.A2(n_1051),
.B(n_1038),
.C(n_1098),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1129),
.A2(n_1059),
.B(n_1058),
.C(n_1061),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_SL g1190 ( 
.A(n_1153),
.B(n_1135),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1132),
.B(n_1010),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1144),
.A2(n_1072),
.B(n_1080),
.C(n_1085),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1151),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1116),
.B(n_1013),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1115),
.A2(n_1078),
.B1(n_1096),
.B2(n_1046),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1143),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1159),
.B(n_1068),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1150),
.B(n_1043),
.Y(n_1198)
);

CKINVDCx11_ASAP7_75t_R g1199 ( 
.A(n_1159),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1179),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1182),
.A2(n_1157),
.B1(n_1154),
.B2(n_1166),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_L g1202 ( 
.A1(n_1182),
.A2(n_1157),
.B1(n_1130),
.B2(n_1120),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1179),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1184),
.B(n_1139),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1172),
.B(n_1123),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1176),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1194),
.B(n_1122),
.Y(n_1207)
);

INVx4_ASAP7_75t_L g1208 ( 
.A(n_1199),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1196),
.B(n_1067),
.C(n_1015),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1170),
.A2(n_1136),
.B1(n_1153),
.B2(n_1140),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1175),
.A2(n_1124),
.B1(n_1138),
.B2(n_1149),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1179),
.Y(n_1212)
);

OAI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1170),
.A2(n_1068),
.B1(n_1162),
.B2(n_1142),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1190),
.B(n_1152),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1199),
.A2(n_1165),
.B1(n_1131),
.B2(n_1096),
.Y(n_1215)
);

AND2x4_ASAP7_75t_L g1216 ( 
.A(n_1174),
.B(n_1152),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1173),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1192),
.A2(n_1141),
.A3(n_1156),
.B(n_1053),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1177),
.A2(n_1131),
.B1(n_1096),
.B2(n_1078),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1188),
.A2(n_1018),
.B(n_1054),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1177),
.A2(n_1125),
.B1(n_1046),
.B2(n_1104),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1214),
.Y(n_1222)
);

INVx4_ASAP7_75t_L g1223 ( 
.A(n_1208),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1207),
.B(n_1169),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1208),
.A2(n_1197),
.B1(n_1191),
.B2(n_1186),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1206),
.Y(n_1226)
);

OAI211xp5_ASAP7_75t_L g1227 ( 
.A1(n_1202),
.A2(n_1195),
.B(n_1187),
.C(n_1167),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1204),
.B(n_1171),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1205),
.B(n_1180),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1201),
.A2(n_1208),
.B1(n_1211),
.B2(n_1220),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1210),
.A2(n_1197),
.B1(n_1183),
.B2(n_1193),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_1209),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1211),
.A2(n_1195),
.B1(n_1197),
.B2(n_1104),
.Y(n_1233)
);

AOI221xp5_ASAP7_75t_L g1234 ( 
.A1(n_1213),
.A2(n_1188),
.B1(n_1189),
.B2(n_1094),
.C(n_1168),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_L g1235 ( 
.A1(n_1221),
.A2(n_1185),
.B1(n_1198),
.B2(n_1183),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1219),
.A2(n_1185),
.B1(n_1161),
.B2(n_1168),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1216),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_SL g1238 ( 
.A1(n_1216),
.A2(n_1181),
.B1(n_1043),
.B2(n_1163),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1215),
.A2(n_1181),
.B1(n_1173),
.B2(n_1160),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1222),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1222),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1226),
.Y(n_1242)
);

OAI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1223),
.A2(n_1163),
.B1(n_1203),
.B2(n_1200),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1224),
.Y(n_1244)
);

CKINVDCx14_ASAP7_75t_R g1245 ( 
.A(n_1223),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1237),
.B(n_1212),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1222),
.B(n_1212),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1228),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1222),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1229),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1225),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1239),
.B(n_1217),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1227),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1235),
.Y(n_1254)
);

OAI31xp33_ASAP7_75t_L g1255 ( 
.A1(n_1245),
.A2(n_1230),
.A3(n_1231),
.B(n_1235),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1244),
.B(n_1230),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1242),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1245),
.A2(n_1233),
.B1(n_1234),
.B2(n_1238),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1250),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1248),
.B(n_1217),
.Y(n_1260)
);

AOI221xp5_ASAP7_75t_L g1261 ( 
.A1(n_1253),
.A2(n_1232),
.B1(n_1236),
.B2(n_1178),
.C(n_1035),
.Y(n_1261)
);

AOI22xp5_ASAP7_75t_SL g1262 ( 
.A1(n_1251),
.A2(n_1031),
.B1(n_1173),
.B2(n_1021),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1254),
.A2(n_1073),
.B1(n_1071),
.B2(n_1095),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1257),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1255),
.B(n_1258),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1259),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1260),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1263),
.B(n_1252),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1262),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1263),
.Y(n_1270)
);

INVxp67_ASAP7_75t_L g1271 ( 
.A(n_1261),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1256),
.B(n_1246),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1270),
.B(n_1246),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1264),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1265),
.B(n_1240),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1274),
.Y(n_1276)
);

OR2x2_ASAP7_75t_L g1277 ( 
.A(n_1273),
.B(n_1267),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1276),
.A2(n_1265),
.B1(n_1275),
.B2(n_1269),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1278),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1279),
.B(n_1277),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1279),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1279),
.Y(n_1282)
);

AND4x1_ASAP7_75t_L g1283 ( 
.A(n_1281),
.B(n_1268),
.C(n_1271),
.D(n_1272),
.Y(n_1283)
);

NAND3xp33_ASAP7_75t_L g1284 ( 
.A(n_1282),
.B(n_1266),
.C(n_1107),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1280),
.Y(n_1285)
);

NOR3x1_ASAP7_75t_L g1286 ( 
.A(n_1281),
.B(n_1240),
.C(n_1241),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1282),
.A2(n_1249),
.B1(n_1247),
.B2(n_1243),
.Y(n_1287)
);

AO22x2_ASAP7_75t_L g1288 ( 
.A1(n_1284),
.A2(n_70),
.B1(n_67),
.B2(n_68),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1283),
.B(n_70),
.Y(n_1289)
);

NAND4xp25_ASAP7_75t_L g1290 ( 
.A(n_1286),
.B(n_75),
.C(n_72),
.D(n_73),
.Y(n_1290)
);

OAI211xp5_ASAP7_75t_SL g1291 ( 
.A1(n_1287),
.A2(n_79),
.B(n_80),
.C(n_81),
.Y(n_1291)
);

OAI21xp33_ASAP7_75t_L g1292 ( 
.A1(n_1285),
.A2(n_79),
.B(n_80),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_R g1293 ( 
.A(n_1289),
.B(n_83),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1288),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1290),
.B(n_89),
.Y(n_1295)
);

OAI211xp5_ASAP7_75t_L g1296 ( 
.A1(n_1291),
.A2(n_90),
.B(n_91),
.C(n_92),
.Y(n_1296)
);

XOR2xp5_ASAP7_75t_L g1297 ( 
.A(n_1290),
.B(n_94),
.Y(n_1297)
);

A2O1A1Ixp33_ASAP7_75t_L g1298 ( 
.A1(n_1292),
.A2(n_96),
.B(n_97),
.C(n_98),
.Y(n_1298)
);

AO22x1_ASAP7_75t_L g1299 ( 
.A1(n_1294),
.A2(n_1128),
.B1(n_1218),
.B2(n_1174),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1297),
.B(n_1174),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1293),
.Y(n_1301)
);

NOR3xp33_ASAP7_75t_L g1302 ( 
.A(n_1296),
.B(n_115),
.C(n_116),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1295),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1295),
.Y(n_1304)
);

O2A1O1Ixp33_ASAP7_75t_L g1305 ( 
.A1(n_1298),
.A2(n_118),
.B(n_119),
.C(n_121),
.Y(n_1305)
);

HB1xp67_ASAP7_75t_L g1306 ( 
.A(n_1303),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1304),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1301),
.Y(n_1308)
);

NAND4xp25_ASAP7_75t_L g1309 ( 
.A(n_1302),
.B(n_125),
.C(n_131),
.D(n_132),
.Y(n_1309)
);

NOR3xp33_ASAP7_75t_L g1310 ( 
.A(n_1305),
.B(n_137),
.C(n_138),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1306),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1308),
.Y(n_1312)
);

NOR2x1_ASAP7_75t_L g1313 ( 
.A(n_1307),
.B(n_1300),
.Y(n_1313)
);

OR3x1_ASAP7_75t_L g1314 ( 
.A(n_1309),
.B(n_1299),
.C(n_143),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1311),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1312),
.B(n_1310),
.C(n_147),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1314),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1313),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1315),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1317),
.A2(n_1318),
.B(n_1316),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1319),
.Y(n_1321)
);

INVxp67_ASAP7_75t_L g1322 ( 
.A(n_1320),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1321),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1322),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1323),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1324),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1326),
.B(n_281),
.Y(n_1327)
);

AOI322xp5_ASAP7_75t_L g1328 ( 
.A1(n_1325),
.A2(n_153),
.A3(n_160),
.B1(n_161),
.B2(n_163),
.C1(n_164),
.C2(n_165),
.Y(n_1328)
);

AOI221xp5_ASAP7_75t_L g1329 ( 
.A1(n_1327),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.C(n_172),
.Y(n_1329)
);

AOI211xp5_ASAP7_75t_L g1330 ( 
.A1(n_1329),
.A2(n_1328),
.B(n_174),
.C(n_179),
.Y(n_1330)
);


endmodule