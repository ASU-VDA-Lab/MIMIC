module fake_jpeg_21972_n_262 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_262);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_262;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_40),
.B(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_23),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_33),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_48),
.Y(n_81)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_41),
.A2(n_23),
.B1(n_31),
.B2(n_35),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_53),
.B1(n_60),
.B2(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_26),
.Y(n_51)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_61),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_23),
.B1(n_31),
.B2(n_48),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_26),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_54),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_57),
.A2(n_59),
.B1(n_68),
.B2(n_76),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_20),
.B1(n_32),
.B2(n_29),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_20),
.B1(n_36),
.B2(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_62),
.B(n_79),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_20),
.B(n_36),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_80),
.B(n_27),
.Y(n_110)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_65),
.Y(n_97)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_36),
.B1(n_26),
.B2(n_29),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_72),
.B(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_19),
.B1(n_28),
.B2(n_22),
.Y(n_73)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_16),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_46),
.A2(n_22),
.B1(n_19),
.B2(n_25),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_77),
.A2(n_83),
.B1(n_61),
.B2(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_78),
.Y(n_108)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_34),
.C(n_27),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_87),
.B(n_58),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_41),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_83)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_87),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_0),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_34),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_101),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_100),
.Y(n_124)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_96),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_24),
.B1(n_18),
.B2(n_71),
.Y(n_135)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_104),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_66),
.B(n_0),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_34),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_34),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_103),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_34),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_61),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_75),
.B(n_1),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_107),
.B(n_85),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_117),
.C(n_18),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_18),
.B(n_4),
.Y(n_137)
);

OR2x2_ASAP7_75t_SL g117 ( 
.A(n_65),
.B(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_121),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_137),
.B(n_91),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_111),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_79),
.C(n_62),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_138),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_56),
.B(n_67),
.C(n_85),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_126),
.B1(n_130),
.B2(n_93),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_125),
.B(n_132),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_82),
.B1(n_73),
.B2(n_70),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_69),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_129),
.C(n_98),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_58),
.C(n_64),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_96),
.A2(n_70),
.B1(n_74),
.B2(n_24),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_135),
.A2(n_146),
.B1(n_107),
.B2(n_95),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_2),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_8),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_18),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_142),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_116),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_140),
.Y(n_163)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_141),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_2),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_4),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_7),
.Y(n_165)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_105),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_108),
.B(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_145),
.B(n_147),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_108),
.B(n_5),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_144),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_SL g187 ( 
.A1(n_149),
.A2(n_155),
.B(n_169),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_150),
.A2(n_152),
.B1(n_160),
.B2(n_166),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_131),
.A2(n_94),
.B1(n_109),
.B2(n_117),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_120),
.B(n_128),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_157),
.A2(n_172),
.B(n_173),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_127),
.B(n_90),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_109),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_161),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_112),
.B1(n_115),
.B2(n_98),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_115),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_169),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_143),
.B1(n_139),
.B2(n_129),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_98),
.B1(n_10),
.B2(n_12),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_167),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_140),
.A2(n_123),
.B1(n_130),
.B2(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_121),
.A2(n_8),
.B(n_12),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_154),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_179),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_156),
.B(n_142),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_178),
.B(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_163),
.A2(n_141),
.B1(n_136),
.B2(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_181),
.A2(n_168),
.B(n_151),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_184),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_164),
.B(n_125),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_185),
.A2(n_194),
.B1(n_169),
.B2(n_162),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_136),
.B(n_14),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_188),
.A2(n_173),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_191),
.Y(n_206)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_124),
.C(n_13),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_185),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_195),
.A2(n_198),
.B(n_202),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_189),
.B(n_166),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_201),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g201 ( 
.A(n_189),
.B(n_158),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_174),
.B(n_157),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_172),
.C(n_155),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_207),
.Y(n_218)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_181),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_191),
.C(n_179),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_174),
.A2(n_149),
.B(n_160),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_152),
.B(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_209),
.B(n_170),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_198),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_186),
.B1(n_194),
.B2(n_182),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_214),
.A2(n_223),
.B(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_219),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_187),
.B1(n_186),
.B2(n_177),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_216),
.A2(n_222),
.B1(n_214),
.B2(n_225),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_222),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_165),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_181),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_171),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_229),
.B1(n_216),
.B2(n_219),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_199),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_236),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_206),
.B1(n_202),
.B2(n_196),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_195),
.B(n_210),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_237),
.B(n_188),
.Y(n_244)
);

XNOR2x1_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_236),
.Y(n_243)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_235),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_181),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_197),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_244),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_245),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_229),
.B(n_235),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_221),
.C(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_237),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_231),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_247),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_252),
.B(n_253),
.Y(n_257)
);

OAI21x1_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_243),
.B(n_233),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_255),
.A2(n_245),
.B(n_249),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_251),
.Y(n_256)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_256),
.Y(n_259)
);

AOI211xp5_ASAP7_75t_L g260 ( 
.A1(n_257),
.A2(n_258),
.B(n_226),
.C(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_228),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_259),
.Y(n_262)
);


endmodule