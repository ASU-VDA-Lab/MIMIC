module fake_jpeg_9511_n_329 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_329);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_329;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_46),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_45),
.A2(n_23),
.B1(n_20),
.B2(n_30),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_49),
.A2(n_27),
.B1(n_24),
.B2(n_38),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_44),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_50),
.B(n_55),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_52),
.A2(n_53),
.B1(n_64),
.B2(n_66),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_22),
.B1(n_30),
.B2(n_18),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_17),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_61),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_35),
.B1(n_27),
.B2(n_24),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_69),
.B1(n_71),
.B2(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_56),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_37),
.A2(n_17),
.B1(n_18),
.B2(n_33),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_37),
.A2(n_17),
.B1(n_33),
.B2(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_20),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_73),
.C(n_55),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_37),
.A2(n_34),
.B1(n_25),
.B2(n_23),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_42),
.A2(n_33),
.B1(n_32),
.B2(n_35),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_32),
.B1(n_24),
.B2(n_35),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_23),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_20),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_75),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_76),
.A2(n_80),
.B1(n_81),
.B2(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_42),
.B1(n_45),
.B2(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_88),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_107),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_51),
.A2(n_46),
.B1(n_41),
.B2(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_92),
.Y(n_124)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_41),
.B(n_36),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_108),
.B(n_31),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_91),
.B(n_95),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_51),
.A2(n_26),
.B1(n_19),
.B2(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_31),
.Y(n_93)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_31),
.Y(n_96)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_100),
.B(n_105),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_101),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_29),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_57),
.B1(n_61),
.B2(n_59),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_57),
.B(n_29),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_63),
.B(n_43),
.C(n_26),
.Y(n_107)
);

AO22x1_ASAP7_75t_SL g108 ( 
.A1(n_54),
.A2(n_43),
.B1(n_31),
.B2(n_3),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_48),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_57),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_72),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_113),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_60),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_119),
.B(n_76),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_96),
.A3(n_93),
.B1(n_82),
.B2(n_75),
.Y(n_119)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_126),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_60),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_43),
.Y(n_164)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_125),
.Y(n_146)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx13_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_135),
.Y(n_144)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_97),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_88),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_107),
.C(n_86),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_171),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_79),
.B(n_77),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_145),
.B(n_154),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_81),
.B(n_91),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_153),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_150),
.A2(n_160),
.B1(n_163),
.B2(n_136),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_130),
.B(n_106),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_128),
.A2(n_74),
.B1(n_108),
.B2(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OAI32xp33_ASAP7_75t_L g157 ( 
.A1(n_111),
.A2(n_106),
.A3(n_108),
.B1(n_92),
.B2(n_80),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_48),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_78),
.B(n_105),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_162),
.B1(n_159),
.B2(n_146),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_83),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_137),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_168),
.B1(n_170),
.B2(n_134),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_101),
.B(n_31),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_117),
.B(n_99),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_165),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_123),
.B(n_43),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_118),
.B(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_117),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_124),
.A2(n_84),
.B1(n_94),
.B2(n_99),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_169),
.A2(n_133),
.B1(n_94),
.B2(n_112),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_125),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_131),
.B(n_68),
.C(n_61),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_152),
.B(n_119),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_175),
.B(n_188),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_128),
.B1(n_131),
.B2(n_138),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_176),
.B(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_151),
.B(n_138),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_189),
.Y(n_215)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_124),
.B(n_115),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_180),
.A2(n_191),
.B1(n_200),
.B2(n_161),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_183),
.B(n_193),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_126),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_168),
.A2(n_127),
.B1(n_121),
.B2(n_125),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_185),
.A2(n_190),
.B1(n_194),
.B2(n_197),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_149),
.Y(n_186)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_187),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_98),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_151),
.B(n_133),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_127),
.B1(n_135),
.B2(n_84),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_167),
.B(n_68),
.Y(n_193)
);

OAI22x1_ASAP7_75t_L g233 ( 
.A1(n_195),
.A2(n_154),
.B1(n_169),
.B2(n_162),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_142),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_205),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_48),
.B1(n_134),
.B2(n_3),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_198),
.B(n_141),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_199),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_141),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_194),
.B1(n_160),
.B2(n_178),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_139),
.B(n_164),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_166),
.C(n_171),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_165),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_184),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_217),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_143),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_225),
.C(n_228),
.Y(n_238)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_226),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_192),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_170),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_158),
.B(n_145),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_233),
.B1(n_175),
.B2(n_173),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_221),
.B(n_173),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_230),
.Y(n_236)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_224),
.B(n_183),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_153),
.C(n_171),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_182),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_231),
.Y(n_255)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_237),
.B(n_247),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_181),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_240),
.C(n_243),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_172),
.C(n_193),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_181),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_251),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_188),
.C(n_197),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_246),
.B(n_249),
.C(n_254),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_202),
.B1(n_177),
.B2(n_188),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_248),
.A2(n_233),
.B1(n_211),
.B2(n_223),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_177),
.C(n_145),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_208),
.A2(n_154),
.B1(n_140),
.B2(n_148),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_232),
.A2(n_11),
.B(n_16),
.Y(n_251)
);

XOR2x2_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_140),
.Y(n_253)
);

OAI31xp33_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_212),
.A3(n_214),
.B(n_223),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_140),
.C(n_134),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_208),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_220),
.Y(n_260)
);

INVx11_ASAP7_75t_L g257 ( 
.A(n_253),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_267),
.B1(n_10),
.B2(n_15),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_258),
.A2(n_249),
.B1(n_235),
.B2(n_246),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_245),
.B(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_230),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_265),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_241),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_226),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_215),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_217),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_273),
.Y(n_290)
);

OAI222xp33_ASAP7_75t_L g272 ( 
.A1(n_247),
.A2(n_214),
.B1(n_224),
.B2(n_219),
.C1(n_206),
.C2(n_211),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_255),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_213),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_207),
.C(n_227),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_238),
.Y(n_282)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_277),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_270),
.B1(n_266),
.B2(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_243),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_282),
.C(n_286),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_254),
.B(n_251),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_266),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_237),
.B1(n_239),
.B2(n_240),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_284),
.A2(n_287),
.B1(n_289),
.B2(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_288),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_269),
.A2(n_262),
.B1(n_272),
.B2(n_264),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_226),
.Y(n_288)
);

OAI321xp33_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_267),
.A3(n_261),
.B1(n_259),
.B2(n_258),
.C(n_264),
.Y(n_291)
);

AOI21x1_ASAP7_75t_SL g304 ( 
.A1(n_291),
.A2(n_287),
.B(n_281),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_292),
.A2(n_13),
.B(n_15),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_293),
.A2(n_300),
.B(n_14),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_270),
.B1(n_263),
.B2(n_268),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_268),
.C(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_10),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_9),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_9),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_12),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_303),
.B(n_13),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_309),
.B(n_310),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_296),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_307),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_299),
.B(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_312),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_294),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_295),
.Y(n_318)
);

O2A1O1Ixp33_ASAP7_75t_SL g321 ( 
.A1(n_318),
.A2(n_319),
.B(n_312),
.C(n_292),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

OAI21xp33_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_323),
.B(n_315),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_320),
.A2(n_295),
.B1(n_14),
.B2(n_16),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_5),
.C(n_6),
.Y(n_326)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g323 ( 
.A1(n_316),
.A2(n_5),
.B(n_6),
.C(n_7),
.D(n_8),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_325),
.B(n_326),
.C(n_323),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_SL g328 ( 
.A1(n_327),
.A2(n_324),
.B(n_7),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_7),
.Y(n_329)
);


endmodule