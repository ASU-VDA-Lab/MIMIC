module fake_jpeg_1663_n_700 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_700);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_700;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_544;
wire n_455;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_588;
wire n_670;
wire n_168;
wire n_384;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVxp33_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_59),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_11),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_63),
.B(n_71),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_64),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_66),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_67),
.Y(n_161)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_68),
.Y(n_134)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_70),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_11),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_73),
.Y(n_195)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_74),
.Y(n_188)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx11_ASAP7_75t_L g229 ( 
.A(n_75),
.Y(n_229)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_76),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_40),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_82),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_34),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_83),
.Y(n_218)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_84),
.Y(n_227)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_20),
.Y(n_89)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_90),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_34),
.Y(n_91)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_91),
.Y(n_156)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_56),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g183 ( 
.A(n_94),
.Y(n_183)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_25),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_96),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_25),
.Y(n_97)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_97),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_98),
.Y(n_158)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_101),
.Y(n_168)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_46),
.Y(n_102)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_103),
.Y(n_208)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_104),
.Y(n_219)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx8_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_106),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_26),
.Y(n_108)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_43),
.B(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_117),
.Y(n_145)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_110),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_54),
.Y(n_111)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_111),
.Y(n_224)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_112),
.Y(n_231)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_26),
.Y(n_113)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_114),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_116),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_47),
.B(n_10),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_118),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_37),
.B(n_12),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_38),
.B(n_12),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_38),
.B(n_12),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_126),
.Y(n_146)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_131),
.Y(n_200)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

INVx6_ASAP7_75t_SL g126 ( 
.A(n_27),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_27),
.Y(n_127)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_127),
.Y(n_220)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_48),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_130),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_32),
.B(n_19),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_33),
.Y(n_132)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_48),
.B(n_8),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_50),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_71),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_147),
.B(n_206),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_50),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_148),
.B(n_171),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_22),
.B1(n_41),
.B2(n_39),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_150),
.A2(n_153),
.B1(n_164),
.B2(n_169),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_22),
.B1(n_41),
.B2(n_39),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_160),
.B(n_225),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_120),
.A2(n_41),
.B1(n_28),
.B2(n_39),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_117),
.A2(n_22),
.B1(n_28),
.B2(n_58),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_52),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_58),
.B1(n_28),
.B2(n_36),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_175),
.A2(n_184),
.B1(n_205),
.B2(n_209),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_90),
.B(n_44),
.C(n_55),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_198),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_96),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_180),
.B(n_187),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_123),
.A2(n_58),
.B1(n_55),
.B2(n_33),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_108),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_74),
.B(n_52),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_189),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_61),
.A2(n_36),
.B1(n_42),
.B2(n_21),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_193),
.A2(n_213),
.B1(n_100),
.B2(n_98),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_80),
.B(n_55),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_105),
.A2(n_42),
.B1(n_36),
.B2(n_44),
.Y(n_205)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_110),
.A2(n_45),
.B1(n_35),
.B2(n_24),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_65),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_66),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_212),
.B(n_216),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_67),
.A2(n_45),
.B1(n_35),
.B2(n_24),
.Y(n_213)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_87),
.B(n_24),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_64),
.A2(n_35),
.B1(n_21),
.B2(n_14),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_217),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_72),
.B(n_21),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_221),
.B(n_219),
.Y(n_316)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_73),
.Y(n_223)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_77),
.B(n_7),
.Y(n_225)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_83),
.Y(n_230)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_230),
.Y(n_254)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_88),
.Y(n_232)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_232),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_91),
.A2(n_115),
.B1(n_111),
.B2(n_106),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_234),
.A2(n_209),
.B1(n_150),
.B2(n_169),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_236),
.A2(n_267),
.B1(n_204),
.B2(n_218),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_222),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_237),
.B(n_239),
.Y(n_351)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_147),
.A2(n_85),
.B(n_13),
.C(n_15),
.Y(n_239)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_201),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_240),
.Y(n_369)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_241),
.Y(n_353)
);

INVx3_ASAP7_75t_SL g242 ( 
.A(n_226),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g380 ( 
.A(n_242),
.Y(n_380)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_243),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_0),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_244),
.B(n_268),
.Y(n_330)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_247),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_188),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_249),
.B(n_250),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_222),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_193),
.Y(n_251)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

AND2x4_ASAP7_75t_SL g252 ( 
.A(n_177),
.B(n_0),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g342 ( 
.A(n_252),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_139),
.A2(n_7),
.B1(n_18),
.B2(n_17),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_255),
.A2(n_290),
.B1(n_296),
.B2(n_309),
.Y(n_331)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_257),
.Y(n_375)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_259),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_188),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_260),
.B(n_271),
.Y(n_327)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_261),
.Y(n_348)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_136),
.Y(n_264)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_264),
.Y(n_332)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_173),
.Y(n_265)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_265),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_266),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_175),
.B(n_162),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_270),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_192),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_272),
.Y(n_386)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_273),
.Y(n_359)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_201),
.Y(n_275)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_275),
.Y(n_350)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_167),
.Y(n_277)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_277),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_192),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_278),
.B(n_293),
.Y(n_329)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g354 ( 
.A(n_279),
.Y(n_354)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_174),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_159),
.Y(n_281)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_281),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_164),
.A2(n_7),
.B(n_18),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_282),
.Y(n_335)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_283),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_228),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_284),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_153),
.A2(n_7),
.B(n_17),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_285),
.B(n_288),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_143),
.B(n_1),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_286),
.B(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_140),
.Y(n_287)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_287),
.Y(n_379)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_231),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_145),
.A2(n_5),
.B1(n_16),
.B2(n_13),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_146),
.A2(n_5),
.B1(n_19),
.B2(n_3),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_291),
.A2(n_297),
.B1(n_305),
.B2(n_315),
.Y(n_333)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_292),
.B(n_294),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_137),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_183),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_197),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_307),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_203),
.A2(n_234),
.B1(n_149),
.B2(n_214),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_199),
.A2(n_5),
.B1(n_19),
.B2(n_3),
.Y(n_297)
);

INVx3_ASAP7_75t_SL g298 ( 
.A(n_226),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_298),
.B(n_299),
.Y(n_366)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_138),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_141),
.B(n_1),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_168),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_301),
.B(n_306),
.Y(n_376)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_144),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_302),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_214),
.B(n_5),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_303),
.B(n_304),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_135),
.B(n_4),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_154),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_228),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_308),
.B(n_284),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_227),
.A2(n_2),
.B1(n_4),
.B2(n_155),
.Y(n_309)
);

BUFx2_ASAP7_75t_SL g310 ( 
.A(n_144),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g360 ( 
.A(n_310),
.Y(n_360)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_191),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_311),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_163),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_313),
.B(n_316),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_163),
.A2(n_229),
.B1(n_151),
.B2(n_134),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_220),
.A2(n_165),
.B1(n_185),
.B2(n_190),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_317),
.A2(n_161),
.B1(n_170),
.B2(n_172),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_210),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_319),
.Y(n_364)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_157),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_137),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_320),
.B(n_321),
.Y(n_365)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_196),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_156),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_322),
.B(n_264),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_259),
.A2(n_210),
.B1(n_208),
.B2(n_195),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_326),
.A2(n_313),
.B(n_242),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_261),
.A2(n_178),
.B1(n_156),
.B2(n_158),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_328),
.A2(n_346),
.B1(n_355),
.B2(n_358),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_155),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_339),
.B(n_373),
.C(n_374),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_L g341 ( 
.A1(n_263),
.A2(n_217),
.B(n_158),
.C(n_207),
.Y(n_341)
);

O2A1O1Ixp33_ASAP7_75t_L g423 ( 
.A1(n_341),
.A2(n_240),
.B(n_275),
.C(n_258),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_256),
.A2(n_224),
.B1(n_207),
.B2(n_178),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_352),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_256),
.A2(n_224),
.B1(n_170),
.B2(n_172),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_251),
.A2(n_161),
.B1(n_195),
.B2(n_204),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_361),
.A2(n_370),
.B1(n_252),
.B2(n_298),
.Y(n_403)
);

OAI32xp33_ASAP7_75t_L g367 ( 
.A1(n_253),
.A2(n_218),
.A3(n_251),
.B1(n_244),
.B2(n_286),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_367),
.B(n_239),
.Y(n_396)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_236),
.A2(n_282),
.B1(n_267),
.B2(n_274),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_312),
.B(n_238),
.C(n_300),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_245),
.B(n_248),
.C(n_299),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_276),
.B(n_283),
.C(n_281),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_377),
.B(n_374),
.C(n_371),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_382),
.Y(n_400)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_285),
.A2(n_262),
.B1(n_301),
.B2(n_292),
.Y(n_383)
);

OAI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_383),
.A2(n_326),
.B1(n_380),
.B2(n_337),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_361),
.A2(n_309),
.B1(n_290),
.B2(n_314),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_387),
.A2(n_390),
.B1(n_403),
.B2(n_406),
.Y(n_465)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_330),
.B(n_252),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_398),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_340),
.A2(n_306),
.B1(n_322),
.B2(n_302),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_338),
.B(n_330),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g452 ( 
.A(n_392),
.B(n_393),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_378),
.B(n_347),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_329),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_395),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_396),
.B(n_431),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_339),
.B(n_289),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_340),
.B(n_246),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_428),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_327),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_417),
.Y(n_440)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_402),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_265),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_410),
.Y(n_459)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_348),
.A2(n_334),
.B1(n_370),
.B2(n_335),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_362),
.Y(n_407)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_342),
.A2(n_308),
.B(n_243),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_408),
.A2(n_414),
.B(n_418),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_357),
.A2(n_241),
.B(n_247),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_409),
.A2(n_360),
.B(n_356),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_348),
.A2(n_288),
.B1(n_307),
.B2(n_272),
.Y(n_410)
);

BUFx2_ASAP7_75t_SL g412 ( 
.A(n_354),
.Y(n_412)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_412),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_373),
.B(n_235),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_413),
.B(n_419),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_235),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_415),
.B(n_420),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_354),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_351),
.A2(n_294),
.B(n_254),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_270),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_377),
.B(n_269),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_376),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_421),
.B(n_435),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_334),
.A2(n_254),
.B1(n_258),
.B2(n_257),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_422),
.A2(n_325),
.B1(n_337),
.B2(n_372),
.Y(n_457)
);

OAI22xp33_ASAP7_75t_SL g471 ( 
.A1(n_423),
.A2(n_434),
.B1(n_325),
.B2(n_380),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_424),
.B(n_381),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_L g425 ( 
.A1(n_357),
.A2(n_319),
.B(n_279),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_425),
.A2(n_409),
.B(n_408),
.Y(n_466)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g427 ( 
.A1(n_385),
.A2(n_311),
.B1(n_280),
.B2(n_321),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_427),
.Y(n_467)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_354),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_429),
.B(n_433),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_365),
.B(n_357),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_432),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_382),
.B(n_346),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_355),
.B(n_363),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_331),
.A2(n_341),
.B1(n_385),
.B2(n_333),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_366),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_366),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_437),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_364),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_399),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_444),
.B(n_445),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_399),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_399),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_446),
.B(n_447),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_399),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_363),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_411),
.C(n_389),
.Y(n_490)
);

NAND2x1_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_366),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_SL g514 ( 
.A1(n_456),
.A2(n_354),
.B(n_417),
.C(n_428),
.Y(n_514)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_390),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_458),
.B(n_460),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_400),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_415),
.A2(n_331),
.B1(n_358),
.B2(n_328),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_463),
.A2(n_475),
.B1(n_478),
.B2(n_394),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g488 ( 
.A1(n_466),
.A2(n_469),
.B(n_473),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_396),
.A2(n_336),
.B(n_359),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_379),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_470),
.B(n_481),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_471),
.A2(n_444),
.B1(n_445),
.B2(n_447),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_418),
.A2(n_343),
.B(n_356),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_403),
.A2(n_379),
.B1(n_359),
.B2(n_332),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_410),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_477),
.B(n_380),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_432),
.A2(n_386),
.B1(n_376),
.B2(n_375),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_479),
.A2(n_428),
.B(n_343),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_404),
.B(n_371),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_480),
.B(n_376),
.Y(n_513)
);

XOR2x2_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_398),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_482),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_462),
.A2(n_397),
.B1(n_420),
.B2(n_434),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_483),
.A2(n_494),
.B1(n_496),
.B2(n_498),
.Y(n_547)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_442),
.Y(n_485)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_485),
.Y(n_541)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_487),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_439),
.B(n_411),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_489),
.B(n_454),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_490),
.B(n_461),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_443),
.B(n_429),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_491),
.B(n_492),
.C(n_497),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_443),
.B(n_413),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_462),
.A2(n_397),
.B1(n_416),
.B2(n_433),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_450),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_495),
.B(n_450),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_465),
.A2(n_433),
.B1(n_406),
.B2(n_387),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_439),
.B(n_389),
.C(n_395),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_465),
.A2(n_391),
.B1(n_421),
.B2(n_419),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_452),
.A2(n_393),
.B1(n_391),
.B2(n_407),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_499),
.A2(n_500),
.B1(n_507),
.B2(n_509),
.Y(n_531)
);

AOI22x1_ASAP7_75t_L g500 ( 
.A1(n_471),
.A2(n_423),
.B1(n_414),
.B2(n_436),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_451),
.Y(n_501)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_501),
.Y(n_554)
);

A2O1A1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_469),
.A2(n_423),
.B(n_405),
.C(n_426),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_502),
.B(n_513),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_439),
.B(n_435),
.C(n_402),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_508),
.C(n_510),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_448),
.B(n_456),
.C(n_468),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_463),
.A2(n_422),
.B1(n_388),
.B2(n_386),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_448),
.B(n_372),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_438),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_511),
.Y(n_539)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_459),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_512),
.A2(n_516),
.B1(n_517),
.B2(n_521),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_514),
.A2(n_519),
.B(n_472),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_456),
.B(n_343),
.C(n_369),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_472),
.C(n_466),
.Y(n_529)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_459),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_518),
.A2(n_472),
.B1(n_479),
.B2(n_453),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_SL g520 ( 
.A(n_468),
.B(n_412),
.C(n_350),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_SL g530 ( 
.A(n_520),
.B(n_472),
.Y(n_530)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_438),
.Y(n_521)
);

NOR2x1_ASAP7_75t_R g522 ( 
.A(n_449),
.B(n_381),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_522),
.B(n_514),
.Y(n_560)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_497),
.B(n_452),
.C(n_470),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_523),
.B(n_530),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_524),
.B(n_529),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_507),
.A2(n_474),
.B1(n_458),
.B2(n_477),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_527),
.A2(n_536),
.B1(n_502),
.B2(n_517),
.Y(n_562)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_532),
.B(n_537),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_461),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_533),
.B(n_535),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_484),
.A2(n_474),
.B1(n_460),
.B2(n_446),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_505),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_537),
.B(n_549),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_489),
.B(n_456),
.C(n_449),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_538),
.B(n_558),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g540 ( 
.A1(n_484),
.A2(n_440),
.B1(n_454),
.B2(n_450),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_540),
.A2(n_551),
.B1(n_556),
.B2(n_561),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_482),
.B(n_440),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_542),
.B(n_508),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g543 ( 
.A1(n_488),
.A2(n_486),
.B(n_504),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g583 ( 
.A1(n_543),
.A2(n_544),
.B(n_546),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_492),
.B(n_441),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_SL g593 ( 
.A(n_545),
.B(n_457),
.Y(n_593)
);

CKINVDCx14_ASAP7_75t_R g591 ( 
.A(n_548),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_519),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_496),
.A2(n_475),
.B1(n_478),
.B2(n_480),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_490),
.B(n_481),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_553),
.B(n_522),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_488),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_518),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_483),
.A2(n_455),
.B1(n_453),
.B2(n_476),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_503),
.B(n_476),
.C(n_455),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_498),
.B(n_350),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g588 ( 
.A(n_559),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_560),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_509),
.A2(n_467),
.B1(n_473),
.B2(n_441),
.Y(n_561)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_562),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_531),
.A2(n_527),
.B1(n_494),
.B2(n_547),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_563),
.A2(n_569),
.B1(n_581),
.B2(n_594),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_547),
.A2(n_512),
.B1(n_515),
.B2(n_520),
.Y(n_569)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_571),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_590),
.Y(n_614)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_524),
.B(n_510),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_574),
.B(n_593),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_539),
.Y(n_575)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_575),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_543),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_576),
.B(n_578),
.Y(n_601)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g579 ( 
.A1(n_556),
.A2(n_500),
.B1(n_501),
.B2(n_485),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_579),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_551),
.A2(n_500),
.B1(n_521),
.B2(n_511),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_580),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_536),
.A2(n_560),
.B1(n_555),
.B2(n_557),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_558),
.B(n_345),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_582),
.B(n_585),
.Y(n_602)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_554),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_586),
.B(n_587),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_534),
.B(n_514),
.Y(n_587)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_554),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_589),
.B(n_552),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_526),
.B(n_514),
.Y(n_590)
);

CKINVDCx16_ASAP7_75t_R g592 ( 
.A(n_557),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_552),
.Y(n_605)
);

AOI211xp5_ASAP7_75t_L g594 ( 
.A1(n_549),
.A2(n_464),
.B(n_369),
.C(n_345),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_565),
.B(n_526),
.C(n_528),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_595),
.B(n_606),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_563),
.A2(n_525),
.B1(n_545),
.B2(n_544),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_603),
.A2(n_615),
.B1(n_566),
.B2(n_590),
.Y(n_625)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_605),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_591),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_565),
.B(n_528),
.C(n_535),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_607),
.B(n_609),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_567),
.B(n_568),
.C(n_572),
.Y(n_609)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_610),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_564),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_611),
.B(n_616),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_564),
.B(n_533),
.Y(n_612)
);

CKINVDCx14_ASAP7_75t_R g633 ( 
.A(n_612),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_562),
.A2(n_525),
.B1(n_550),
.B2(n_542),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_538),
.C(n_529),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_568),
.B(n_550),
.C(n_369),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_618),
.B(n_621),
.Y(n_640)
);

AO21x2_ASAP7_75t_L g620 ( 
.A1(n_587),
.A2(n_464),
.B(n_344),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_620),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_575),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_618),
.B(n_583),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_622),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_599),
.A2(n_569),
.B1(n_581),
.B2(n_570),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_624),
.A2(n_620),
.B1(n_613),
.B2(n_617),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_625),
.B(n_628),
.Y(n_648)
);

MAJx2_ASAP7_75t_L g626 ( 
.A(n_614),
.B(n_600),
.C(n_609),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_626),
.B(n_636),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_614),
.B(n_574),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_601),
.Y(n_630)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_630),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g631 ( 
.A1(n_601),
.A2(n_571),
.B(n_583),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_631),
.B(n_634),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_595),
.B(n_593),
.C(n_584),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_607),
.B(n_584),
.C(n_588),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_635),
.B(n_620),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g636 ( 
.A(n_615),
.B(n_594),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_600),
.B(n_573),
.Y(n_637)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_637),
.B(n_642),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_604),
.B(n_608),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_638),
.B(n_620),
.Y(n_653)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_608),
.A2(n_577),
.B(n_586),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g646 ( 
.A1(n_641),
.A2(n_604),
.B(n_610),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g642 ( 
.A(n_616),
.B(n_589),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_642),
.B(n_598),
.C(n_597),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_645),
.B(n_649),
.Y(n_673)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_646),
.Y(n_664)
);

OAI21xp5_ASAP7_75t_L g647 ( 
.A1(n_638),
.A2(n_598),
.B(n_596),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g675 ( 
.A1(n_647),
.A2(n_656),
.B(n_659),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_596),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g652 ( 
.A(n_622),
.B(n_603),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g670 ( 
.A(n_652),
.B(n_636),
.Y(n_670)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_SL g654 ( 
.A(n_629),
.B(n_602),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_654),
.B(n_655),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g655 ( 
.A(n_643),
.B(n_635),
.C(n_634),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_639),
.B(n_619),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_658),
.B(n_653),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_630),
.A2(n_620),
.B(n_613),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_SL g662 ( 
.A(n_661),
.B(n_638),
.Y(n_662)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_662),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_623),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_663),
.B(n_665),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_656),
.A2(n_627),
.B1(n_641),
.B2(n_633),
.Y(n_665)
);

XNOR2xp5_ASAP7_75t_SL g666 ( 
.A(n_652),
.B(n_625),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g679 ( 
.A(n_666),
.B(n_669),
.Y(n_679)
);

XNOR2xp5_ASAP7_75t_L g677 ( 
.A(n_667),
.B(n_670),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_657),
.B(n_626),
.C(n_628),
.Y(n_668)
);

NOR2xp67_ASAP7_75t_SL g685 ( 
.A(n_668),
.B(n_650),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_645),
.B(n_624),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_647),
.A2(n_646),
.B(n_659),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_671),
.A2(n_637),
.B(n_648),
.Y(n_682)
);

NAND3xp33_ASAP7_75t_SL g676 ( 
.A(n_675),
.B(n_660),
.C(n_658),
.Y(n_676)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_676),
.A2(n_682),
.B(n_683),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_SL g680 ( 
.A1(n_664),
.A2(n_651),
.B1(n_644),
.B2(n_640),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_680),
.B(n_681),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_673),
.B(n_648),
.Y(n_681)
);

AOI21x1_ASAP7_75t_L g683 ( 
.A1(n_672),
.A2(n_650),
.B(n_353),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_685),
.B(n_666),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_678),
.B(n_668),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g693 ( 
.A1(n_687),
.A2(n_688),
.B(n_690),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g688 ( 
.A1(n_679),
.A2(n_675),
.B(n_671),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_684),
.A2(n_674),
.B(n_670),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_691),
.B(n_689),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_686),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_692),
.B(n_694),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_693),
.A2(n_676),
.B(n_677),
.Y(n_696)
);

AO22x1_ASAP7_75t_L g697 ( 
.A1(n_696),
.A2(n_677),
.B1(n_667),
.B2(n_353),
.Y(n_697)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_697),
.B(n_695),
.C(n_344),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_698),
.A2(n_349),
.B(n_384),
.Y(n_699)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_699),
.B(n_349),
.C(n_384),
.Y(n_700)
);


endmodule