module fake_jpeg_1613_n_305 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_305);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_107;
wire n_39;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_282;
wire n_258;
wire n_96;

INVx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_33),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_43),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_47),
.Y(n_98)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_48),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

NAND2xp67_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_0),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_65),
.Y(n_92)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_59),
.Y(n_100)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_19),
.A2(n_0),
.B(n_1),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_5),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_62),
.B(n_68),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_71),
.Y(n_93)
);

AOI21xp33_ASAP7_75t_L g68 ( 
.A1(n_24),
.A2(n_1),
.B(n_2),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_25),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_70),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_1),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_107),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_27),
.C(n_42),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g135 ( 
.A(n_77),
.B(n_10),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_39),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_39),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_38),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g144 ( 
.A(n_85),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_46),
.A2(n_40),
.B1(n_20),
.B2(n_36),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_101),
.B1(n_103),
.B2(n_108),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_42),
.B1(n_41),
.B2(n_35),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_88),
.A2(n_92),
.B1(n_87),
.B2(n_106),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_55),
.B(n_38),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_89),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_20),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_57),
.B(n_36),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_52),
.B(n_41),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_60),
.A2(n_40),
.B1(n_35),
.B2(n_31),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_49),
.A2(n_30),
.B1(n_29),
.B2(n_26),
.Y(n_104)
);

AO22x1_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_26),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_58),
.B(n_4),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_50),
.B(n_5),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_111),
.B(n_10),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_67),
.B1(n_64),
.B2(n_63),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_53),
.B1(n_7),
.B2(n_8),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_142),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_72),
.Y(n_122)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_123),
.B(n_85),
.Y(n_160)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_134),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_137),
.Y(n_157)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_136),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_138),
.B(n_76),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_148),
.Y(n_153)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_L g142 ( 
.A1(n_101),
.A2(n_11),
.B1(n_13),
.B2(n_86),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_74),
.A2(n_77),
.B1(n_104),
.B2(n_72),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_143),
.A2(n_147),
.B1(n_109),
.B2(n_73),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_146),
.Y(n_152)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_109),
.A2(n_106),
.B1(n_87),
.B2(n_88),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_85),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_150),
.Y(n_161)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_73),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_156),
.B(n_160),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_159),
.B(n_169),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_100),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_84),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_114),
.B(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_168),
.B(n_174),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_139),
.A2(n_84),
.B1(n_91),
.B2(n_112),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_172),
.A2(n_146),
.B1(n_141),
.B2(n_118),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_115),
.B(n_112),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_144),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_102),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_132),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_177),
.B(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_102),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_180),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_124),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_158),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_128),
.C(n_144),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_127),
.C(n_170),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_129),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_SL g229 ( 
.A1(n_190),
.A2(n_192),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_182),
.A2(n_142),
.B1(n_137),
.B2(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_193),
.A2(n_198),
.B1(n_200),
.B2(n_175),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_161),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_201),
.Y(n_211)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_152),
.A2(n_136),
.B1(n_125),
.B2(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_202),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_157),
.A2(n_137),
.B1(n_122),
.B2(n_134),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_181),
.Y(n_203)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_155),
.B(n_165),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_166),
.B(n_149),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_172),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_171),
.A2(n_151),
.B(n_157),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_206),
.A2(n_169),
.B(n_160),
.Y(n_216)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_157),
.A3(n_173),
.B1(n_171),
.B2(n_162),
.C1(n_176),
.C2(n_151),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_202),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_206),
.A2(n_177),
.B(n_176),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

AOI21xp33_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_162),
.B(n_156),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_218),
.C(n_224),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_216),
.B(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

OA21x2_ASAP7_75t_L g220 ( 
.A1(n_190),
.A2(n_159),
.B(n_181),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_220),
.A2(n_229),
.B1(n_214),
.B2(n_207),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_221),
.A2(n_228),
.B1(n_207),
.B2(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_165),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_227),
.C(n_188),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_170),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_187),
.A2(n_170),
.B1(n_201),
.B2(n_193),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_239),
.C(n_251),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_236),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_213),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_185),
.C(n_186),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_211),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_219),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_243),
.A2(n_244),
.B1(n_246),
.B2(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_249),
.B(n_216),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_189),
.C(n_209),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_260),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_220),
.B1(n_231),
.B2(n_233),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_257),
.A2(n_232),
.B1(n_249),
.B2(n_230),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_233),
.Y(n_259)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_237),
.B(n_222),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_261),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_223),
.B(n_228),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_262),
.A2(n_238),
.B(n_221),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_217),
.C(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_239),
.C(n_184),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_251),
.Y(n_267)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_267),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_238),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_268),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_244),
.B1(n_220),
.B2(n_237),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_272),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_271),
.A2(n_253),
.B(n_261),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_264),
.C(n_265),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_203),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_254),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_250),
.B1(n_200),
.B2(n_183),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_259),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_277),
.A2(n_285),
.B(n_268),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_264),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_281),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_255),
.C(n_260),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_283),
.B(n_284),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_280),
.A2(n_268),
.B(n_269),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_292),
.B(n_285),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_276),
.B1(n_266),
.B2(n_275),
.Y(n_288)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_292),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_279),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_294),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_296),
.C(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_291),
.B(n_258),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_298),
.B(n_300),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_293),
.C(n_270),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_272),
.B(n_290),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_301),
.A2(n_271),
.B(n_199),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_302),
.B(n_196),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_304),
.B(n_208),
.Y(n_305)
);


endmodule