module fake_jpeg_13200_n_465 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_465);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_465;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_0),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g134 ( 
.A(n_50),
.Y(n_134)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_52),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_54),
.Y(n_123)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g150 ( 
.A(n_59),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_23),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_89),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_75),
.Y(n_98)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_28),
.Y(n_77)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_82),
.B(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_87),
.Y(n_99)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_92),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_16),
.B(n_0),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_96),
.Y(n_111)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_94),
.B(n_95),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_16),
.B(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_89),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_97),
.B(n_36),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_22),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_103),
.B(n_117),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_57),
.B1(n_90),
.B2(n_53),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_104),
.A2(n_106),
.B1(n_29),
.B2(n_37),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_58),
.A2(n_48),
.B1(n_32),
.B2(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_60),
.A2(n_17),
.B1(n_48),
.B2(n_32),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_110),
.A2(n_120),
.B1(n_141),
.B2(n_124),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_47),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_70),
.A2(n_17),
.B1(n_25),
.B2(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_47),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_129),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_45),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_36),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_143),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_88),
.A2(n_41),
.B1(n_43),
.B2(n_86),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_59),
.B(n_45),
.Y(n_143)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_152),
.Y(n_242)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_155),
.B(n_165),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_157),
.Y(n_234)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_160),
.Y(n_235)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_161),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_107),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_164),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_105),
.Y(n_167)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_149),
.A2(n_68),
.B1(n_80),
.B2(n_79),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_197),
.B1(n_199),
.B2(n_124),
.Y(n_209)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_22),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_180),
.Y(n_205)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g240 ( 
.A(n_173),
.B(n_176),
.Y(n_240)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_44),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_181),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_109),
.B(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_147),
.Y(n_178)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_179),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_111),
.B(n_44),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_102),
.B(n_23),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_182),
.Y(n_236)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_183),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_29),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_184),
.B(n_185),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_33),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_186),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_104),
.A2(n_85),
.B1(n_73),
.B2(n_65),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_189),
.B1(n_120),
.B2(n_148),
.Y(n_210)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_188),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_138),
.A2(n_62),
.B1(n_61),
.B2(n_33),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_211)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_128),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_191),
.Y(n_231)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_138),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_192),
.Y(n_233)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_112),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_114),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_134),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_196),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_241)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_141),
.A2(n_43),
.B1(n_41),
.B2(n_2),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_218),
.B1(n_222),
.B2(n_100),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_168),
.A2(n_134),
.B(n_142),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_159),
.B(n_133),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_148),
.B1(n_140),
.B2(n_145),
.Y(n_218)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_162),
.B(n_139),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_145),
.B1(n_121),
.B2(n_139),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_158),
.B(n_130),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_126),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_151),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_126),
.C(n_119),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_195),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_173),
.A2(n_115),
.B1(n_119),
.B2(n_43),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

AO21x1_ASAP7_75t_L g245 ( 
.A1(n_226),
.A2(n_181),
.B(n_166),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_245),
.A2(n_239),
.B(n_202),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_247),
.B(n_251),
.Y(n_303)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_214),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_209),
.A2(n_211),
.B1(n_216),
.B2(n_226),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_252),
.A2(n_255),
.B1(n_270),
.B2(n_271),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_253),
.A2(n_213),
.B1(n_236),
.B2(n_217),
.Y(n_287)
);

CKINVDCx6p67_ASAP7_75t_R g254 ( 
.A(n_223),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_254),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_226),
.A2(n_229),
.B1(n_232),
.B2(n_189),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_256),
.B(n_260),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_231),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_276),
.Y(n_285)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_223),
.B(n_176),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_174),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_261),
.B(n_263),
.Y(n_295)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_242),
.B(n_167),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_206),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_264),
.A2(n_274),
.B1(n_281),
.B2(n_243),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_232),
.A2(n_156),
.B1(n_115),
.B2(n_153),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_317)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_207),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_207),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_269),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_205),
.A2(n_198),
.B1(n_164),
.B2(n_163),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_205),
.A2(n_193),
.B1(n_182),
.B2(n_41),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_222),
.A2(n_41),
.B1(n_1),
.B2(n_2),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_272),
.A2(n_277),
.B1(n_243),
.B2(n_208),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_213),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_240),
.B(n_227),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_219),
.B(n_1),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_227),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_225),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_280),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

NOR2x1p5_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_3),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_218),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_213),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_282),
.B(n_235),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_219),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_283),
.B(n_289),
.C(n_307),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_299),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_287),
.A2(n_306),
.B1(n_309),
.B2(n_311),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_230),
.C(n_228),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_292),
.A2(n_275),
.B(n_261),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_253),
.A2(n_273),
.B1(n_248),
.B2(n_246),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_294),
.A2(n_298),
.B1(n_249),
.B2(n_206),
.Y(n_333)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_280),
.B(n_230),
.CI(n_228),
.CON(n_297),
.SN(n_297)
);

FAx1_ASAP7_75t_SL g345 ( 
.A(n_297),
.B(n_9),
.CI(n_10),
.CON(n_345),
.SN(n_345)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_246),
.A2(n_241),
.B1(n_203),
.B2(n_237),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_254),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_301),
.B1(n_264),
.B2(n_274),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_202),
.B(n_208),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_314),
.B(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_217),
.B1(n_237),
.B2(n_220),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_224),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_255),
.A2(n_224),
.B1(n_220),
.B2(n_221),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g343 ( 
.A(n_310),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_267),
.A2(n_270),
.B1(n_272),
.B2(n_271),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_257),
.A2(n_267),
.B1(n_276),
.B2(n_280),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_254),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_258),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_235),
.B(n_234),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_260),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_318),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_319),
.B(n_322),
.Y(n_353)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_320),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_298),
.A2(n_247),
.B1(n_256),
.B2(n_251),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_321),
.A2(n_333),
.B1(n_342),
.B2(n_347),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_303),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_304),
.A2(n_265),
.B1(n_259),
.B2(n_262),
.Y(n_323)
);

XOR2x1_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_326),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_263),
.Y(n_324)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_325),
.B(n_331),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_294),
.A2(n_254),
.B1(n_277),
.B2(n_250),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_327),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_288),
.B(n_278),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_329),
.B(n_346),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_269),
.C(n_268),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_336),
.C(n_344),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_303),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_332),
.A2(n_315),
.B1(n_287),
.B2(n_295),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_307),
.B(n_234),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_337),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_317),
.A2(n_221),
.B(n_274),
.Y(n_340)
);

AO22x1_ASAP7_75t_L g360 ( 
.A1(n_340),
.A2(n_341),
.B1(n_345),
.B2(n_284),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_317),
.A2(n_8),
.B(n_9),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_316),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_288),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_286),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_347)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_352),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_330),
.C(n_344),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_358),
.C(n_365),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_328),
.B(n_314),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_361),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_310),
.C(n_285),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_360),
.B(n_367),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_318),
.B(n_285),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_339),
.B(n_295),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_368),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_364),
.A2(n_348),
.B1(n_356),
.B2(n_351),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_291),
.C(n_286),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_322),
.B(n_302),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_291),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_331),
.B(n_290),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_370),
.B(n_347),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_334),
.A2(n_313),
.B1(n_311),
.B2(n_306),
.Y(n_371)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_371),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_354),
.A2(n_334),
.B1(n_343),
.B2(n_318),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_357),
.B(n_324),
.Y(n_375)
);

XNOR2x1_ASAP7_75t_L g411 ( 
.A(n_375),
.B(n_376),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_365),
.A2(n_333),
.B1(n_326),
.B2(n_346),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_353),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_383),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_338),
.C(n_335),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_379),
.B(n_384),
.C(n_389),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_369),
.A2(n_325),
.B(n_340),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_380),
.A2(n_394),
.B(n_371),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_351),
.A2(n_337),
.B1(n_327),
.B2(n_341),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_363),
.C(n_358),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_353),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_387),
.B(n_392),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_323),
.C(n_296),
.Y(n_389)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_297),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_373),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_356),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_345),
.Y(n_412)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_352),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_308),
.Y(n_396)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_396),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_377),
.B(n_348),
.C(n_361),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_406),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_403),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_379),
.B(n_359),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_400),
.B(n_381),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_384),
.B(n_373),
.C(n_372),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_405),
.C(n_394),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_350),
.B1(n_360),
.B2(n_312),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_309),
.C(n_312),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_388),
.C(n_391),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_308),
.C(n_342),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_409),
.B(n_380),
.C(n_390),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_300),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_410),
.B(n_412),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g413 ( 
.A(n_407),
.B(n_382),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_413),
.B(n_414),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_375),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_417),
.B(n_420),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_376),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_418),
.B(n_426),
.Y(n_438)
);

BUFx24_ASAP7_75t_SL g423 ( 
.A(n_402),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_423),
.B(n_424),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_374),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_425),
.B(n_397),
.C(n_409),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_386),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_438),
.C(n_428),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_408),
.C(n_411),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_431),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_422),
.A2(n_408),
.B1(n_420),
.B2(n_419),
.Y(n_430)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_430),
.Y(n_448)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_411),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_433),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_399),
.Y(n_433)
);

INVx13_ASAP7_75t_L g434 ( 
.A(n_426),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_437),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_421),
.A2(n_385),
.B1(n_416),
.B2(n_383),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_439),
.B(n_440),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_435),
.A2(n_385),
.B(n_345),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_297),
.C(n_13),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_442),
.B(n_444),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_297),
.C(n_13),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_12),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_14),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_14),
.Y(n_447)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_447),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_SL g449 ( 
.A1(n_445),
.A2(n_431),
.B(n_437),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_449),
.A2(n_452),
.B(n_443),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_436),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_454),
.B(n_430),
.Y(n_455)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_452),
.B(n_443),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_460),
.A2(n_457),
.B(n_459),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_453),
.B1(n_451),
.B2(n_458),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_441),
.C(n_432),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_441),
.C(n_433),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_464),
.B(n_434),
.Y(n_465)
);


endmodule