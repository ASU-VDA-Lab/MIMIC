module fake_netlist_5_2178_n_2936 (n_137, n_294, n_431, n_318, n_380, n_419, n_611, n_444, n_469, n_615, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_619, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_605, n_74, n_515, n_57, n_353, n_351, n_367, n_620, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_629, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_625, n_621, n_100, n_455, n_417, n_612, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_606, n_559, n_275, n_252, n_624, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_610, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_618, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_603, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_636, n_600, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_635, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_622, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_614, n_50, n_337, n_430, n_313, n_631, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_613, n_241, n_357, n_598, n_608, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_609, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_595, n_502, n_239, n_466, n_420, n_630, n_489, n_632, n_55, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_601, n_279, n_70, n_253, n_261, n_174, n_289, n_627, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_628, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_607, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_602, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_623, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_596, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_599, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_594, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_634, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_626, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2936);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_611;
input n_444;
input n_469;
input n_615;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_619;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_629;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_625;
input n_621;
input n_100;
input n_455;
input n_417;
input n_612;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_606;
input n_559;
input n_275;
input n_252;
input n_624;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_610;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_618;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_603;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_636;
input n_600;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_635;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_614;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_613;
input n_241;
input n_357;
input n_598;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_609;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_502;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_55;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_601;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_627;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_628;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_607;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_623;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_599;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_594;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_634;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_626;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2936;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_1462;
wire n_854;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1107;
wire n_1728;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_777;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1071;
wire n_1165;
wire n_1561;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2267;
wire n_2218;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2529;
wire n_2195;
wire n_2698;
wire n_809;
wire n_931;
wire n_870;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_744;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2320;
wire n_2038;
wire n_2473;
wire n_2137;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_968;
wire n_912;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_762;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_2935;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_990;
wire n_836;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_756;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_1546;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2335;
wire n_2135;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g637 ( 
.A(n_173),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_310),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_175),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_287),
.Y(n_640)
);

CKINVDCx20_ASAP7_75t_R g641 ( 
.A(n_588),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_337),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_219),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_429),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_288),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_102),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_224),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_562),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_221),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_417),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_249),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_113),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_526),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_205),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_107),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_563),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_283),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_237),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_403),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_272),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_482),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_602),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_528),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_474),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_440),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_630),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_438),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_442),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_93),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_108),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_614),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_324),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_623),
.Y(n_673)
);

BUFx5_ASAP7_75t_L g674 ( 
.A(n_349),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_235),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_414),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_295),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_162),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_351),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_247),
.Y(n_680)
);

CKINVDCx16_ASAP7_75t_R g681 ( 
.A(n_384),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_550),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_296),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_106),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_510),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_288),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_431),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_400),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_436),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g690 ( 
.A(n_31),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_308),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_120),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_610),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_469),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_227),
.Y(n_695)
);

CKINVDCx20_ASAP7_75t_R g696 ( 
.A(n_179),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_87),
.Y(n_697)
);

BUFx2_ASAP7_75t_L g698 ( 
.A(n_14),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_421),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_22),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_99),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_603),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_422),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_397),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_478),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_8),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_406),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_216),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_226),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_308),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_572),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_155),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_565),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_552),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_415),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_270),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_127),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_139),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_205),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_400),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_164),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_376),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_456),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_576),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_101),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_564),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_434),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_425),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_484),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_426),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_577),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_475),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_242),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_310),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_286),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_68),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_199),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_575),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_472),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_73),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_28),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_607),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_462),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_547),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_43),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_109),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_74),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_59),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_37),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_66),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_144),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_371),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_477),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_61),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_248),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_433),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_46),
.Y(n_757)
);

CKINVDCx16_ASAP7_75t_R g758 ( 
.A(n_226),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_435),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_380),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_594),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_5),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_38),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_362),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_296),
.Y(n_765)
);

INVxp33_ASAP7_75t_SL g766 ( 
.A(n_86),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_191),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_432),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_388),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_437),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_430),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_591),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_422),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_428),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_90),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_119),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_316),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_438),
.Y(n_778)
);

BUFx10_ASAP7_75t_L g779 ( 
.A(n_412),
.Y(n_779)
);

BUFx8_ASAP7_75t_SL g780 ( 
.A(n_65),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_342),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_43),
.Y(n_782)
);

BUFx10_ASAP7_75t_L g783 ( 
.A(n_150),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_124),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_570),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_483),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_420),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_31),
.Y(n_788)
);

CKINVDCx14_ASAP7_75t_R g789 ( 
.A(n_458),
.Y(n_789)
);

BUFx3_ASAP7_75t_L g790 ( 
.A(n_137),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_479),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_106),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_305),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_541),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_446),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_4),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_34),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_419),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_305),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_229),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_551),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_427),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_634),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_257),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_343),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_491),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_628),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_394),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_281),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_497),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_29),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_383),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_405),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_215),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_523),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_282),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_499),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_231),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_556),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_307),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_218),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_540),
.Y(n_822)
);

CKINVDCx20_ASAP7_75t_R g823 ( 
.A(n_299),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_245),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_23),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_129),
.Y(n_826)
);

BUFx2_ASAP7_75t_SL g827 ( 
.A(n_539),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_606),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_402),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_553),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_336),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_372),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_402),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_101),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_300),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_292),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_486),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_98),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_430),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_580),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_133),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_381),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_416),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_133),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_201),
.Y(n_845)
);

INVx1_ASAP7_75t_SL g846 ( 
.A(n_40),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_189),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_424),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_198),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_210),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_334),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_408),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_287),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_362),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_277),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_423),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_426),
.Y(n_857)
);

CKINVDCx20_ASAP7_75t_R g858 ( 
.A(n_121),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_116),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_241),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_154),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_476),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_465),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_117),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_340),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_601),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_622),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_407),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_282),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_592),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_455),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_521),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_245),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_560),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_4),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_110),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_626),
.Y(n_877)
);

CKINVDCx5p33_ASAP7_75t_R g878 ( 
.A(n_200),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_200),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_418),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_636),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_574),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_236),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_139),
.Y(n_884)
);

BUFx10_ASAP7_75t_L g885 ( 
.A(n_151),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_234),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_698),
.Y(n_887)
);

CKINVDCx16_ASAP7_75t_R g888 ( 
.A(n_681),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_718),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_674),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_674),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_674),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_780),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_753),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_780),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_674),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_805),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_674),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_674),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_661),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_694),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_674),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_758),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_675),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_675),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_722),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_722),
.Y(n_907)
);

CKINVDCx20_ASAP7_75t_R g908 ( 
.A(n_641),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_662),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_740),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_740),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_741),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_741),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_774),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_774),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_790),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_790),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_639),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_690),
.Y(n_919)
);

HB1xp67_ASAP7_75t_L g920 ( 
.A(n_873),
.Y(n_920)
);

INVx1_ASAP7_75t_SL g921 ( 
.A(n_875),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_694),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_663),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_639),
.Y(n_924)
);

INVxp67_ASAP7_75t_L g925 ( 
.A(n_876),
.Y(n_925)
);

INVxp33_ASAP7_75t_L g926 ( 
.A(n_730),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_664),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_665),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_639),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_639),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_652),
.Y(n_931)
);

INVxp67_ASAP7_75t_SL g932 ( 
.A(n_652),
.Y(n_932)
);

CKINVDCx20_ASAP7_75t_R g933 ( 
.A(n_641),
.Y(n_933)
);

BUFx2_ASAP7_75t_L g934 ( 
.A(n_638),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_668),
.Y(n_935)
);

CKINVDCx20_ASAP7_75t_R g936 ( 
.A(n_690),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_671),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_652),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_652),
.Y(n_939)
);

CKINVDCx20_ASAP7_75t_R g940 ( 
.A(n_696),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_660),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_679),
.Y(n_942)
);

BUFx6f_ASAP7_75t_SL g943 ( 
.A(n_660),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_679),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_673),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_679),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_679),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_778),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_778),
.Y(n_949)
);

CKINVDCx16_ASAP7_75t_R g950 ( 
.A(n_789),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_778),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_682),
.Y(n_952)
);

BUFx5_ASAP7_75t_L g953 ( 
.A(n_653),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_778),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_648),
.Y(n_955)
);

CKINVDCx20_ASAP7_75t_R g956 ( 
.A(n_648),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_861),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_693),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_861),
.Y(n_959)
);

INVxp67_ASAP7_75t_SL g960 ( 
.A(n_861),
.Y(n_960)
);

INVx2_ASAP7_75t_L g961 ( 
.A(n_861),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_660),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_702),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_637),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_642),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_649),
.Y(n_966)
);

NOR2xp67_ASAP7_75t_L g967 ( 
.A(n_709),
.B(n_0),
.Y(n_967)
);

INVxp67_ASAP7_75t_SL g968 ( 
.A(n_730),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_744),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_654),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_694),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_705),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_667),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_672),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_683),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_684),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_713),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_809),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_687),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_809),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_714),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_723),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_688),
.Y(n_983)
);

INVxp33_ASAP7_75t_SL g984 ( 
.A(n_640),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_724),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_691),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_697),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_701),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_812),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_710),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_932),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_900),
.Y(n_992)
);

INVxp67_ASAP7_75t_SL g993 ( 
.A(n_932),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_908),
.Y(n_994)
);

CKINVDCx20_ASAP7_75t_R g995 ( 
.A(n_933),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_960),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_909),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_960),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_951),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_888),
.Y(n_1000)
);

CKINVDCx16_ASAP7_75t_R g1001 ( 
.A(n_903),
.Y(n_1001)
);

CKINVDCx20_ASAP7_75t_R g1002 ( 
.A(n_955),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_924),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_929),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_894),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_930),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_923),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_951),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_931),
.Y(n_1010)
);

INVxp67_ASAP7_75t_L g1011 ( 
.A(n_934),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_938),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_939),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_927),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_956),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_928),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_935),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_937),
.Y(n_1018)
);

INVxp67_ASAP7_75t_SL g1019 ( 
.A(n_894),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_984),
.B(n_977),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_969),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_945),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_919),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_919),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_952),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_958),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_942),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_944),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_936),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_963),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_972),
.B(n_753),
.Y(n_1031)
);

INVxp33_ASAP7_75t_SL g1032 ( 
.A(n_893),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_981),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_901),
.Y(n_1034)
);

INVxp67_ASAP7_75t_SL g1035 ( 
.A(n_901),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_946),
.Y(n_1036)
);

INVxp67_ASAP7_75t_L g1037 ( 
.A(n_962),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_947),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_961),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_948),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_949),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_954),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_957),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_982),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_985),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_936),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_940),
.Y(n_1047)
);

CKINVDCx20_ASAP7_75t_R g1048 ( 
.A(n_940),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_959),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_895),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_943),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_943),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_897),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_961),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_968),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_920),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_950),
.B(n_807),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1006),
.B(n_810),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_1001),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_991),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_999),
.Y(n_1061)
);

BUFx3_ASAP7_75t_L g1062 ( 
.A(n_996),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_999),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1053),
.B(n_921),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_998),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_993),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1003),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1009),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_1009),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_1039),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1004),
.Y(n_1071)
);

NAND2xp33_ASAP7_75t_R g1072 ( 
.A(n_1045),
.B(n_766),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_1055),
.B(n_666),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_1039),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1019),
.B(n_926),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1034),
.B(n_953),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_1031),
.A2(n_891),
.B(n_890),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_SL g1078 ( 
.A(n_1045),
.B(n_744),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1054),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_1005),
.A2(n_896),
.B(n_892),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1035),
.B(n_953),
.Y(n_1081)
);

BUFx8_ASAP7_75t_L g1082 ( 
.A(n_1007),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1010),
.B(n_953),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1012),
.Y(n_1084)
);

NAND2xp33_ASAP7_75t_R g1085 ( 
.A(n_1050),
.B(n_904),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1013),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1057),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_1056),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1027),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1028),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_1036),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1038),
.B(n_953),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_1023),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1011),
.B(n_926),
.Y(n_1094)
);

AND2x6_ASAP7_75t_L g1095 ( 
.A(n_1020),
.B(n_666),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1040),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_1041),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1042),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1043),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_1049),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1037),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_992),
.B(n_887),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_997),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1008),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_1014),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_1016),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_1017),
.B(n_819),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1018),
.Y(n_1108)
);

INVx5_ASAP7_75t_L g1109 ( 
.A(n_1015),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_1022),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1025),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1026),
.B(n_953),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_1030),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1033),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1044),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_R g1116 ( 
.A(n_1050),
.B(n_905),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1000),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1052),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1051),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_994),
.Y(n_1120)
);

AND2x4_ASAP7_75t_L g1121 ( 
.A(n_994),
.B(n_810),
.Y(n_1121)
);

XNOR2xp5_ASAP7_75t_L g1122 ( 
.A(n_995),
.B(n_874),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_1032),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1032),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_995),
.B(n_978),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1002),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_1002),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1021),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1021),
.Y(n_1129)
);

OR2x2_ASAP7_75t_L g1130 ( 
.A(n_1023),
.B(n_941),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1024),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1048),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1048),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1024),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1029),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1029),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1046),
.Y(n_1137)
);

INVx4_ASAP7_75t_L g1138 ( 
.A(n_1046),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1047),
.B(n_953),
.Y(n_1139)
);

CKINVDCx20_ASAP7_75t_R g1140 ( 
.A(n_1047),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_991),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_991),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_991),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1053),
.B(n_925),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_991),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_991),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1060),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1061),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_1075),
.B(n_694),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_1064),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1061),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1125),
.Y(n_1152)
);

BUFx6f_ASAP7_75t_SL g1153 ( 
.A(n_1110),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1068),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_1087),
.B(n_867),
.Y(n_1155)
);

INVxp33_ASAP7_75t_SL g1156 ( 
.A(n_1078),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1076),
.A2(n_899),
.B(n_898),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1063),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1125),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1068),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_1109),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1065),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1141),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1069),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_1094),
.B(n_889),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_SL g1166 ( 
.A(n_1110),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_1080),
.Y(n_1167)
);

AND3x2_ASAP7_75t_L g1168 ( 
.A(n_1088),
.B(n_731),
.C(n_920),
.Y(n_1168)
);

INVx4_ASAP7_75t_L g1169 ( 
.A(n_1070),
.Y(n_1169)
);

NAND2xp33_ASAP7_75t_SL g1170 ( 
.A(n_1139),
.B(n_874),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1069),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1063),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1066),
.B(n_819),
.Y(n_1173)
);

OAI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1062),
.A2(n_696),
.B1(n_775),
.B2(n_754),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_1062),
.B(n_748),
.Y(n_1175)
);

INVx2_ASAP7_75t_SL g1176 ( 
.A(n_1125),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1142),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1079),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1143),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1079),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1070),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1144),
.B(n_906),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1070),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1070),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1145),
.Y(n_1185)
);

INVx3_ASAP7_75t_L g1186 ( 
.A(n_1074),
.Y(n_1186)
);

AO21x2_ASAP7_75t_L g1187 ( 
.A1(n_1077),
.A2(n_685),
.B(n_656),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1091),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1101),
.B(n_889),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1074),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1146),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1074),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1067),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1112),
.B(n_711),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1095),
.B(n_902),
.Y(n_1195)
);

NOR2xp33_ASAP7_75t_L g1196 ( 
.A(n_1107),
.B(n_846),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1107),
.B(n_853),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1071),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1102),
.Y(n_1199)
);

AND2x2_ASAP7_75t_SL g1200 ( 
.A(n_1121),
.B(n_711),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_1101),
.B(n_864),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1074),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1117),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1086),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1084),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1084),
.Y(n_1206)
);

INVx3_ASAP7_75t_L g1207 ( 
.A(n_1077),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1090),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1089),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1089),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1095),
.B(n_789),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1099),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1098),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1098),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1095),
.B(n_739),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1091),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1058),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1117),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1058),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1091),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1058),
.Y(n_1221)
);

CKINVDCx6p67_ASAP7_75t_R g1222 ( 
.A(n_1109),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1073),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1088),
.B(n_907),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1130),
.B(n_910),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1102),
.B(n_822),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1073),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1091),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1096),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1096),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1108),
.B(n_911),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1096),
.B(n_711),
.Y(n_1232)
);

INVxp33_ASAP7_75t_L g1233 ( 
.A(n_1122),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1096),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1097),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1121),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1097),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1097),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1097),
.Y(n_1239)
);

OR2x6_ASAP7_75t_L g1240 ( 
.A(n_1110),
.B(n_1113),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1100),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1100),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1108),
.B(n_912),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1100),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1083),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1072),
.A2(n_775),
.B1(n_820),
.B2(n_754),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1092),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1081),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1095),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1095),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1121),
.Y(n_1252)
);

INVx8_ASAP7_75t_L g1253 ( 
.A(n_1109),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1105),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1132),
.B(n_913),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1105),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1103),
.Y(n_1257)
);

NOR2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1059),
.B(n_914),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1104),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1114),
.Y(n_1260)
);

BUFx16f_ASAP7_75t_R g1261 ( 
.A(n_1082),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1115),
.Y(n_1262)
);

INVx2_ASAP7_75t_SL g1263 ( 
.A(n_1109),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1118),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1118),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1110),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1085),
.A2(n_726),
.B1(n_732),
.B2(n_729),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1113),
.B(n_711),
.Y(n_1268)
);

AND2x2_ASAP7_75t_SL g1269 ( 
.A(n_1113),
.B(n_882),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1113),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1123),
.B(n_785),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1119),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1124),
.Y(n_1273)
);

NAND2xp33_ASAP7_75t_SL g1274 ( 
.A(n_1085),
.B(n_820),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1106),
.B(n_817),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1124),
.B(n_882),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1124),
.Y(n_1277)
);

INVx6_ASAP7_75t_L g1278 ( 
.A(n_1082),
.Y(n_1278)
);

INVx4_ASAP7_75t_L g1279 ( 
.A(n_1124),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1120),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1106),
.B(n_863),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1111),
.B(n_882),
.Y(n_1282)
);

NAND2xp33_ASAP7_75t_SL g1283 ( 
.A(n_1116),
.B(n_823),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1082),
.Y(n_1284)
);

INVxp67_ASAP7_75t_L g1285 ( 
.A(n_1189),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1178),
.Y(n_1286)
);

BUFx4_ASAP7_75t_L g1287 ( 
.A(n_1261),
.Y(n_1287)
);

AO22x2_ASAP7_75t_L g1288 ( 
.A1(n_1247),
.A2(n_1132),
.B1(n_1134),
.B2(n_1133),
.Y(n_1288)
);

INVx8_ASAP7_75t_L g1289 ( 
.A(n_1253),
.Y(n_1289)
);

AO22x2_ASAP7_75t_L g1290 ( 
.A1(n_1247),
.A2(n_1135),
.B1(n_1137),
.B2(n_1136),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1178),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1180),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1226),
.B(n_1111),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1148),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1150),
.B(n_1257),
.Y(n_1295)
);

INVx3_ASAP7_75t_L g1296 ( 
.A(n_1279),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1180),
.Y(n_1297)
);

AND2x2_ASAP7_75t_SL g1298 ( 
.A(n_1269),
.B(n_1200),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1205),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1153),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1148),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1205),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1151),
.Y(n_1303)
);

OAI21xp33_ASAP7_75t_L g1304 ( 
.A1(n_1226),
.A2(n_644),
.B(n_643),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_1240),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1270),
.B(n_1127),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1279),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_SL g1308 ( 
.A(n_1153),
.B(n_1059),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1206),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1156),
.B(n_1120),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1257),
.B(n_1138),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1249),
.B(n_738),
.Y(n_1312)
);

NAND2xp33_ASAP7_75t_L g1313 ( 
.A(n_1188),
.B(n_742),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1206),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1209),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1209),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1210),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1156),
.B(n_1126),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1225),
.B(n_1128),
.Y(n_1319)
);

AND2x6_ASAP7_75t_L g1320 ( 
.A(n_1250),
.B(n_1251),
.Y(n_1320)
);

AND2x6_ASAP7_75t_L g1321 ( 
.A(n_1248),
.B(n_1127),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1275),
.B(n_1138),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1259),
.B(n_1138),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1210),
.Y(n_1324)
);

INVx3_ASAP7_75t_L g1325 ( 
.A(n_1279),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_SL g1326 ( 
.A(n_1259),
.B(n_1131),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1201),
.B(n_1131),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1151),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1154),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1270),
.B(n_964),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1201),
.B(n_1129),
.Y(n_1331)
);

INVxp67_ASAP7_75t_L g1332 ( 
.A(n_1165),
.Y(n_1332)
);

NOR2xp33_ASAP7_75t_L g1333 ( 
.A(n_1281),
.B(n_1129),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1170),
.A2(n_1116),
.B1(n_1072),
.B2(n_743),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1213),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1240),
.B(n_965),
.Y(n_1336)
);

BUFx6f_ASAP7_75t_L g1337 ( 
.A(n_1240),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1213),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1278),
.B(n_1253),
.Y(n_1339)
);

AND2x4_ASAP7_75t_L g1340 ( 
.A(n_1266),
.B(n_1252),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1260),
.B(n_761),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1222),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1214),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1155),
.B(n_1093),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1252),
.B(n_1273),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1170),
.A2(n_772),
.B1(n_791),
.B2(n_786),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1253),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1154),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1161),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_1260),
.B(n_794),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1160),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1255),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1160),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1164),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1155),
.B(n_1093),
.Y(n_1356)
);

AND2x2_ASAP7_75t_SL g1357 ( 
.A(n_1269),
.B(n_1140),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1164),
.Y(n_1358)
);

INVx4_ASAP7_75t_L g1359 ( 
.A(n_1188),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1166),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1175),
.B(n_915),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1147),
.B(n_795),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1171),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1161),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1162),
.B(n_1163),
.Y(n_1365)
);

AND2x4_ASAP7_75t_L g1366 ( 
.A(n_1252),
.B(n_966),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1188),
.Y(n_1367)
);

AND2x6_ASAP7_75t_L g1368 ( 
.A(n_1254),
.B(n_882),
.Y(n_1368)
);

BUFx4f_ASAP7_75t_L g1369 ( 
.A(n_1222),
.Y(n_1369)
);

INVx4_ASAP7_75t_SL g1370 ( 
.A(n_1166),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1171),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1277),
.B(n_1152),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_L g1373 ( 
.A(n_1199),
.B(n_1140),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1159),
.B(n_970),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1177),
.Y(n_1375)
);

AND2x2_ASAP7_75t_L g1376 ( 
.A(n_1175),
.B(n_1203),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1158),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1188),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1176),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1217),
.A2(n_801),
.B1(n_806),
.B2(n_803),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1172),
.Y(n_1381)
);

AND2x4_ASAP7_75t_L g1382 ( 
.A(n_1236),
.B(n_1219),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1274),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1179),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1182),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1185),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1200),
.B(n_815),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1191),
.B(n_828),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1224),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1193),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_SL g1391 ( 
.A(n_1262),
.Y(n_1391)
);

OR2x6_ASAP7_75t_L g1392 ( 
.A(n_1278),
.B(n_916),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1218),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1198),
.Y(n_1394)
);

BUFx6f_ASAP7_75t_L g1395 ( 
.A(n_1216),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1204),
.Y(n_1396)
);

BUFx3_ASAP7_75t_L g1397 ( 
.A(n_1280),
.Y(n_1397)
);

INVx5_ASAP7_75t_L g1398 ( 
.A(n_1278),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1208),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1231),
.B(n_830),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1172),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1243),
.B(n_1221),
.Y(n_1402)
);

BUFx6f_ASAP7_75t_L g1403 ( 
.A(n_1216),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1220),
.Y(n_1404)
);

AND2x6_ASAP7_75t_L g1405 ( 
.A(n_1256),
.B(n_812),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1158),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1196),
.B(n_917),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1196),
.B(n_968),
.Y(n_1408)
);

INVx4_ASAP7_75t_L g1409 ( 
.A(n_1241),
.Y(n_1409)
);

OAI21xp33_ASAP7_75t_L g1410 ( 
.A1(n_1197),
.A2(n_646),
.B(n_645),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1212),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1220),
.Y(n_1412)
);

INVx3_ASAP7_75t_L g1413 ( 
.A(n_1228),
.Y(n_1413)
);

INVx4_ASAP7_75t_L g1414 ( 
.A(n_1241),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1272),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1181),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1272),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1181),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1228),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

INVx3_ASAP7_75t_L g1421 ( 
.A(n_1229),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_SL g1422 ( 
.A(n_1265),
.B(n_837),
.Y(n_1422)
);

INVx3_ASAP7_75t_L g1423 ( 
.A(n_1229),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1274),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1283),
.Y(n_1425)
);

INVx6_ASAP7_75t_L g1426 ( 
.A(n_1258),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1230),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1263),
.B(n_973),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1230),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1183),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1234),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1199),
.B(n_651),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1199),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1246),
.B(n_840),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1246),
.B(n_862),
.Y(n_1435)
);

AND2x6_ASAP7_75t_L g1436 ( 
.A(n_1207),
.B(n_816),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1234),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1235),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1235),
.Y(n_1439)
);

NAND3xp33_ASAP7_75t_L g1440 ( 
.A(n_1197),
.B(n_967),
.C(n_650),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1283),
.B(n_858),
.Y(n_1441)
);

NOR2xp33_ASAP7_75t_L g1442 ( 
.A(n_1267),
.B(n_823),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1149),
.B(n_866),
.Y(n_1443)
);

AO22x2_ASAP7_75t_L g1444 ( 
.A1(n_1282),
.A2(n_716),
.B1(n_737),
.B2(n_715),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1271),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1237),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1241),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1149),
.B(n_870),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1237),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1282),
.B(n_779),
.Y(n_1450)
);

INVx3_ASAP7_75t_L g1451 ( 
.A(n_1238),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1245),
.A2(n_871),
.B1(n_877),
.B2(n_872),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1173),
.B(n_881),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1284),
.Y(n_1454)
);

OR2x2_ASAP7_75t_L g1455 ( 
.A(n_1233),
.B(n_974),
.Y(n_1455)
);

INVx4_ASAP7_75t_L g1456 ( 
.A(n_1244),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1238),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1239),
.B(n_827),
.Y(n_1458)
);

AND2x6_ASAP7_75t_L g1459 ( 
.A(n_1207),
.B(n_816),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1239),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1242),
.B(n_1244),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1183),
.Y(n_1462)
);

INVxp33_ASAP7_75t_L g1463 ( 
.A(n_1233),
.Y(n_1463)
);

INVx4_ASAP7_75t_L g1464 ( 
.A(n_1186),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1242),
.Y(n_1465)
);

BUFx10_ASAP7_75t_L g1466 ( 
.A(n_1168),
.Y(n_1466)
);

INVx4_ASAP7_75t_SL g1467 ( 
.A(n_1284),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1184),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1184),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1190),
.Y(n_1470)
);

INVxp67_ASAP7_75t_SL g1471 ( 
.A(n_1186),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1190),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1192),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1192),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1202),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1202),
.B(n_975),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1174),
.B(n_829),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1186),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1169),
.B(n_647),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1276),
.B(n_779),
.Y(n_1480)
);

INVx4_ASAP7_75t_L g1481 ( 
.A(n_1169),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1157),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_SL g1483 ( 
.A(n_1169),
.B(n_829),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1232),
.Y(n_1484)
);

INVx4_ASAP7_75t_L g1485 ( 
.A(n_1167),
.Y(n_1485)
);

AND2x6_ASAP7_75t_L g1486 ( 
.A(n_1207),
.B(n_855),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1294),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1408),
.B(n_1276),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1331),
.B(n_1268),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1293),
.B(n_1174),
.Y(n_1490)
);

NOR3xp33_ASAP7_75t_L g1491 ( 
.A(n_1442),
.B(n_1432),
.C(n_1483),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1445),
.B(n_1268),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1415),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1376),
.B(n_1361),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1407),
.B(n_1195),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1389),
.Y(n_1496)
);

INVx6_ASAP7_75t_L g1497 ( 
.A(n_1370),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1306),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1402),
.B(n_1215),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1298),
.B(n_1211),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1301),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1334),
.A2(n_865),
.B1(n_1194),
.B2(n_855),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1303),
.Y(n_1503)
);

INVx3_ASAP7_75t_L g1504 ( 
.A(n_1481),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1417),
.B(n_1194),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1322),
.B(n_1232),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1286),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_L g1508 ( 
.A(n_1289),
.B(n_1167),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1355),
.B(n_1187),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1327),
.B(n_1187),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1291),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1292),
.Y(n_1512)
);

AO221x1_ASAP7_75t_L g1513 ( 
.A1(n_1444),
.A2(n_1290),
.B1(n_1288),
.B2(n_1424),
.C(n_1383),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1433),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1297),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1365),
.B(n_1167),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1310),
.B(n_865),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1328),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1383),
.A2(n_657),
.B1(n_658),
.B2(n_655),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_1357),
.B(n_976),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1400),
.B(n_659),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1375),
.B(n_669),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1384),
.B(n_670),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1299),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1329),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1302),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1351),
.Y(n_1527)
);

NAND2xp33_ASAP7_75t_L g1528 ( 
.A(n_1289),
.B(n_676),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1309),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1353),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1386),
.B(n_677),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1390),
.B(n_678),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1354),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1314),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1352),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1394),
.B(n_680),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_L g1537 ( 
.A(n_1333),
.B(n_686),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1424),
.A2(n_733),
.B1(n_736),
.B2(n_721),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1396),
.B(n_689),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1399),
.B(n_692),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1425),
.A2(n_750),
.B1(n_752),
.B2(n_747),
.Y(n_1541)
);

OAI221xp5_ASAP7_75t_L g1542 ( 
.A1(n_1441),
.A2(n_700),
.B1(n_703),
.B2(n_699),
.C(n_695),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1481),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1411),
.B(n_704),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1312),
.B(n_706),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1425),
.A2(n_708),
.B1(n_712),
.B2(n_707),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1306),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1385),
.B(n_779),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1330),
.B(n_717),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1344),
.B(n_719),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1315),
.Y(n_1551)
);

INVxp33_ASAP7_75t_L g1552 ( 
.A(n_1455),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1330),
.B(n_1366),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1285),
.B(n_783),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1316),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1366),
.B(n_720),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1317),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1434),
.B(n_725),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1324),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1335),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1435),
.B(n_727),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1356),
.B(n_728),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1371),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1338),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1348),
.Y(n_1565)
);

A2O1A1Ixp33_ASAP7_75t_L g1566 ( 
.A1(n_1304),
.A2(n_757),
.B(n_759),
.C(n_755),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1358),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1363),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1381),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1319),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1379),
.B(n_979),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1393),
.Y(n_1572)
);

NOR3xp33_ASAP7_75t_L g1573 ( 
.A(n_1477),
.B(n_986),
.C(n_983),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1409),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_SL g1575 ( 
.A(n_1379),
.B(n_987),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_SL g1576 ( 
.A(n_1347),
.B(n_783),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1401),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1360),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1372),
.B(n_1465),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1372),
.B(n_734),
.Y(n_1580)
);

NOR2xp33_ASAP7_75t_L g1581 ( 
.A(n_1318),
.B(n_735),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1332),
.B(n_1463),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1387),
.A2(n_767),
.B1(n_776),
.B2(n_760),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1465),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1476),
.B(n_745),
.Y(n_1585)
);

NAND2xp33_ASAP7_75t_L g1586 ( 
.A(n_1305),
.B(n_746),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1296),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1476),
.B(n_749),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1420),
.B(n_988),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1379),
.B(n_990),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1397),
.B(n_751),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1307),
.B(n_756),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1305),
.Y(n_1593)
);

AOI22x1_ASAP7_75t_L g1594 ( 
.A1(n_1484),
.A2(n_980),
.B1(n_989),
.B2(n_978),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_SL g1595 ( 
.A(n_1398),
.B(n_784),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1426),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1325),
.B(n_1343),
.Y(n_1597)
);

NOR2xp67_ASAP7_75t_L g1598 ( 
.A(n_1440),
.B(n_439),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1340),
.B(n_762),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1340),
.B(n_763),
.Y(n_1600)
);

NAND3xp33_ASAP7_75t_L g1601 ( 
.A(n_1410),
.B(n_792),
.C(n_788),
.Y(n_1601)
);

NAND2xp33_ASAP7_75t_SL g1602 ( 
.A(n_1305),
.B(n_764),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1472),
.Y(n_1603)
);

AOI221xp5_ASAP7_75t_L g1604 ( 
.A1(n_1288),
.A2(n_1290),
.B1(n_1444),
.B2(n_1450),
.C(n_1391),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1326),
.A2(n_796),
.B(n_798),
.C(n_797),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1337),
.B(n_765),
.Y(n_1606)
);

AOI221xp5_ASAP7_75t_L g1607 ( 
.A1(n_1373),
.A2(n_813),
.B1(n_814),
.B2(n_802),
.C(n_800),
.Y(n_1607)
);

INVxp67_ASAP7_75t_L g1608 ( 
.A(n_1308),
.Y(n_1608)
);

BUFx5_ASAP7_75t_L g1609 ( 
.A(n_1320),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1337),
.B(n_768),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1472),
.B(n_769),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1345),
.B(n_831),
.Y(n_1612)
);

A2O1A1Ixp33_ASAP7_75t_L g1613 ( 
.A1(n_1480),
.A2(n_833),
.B(n_835),
.C(n_832),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1345),
.B(n_841),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1377),
.B(n_843),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1382),
.B(n_770),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1382),
.B(n_771),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1374),
.B(n_773),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1347),
.B(n_783),
.Y(n_1619)
);

BUFx6f_ASAP7_75t_L g1620 ( 
.A(n_1337),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1295),
.B(n_777),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1374),
.B(n_781),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1416),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_SL g1624 ( 
.A(n_1349),
.B(n_782),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1427),
.Y(n_1625)
);

AOI22xp5_ASAP7_75t_L g1626 ( 
.A1(n_1405),
.A2(n_793),
.B1(n_799),
.B2(n_787),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1418),
.Y(n_1627)
);

AO221x1_ASAP7_75t_L g1628 ( 
.A1(n_1395),
.A2(n_879),
.B1(n_880),
.B2(n_850),
.C(n_849),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1428),
.B(n_1336),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1409),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1430),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1429),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1431),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1462),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1349),
.B(n_804),
.Y(n_1635)
);

NAND2x1p5_ASAP7_75t_L g1636 ( 
.A(n_1359),
.B(n_901),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_SL g1637 ( 
.A(n_1349),
.B(n_808),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1311),
.A2(n_886),
.B(n_989),
.C(n_980),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1437),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1405),
.B(n_811),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1362),
.B(n_1388),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1428),
.B(n_818),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1405),
.B(n_821),
.Y(n_1643)
);

NOR2xp67_ASAP7_75t_L g1644 ( 
.A(n_1479),
.B(n_441),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1406),
.B(n_824),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1469),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1364),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1336),
.B(n_825),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1321),
.B(n_1453),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1364),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_SL g1651 ( 
.A(n_1364),
.B(n_826),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1473),
.Y(n_1652)
);

BUFx8_ASAP7_75t_L g1653 ( 
.A(n_1454),
.Y(n_1653)
);

BUFx6f_ASAP7_75t_L g1654 ( 
.A(n_1367),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1370),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1474),
.Y(n_1656)
);

BUFx6f_ASAP7_75t_L g1657 ( 
.A(n_1367),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1438),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1439),
.Y(n_1659)
);

NAND3xp33_ASAP7_75t_L g1660 ( 
.A(n_1346),
.B(n_836),
.C(n_834),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1471),
.A2(n_839),
.B1(n_842),
.B2(n_838),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1359),
.B(n_901),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1321),
.B(n_844),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1446),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1398),
.B(n_845),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1323),
.B(n_847),
.Y(n_1666)
);

BUFx6f_ASAP7_75t_L g1667 ( 
.A(n_1367),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1449),
.Y(n_1668)
);

NOR2xp67_ASAP7_75t_L g1669 ( 
.A(n_1456),
.B(n_443),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1321),
.B(n_848),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1300),
.B(n_851),
.Y(n_1671)
);

BUFx6f_ASAP7_75t_L g1672 ( 
.A(n_1378),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1457),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1475),
.B(n_852),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1378),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1460),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1468),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1470),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1395),
.B(n_1403),
.Y(n_1679)
);

INVxp33_ASAP7_75t_L g1680 ( 
.A(n_1341),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1412),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1395),
.B(n_854),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1426),
.B(n_856),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1350),
.B(n_857),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_SL g1685 ( 
.A(n_1398),
.B(n_859),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1413),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1421),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1422),
.B(n_860),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_SL g1689 ( 
.A(n_1369),
.B(n_885),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1443),
.A2(n_885),
.B1(n_869),
.B2(n_878),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1403),
.B(n_868),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1423),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1403),
.B(n_883),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_SL g1694 ( 
.A(n_1378),
.B(n_884),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1451),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1342),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1494),
.B(n_1448),
.Y(n_1697)
);

AND2x4_ASAP7_75t_L g1698 ( 
.A(n_1629),
.B(n_1339),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1491),
.B(n_1467),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1565),
.Y(n_1700)
);

AND2x6_ASAP7_75t_L g1701 ( 
.A(n_1504),
.B(n_1404),
.Y(n_1701)
);

NAND3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1537),
.B(n_1380),
.C(n_1452),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1507),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1496),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1641),
.B(n_1404),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1490),
.A2(n_1458),
.B(n_1482),
.C(n_1478),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1581),
.B(n_1404),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1511),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1512),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1515),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1567),
.Y(n_1711)
);

AOI22xp5_ASAP7_75t_SL g1712 ( 
.A1(n_1517),
.A2(n_1459),
.B1(n_1486),
.B2(n_1436),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1568),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1489),
.B(n_1392),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1492),
.B(n_1419),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1487),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_SL g1717 ( 
.A(n_1552),
.B(n_1467),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1501),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1550),
.A2(n_1392),
.B1(n_1466),
.B2(n_1313),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1503),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1562),
.B(n_1461),
.C(n_1456),
.Y(n_1721)
);

NAND2x1p5_ASAP7_75t_L g1722 ( 
.A(n_1647),
.B(n_1414),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1584),
.B(n_1419),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1570),
.B(n_1466),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1653),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1524),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1518),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1582),
.B(n_1419),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1525),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1504),
.B(n_1320),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1514),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1653),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1642),
.A2(n_1339),
.B1(n_1459),
.B2(n_1436),
.Y(n_1733)
);

BUFx3_ASAP7_75t_L g1734 ( 
.A(n_1497),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1579),
.B(n_1414),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1495),
.B(n_1447),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1520),
.B(n_1447),
.Y(n_1737)
);

AOI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1591),
.A2(n_1459),
.B1(n_1486),
.B2(n_1436),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1521),
.B(n_1486),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1660),
.A2(n_1502),
.B1(n_1542),
.B2(n_1513),
.Y(n_1740)
);

INVx3_ASAP7_75t_L g1741 ( 
.A(n_1543),
.Y(n_1741)
);

NAND3xp33_ASAP7_75t_SL g1742 ( 
.A(n_1573),
.B(n_1689),
.C(n_1607),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1526),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1493),
.B(n_1464),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1529),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1553),
.B(n_1464),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1534),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1551),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_L g1749 ( 
.A1(n_1506),
.A2(n_1485),
.B1(n_1320),
.B2(n_922),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1527),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1530),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1603),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1533),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1545),
.B(n_1485),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1497),
.Y(n_1755)
);

BUFx3_ASAP7_75t_L g1756 ( 
.A(n_1578),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1558),
.B(n_1368),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1555),
.Y(n_1758)
);

INVx2_ASAP7_75t_SL g1759 ( 
.A(n_1596),
.Y(n_1759)
);

BUFx2_ASAP7_75t_L g1760 ( 
.A(n_1535),
.Y(n_1760)
);

BUFx12f_ASAP7_75t_L g1761 ( 
.A(n_1696),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1561),
.B(n_1368),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1589),
.B(n_885),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1557),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1559),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1655),
.B(n_1287),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1683),
.A2(n_1368),
.B1(n_1287),
.B2(n_971),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1563),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1560),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1593),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1499),
.B(n_1488),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1543),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1564),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1608),
.Y(n_1774)
);

BUFx2_ASAP7_75t_SL g1775 ( 
.A(n_1647),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1612),
.B(n_0),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1660),
.A2(n_971),
.B1(n_922),
.B2(n_3),
.Y(n_1777)
);

BUFx6f_ASAP7_75t_L g1778 ( 
.A(n_1593),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1593),
.Y(n_1779)
);

NOR2x1p5_ASAP7_75t_L g1780 ( 
.A(n_1618),
.B(n_922),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1574),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1625),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1632),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1680),
.B(n_1),
.Y(n_1784)
);

AND2x4_ASAP7_75t_L g1785 ( 
.A(n_1498),
.B(n_444),
.Y(n_1785)
);

BUFx3_ASAP7_75t_L g1786 ( 
.A(n_1620),
.Y(n_1786)
);

INVxp67_ASAP7_75t_SL g1787 ( 
.A(n_1574),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1633),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1589),
.B(n_922),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_L g1790 ( 
.A1(n_1684),
.A2(n_1688),
.B(n_1666),
.C(n_1601),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1612),
.B(n_1),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1614),
.B(n_2),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1614),
.B(n_2),
.Y(n_1793)
);

BUFx6f_ASAP7_75t_L g1794 ( 
.A(n_1620),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1639),
.Y(n_1795)
);

AND2x4_ASAP7_75t_SL g1796 ( 
.A(n_1620),
.B(n_971),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1658),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1572),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1538),
.B(n_3),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1647),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1541),
.B(n_5),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_1654),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1611),
.B(n_1622),
.Y(n_1803)
);

NOR2xp67_ASAP7_75t_L g1804 ( 
.A(n_1682),
.B(n_1691),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1548),
.B(n_6),
.Y(n_1805)
);

INVx5_ASAP7_75t_L g1806 ( 
.A(n_1654),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1673),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1677),
.Y(n_1808)
);

NOR2xp33_ASAP7_75t_L g1809 ( 
.A(n_1621),
.B(n_6),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1615),
.B(n_7),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1689),
.B(n_971),
.Y(n_1811)
);

INVx3_ASAP7_75t_L g1812 ( 
.A(n_1630),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1615),
.B(n_7),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1678),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1693),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1648),
.B(n_8),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1650),
.Y(n_1817)
);

NOR2x2_ASAP7_75t_L g1818 ( 
.A(n_1681),
.B(n_9),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1650),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1671),
.A2(n_11),
.B1(n_9),
.B2(n_10),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1601),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1522),
.B(n_12),
.Y(n_1822)
);

INVx5_ASAP7_75t_L g1823 ( 
.A(n_1654),
.Y(n_1823)
);

INVx8_ASAP7_75t_L g1824 ( 
.A(n_1657),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1659),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1650),
.Y(n_1826)
);

NOR2x1p5_ASAP7_75t_L g1827 ( 
.A(n_1556),
.B(n_445),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1547),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_L g1829 ( 
.A1(n_1516),
.A2(n_448),
.B(n_447),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1657),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1576),
.B(n_13),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1657),
.B(n_449),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1674),
.B(n_13),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1624),
.B(n_450),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1523),
.B(n_1531),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1519),
.B(n_14),
.Y(n_1836)
);

OAI22xp5_ASAP7_75t_SL g1837 ( 
.A1(n_1690),
.A2(n_17),
.B1(n_15),
.B2(n_16),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1664),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1668),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1532),
.B(n_15),
.Y(n_1840)
);

INVx5_ASAP7_75t_L g1841 ( 
.A(n_1667),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1676),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1604),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1843)
);

BUFx2_ASAP7_75t_L g1844 ( 
.A(n_1667),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1549),
.B(n_18),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1602),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1628),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_1847)
);

NOR2xp33_ASAP7_75t_L g1848 ( 
.A(n_1519),
.B(n_19),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1546),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1569),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1577),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1554),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1546),
.B(n_1599),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1536),
.B(n_23),
.Y(n_1854)
);

INVx4_ASAP7_75t_L g1855 ( 
.A(n_1667),
.Y(n_1855)
);

BUFx3_ASAP7_75t_L g1856 ( 
.A(n_1672),
.Y(n_1856)
);

INVx2_ASAP7_75t_SL g1857 ( 
.A(n_1672),
.Y(n_1857)
);

NOR2xp67_ASAP7_75t_L g1858 ( 
.A(n_1663),
.B(n_451),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1623),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1539),
.B(n_24),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_SL g1861 ( 
.A(n_1576),
.B(n_24),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1540),
.B(n_25),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1644),
.A2(n_27),
.B(n_25),
.C(n_26),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1627),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1619),
.B(n_26),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1619),
.B(n_27),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1544),
.B(n_28),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1672),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1631),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1509),
.A2(n_453),
.B(n_452),
.Y(n_1870)
);

AND2x4_ASAP7_75t_L g1871 ( 
.A(n_1635),
.B(n_1637),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1634),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1600),
.B(n_29),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1646),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1652),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1585),
.B(n_30),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1675),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1613),
.B(n_30),
.Y(n_1878)
);

BUFx4f_ASAP7_75t_L g1879 ( 
.A(n_1675),
.Y(n_1879)
);

AND2x6_ASAP7_75t_L g1880 ( 
.A(n_1630),
.B(n_459),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1588),
.B(n_32),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1694),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1675),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1594),
.Y(n_1884)
);

AOI22xp33_ASAP7_75t_L g1885 ( 
.A1(n_1583),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1679),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_SL g1887 ( 
.A(n_1626),
.B(n_1592),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1656),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1686),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1597),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1580),
.B(n_1616),
.Y(n_1891)
);

BUFx4f_ASAP7_75t_L g1892 ( 
.A(n_1687),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1617),
.B(n_35),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1505),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1790),
.A2(n_1508),
.B(n_1500),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1795),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1734),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1731),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1835),
.B(n_1626),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_L g1900 ( 
.A(n_1815),
.B(n_1606),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1807),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1740),
.A2(n_1670),
.B1(n_1587),
.B2(n_1643),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1853),
.B(n_1661),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1771),
.B(n_1661),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1697),
.B(n_1566),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1714),
.B(n_1692),
.Y(n_1906)
);

A2O1A1Ixp33_ASAP7_75t_L g1907 ( 
.A1(n_1809),
.A2(n_1598),
.B(n_1644),
.C(n_1640),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1894),
.B(n_1645),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1703),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1803),
.B(n_1610),
.Y(n_1910)
);

AOI22xp5_ASAP7_75t_L g1911 ( 
.A1(n_1742),
.A2(n_1651),
.B1(n_1586),
.B2(n_1665),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1774),
.B(n_1571),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1700),
.Y(n_1913)
);

NOR3xp33_ASAP7_75t_L g1914 ( 
.A(n_1702),
.B(n_1685),
.C(n_1528),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1894),
.B(n_1575),
.Y(n_1915)
);

BUFx6f_ASAP7_75t_L g1916 ( 
.A(n_1879),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1890),
.B(n_1590),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1891),
.B(n_1695),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_SL g1919 ( 
.A(n_1804),
.B(n_1649),
.Y(n_1919)
);

OAI22xp5_ASAP7_75t_L g1920 ( 
.A1(n_1852),
.A2(n_1719),
.B1(n_1705),
.B2(n_1843),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1887),
.A2(n_1510),
.B(n_1669),
.Y(n_1921)
);

AOI21xp5_ASAP7_75t_L g1922 ( 
.A1(n_1754),
.A2(n_1669),
.B(n_1598),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_1704),
.B(n_1595),
.Y(n_1923)
);

BUFx4f_ASAP7_75t_L g1924 ( 
.A(n_1761),
.Y(n_1924)
);

AOI22xp5_ASAP7_75t_L g1925 ( 
.A1(n_1816),
.A2(n_1609),
.B1(n_1662),
.B2(n_1636),
.Y(n_1925)
);

OR2x6_ASAP7_75t_L g1926 ( 
.A(n_1832),
.B(n_1605),
.Y(n_1926)
);

OAI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1706),
.A2(n_1638),
.B(n_1636),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1890),
.B(n_1609),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1736),
.A2(n_1662),
.B(n_1609),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1707),
.B(n_1609),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1739),
.A2(n_1609),
.B(n_631),
.Y(n_1931)
);

A2O1A1Ixp33_ASAP7_75t_L g1932 ( 
.A1(n_1836),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1932)
);

AOI22x1_ASAP7_75t_L g1933 ( 
.A1(n_1780),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1848),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_1934)
);

AOI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1721),
.A2(n_1749),
.B(n_1757),
.Y(n_1935)
);

OAI22x1_ASAP7_75t_L g1936 ( 
.A1(n_1820),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.Y(n_1936)
);

NOR2xp33_ASAP7_75t_L g1937 ( 
.A(n_1798),
.B(n_454),
.Y(n_1937)
);

AOI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1762),
.A2(n_618),
.B(n_617),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1828),
.B(n_457),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1787),
.A2(n_621),
.B(n_620),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1737),
.B(n_44),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1805),
.B(n_45),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1893),
.B(n_1776),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1756),
.B(n_1698),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1879),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1791),
.B(n_46),
.Y(n_1946)
);

AOI21xp5_ASAP7_75t_L g1947 ( 
.A1(n_1712),
.A2(n_1746),
.B(n_1870),
.Y(n_1947)
);

A2O1A1Ixp33_ASAP7_75t_L g1948 ( 
.A1(n_1833),
.A2(n_1873),
.B(n_1840),
.C(n_1854),
.Y(n_1948)
);

AO21x1_ASAP7_75t_L g1949 ( 
.A1(n_1699),
.A2(n_47),
.B(n_48),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1698),
.B(n_460),
.Y(n_1950)
);

BUFx12f_ASAP7_75t_L g1951 ( 
.A(n_1725),
.Y(n_1951)
);

O2A1O1Ixp33_ASAP7_75t_SL g1952 ( 
.A1(n_1863),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1738),
.A2(n_635),
.B(n_463),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1834),
.B(n_49),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1785),
.B(n_50),
.Y(n_1955)
);

BUFx12f_ASAP7_75t_L g1956 ( 
.A(n_1732),
.Y(n_1956)
);

OAI22xp5_ASAP7_75t_L g1957 ( 
.A1(n_1715),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1766),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1831),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1829),
.A2(n_613),
.B(n_612),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1822),
.A2(n_55),
.B(n_53),
.C(n_54),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1708),
.Y(n_1962)
);

NAND3xp33_ASAP7_75t_L g1963 ( 
.A(n_1821),
.B(n_54),
.C(n_55),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1860),
.B(n_1862),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1793),
.B(n_56),
.Y(n_1965)
);

AOI21xp5_ASAP7_75t_L g1966 ( 
.A1(n_1735),
.A2(n_625),
.B(n_624),
.Y(n_1966)
);

A2O1A1Ixp33_ASAP7_75t_L g1967 ( 
.A1(n_1867),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1711),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1709),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1810),
.B(n_57),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1834),
.B(n_58),
.Y(n_1971)
);

OAI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1881),
.A2(n_1813),
.B(n_1777),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1871),
.B(n_59),
.Y(n_1973)
);

O2A1O1Ixp5_ASAP7_75t_L g1974 ( 
.A1(n_1811),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1974)
);

OAI22xp5_ASAP7_75t_L g1975 ( 
.A1(n_1733),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.Y(n_1975)
);

OAI21xp5_ASAP7_75t_L g1976 ( 
.A1(n_1728),
.A2(n_63),
.B(n_64),
.Y(n_1976)
);

OAI321xp33_ASAP7_75t_L g1977 ( 
.A1(n_1849),
.A2(n_66),
.A3(n_68),
.B1(n_64),
.B2(n_65),
.C(n_67),
.Y(n_1977)
);

INVx5_ASAP7_75t_L g1978 ( 
.A(n_1701),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1752),
.B(n_67),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1871),
.B(n_69),
.Y(n_1980)
);

OAI21xp33_ASAP7_75t_L g1981 ( 
.A1(n_1878),
.A2(n_69),
.B(n_70),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1799),
.A2(n_70),
.B(n_71),
.Y(n_1982)
);

O2A1O1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1861),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1785),
.B(n_72),
.Y(n_1984)
);

AOI21xp5_ASAP7_75t_L g1985 ( 
.A1(n_1741),
.A2(n_464),
.B(n_461),
.Y(n_1985)
);

O2A1O1Ixp33_ASAP7_75t_L g1986 ( 
.A1(n_1865),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_L g1987 ( 
.A(n_1760),
.B(n_466),
.Y(n_1987)
);

NAND2x1p5_ASAP7_75t_L g1988 ( 
.A(n_1806),
.B(n_467),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1806),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1801),
.B(n_75),
.Y(n_1990)
);

O2A1O1Ixp33_ASAP7_75t_L g1991 ( 
.A1(n_1866),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_1991)
);

AOI21xp5_ASAP7_75t_L g1992 ( 
.A1(n_1741),
.A2(n_633),
.B(n_470),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1772),
.A2(n_632),
.B(n_471),
.Y(n_1993)
);

BUFx2_ASAP7_75t_L g1994 ( 
.A(n_1800),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1792),
.B(n_77),
.Y(n_1995)
);

AOI21xp33_ASAP7_75t_L g1996 ( 
.A1(n_1845),
.A2(n_78),
.B(n_79),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1763),
.B(n_468),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1876),
.B(n_473),
.Y(n_1998)
);

O2A1O1Ixp5_ASAP7_75t_L g1999 ( 
.A1(n_1724),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1892),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_2000)
);

OR2x6_ASAP7_75t_L g2001 ( 
.A(n_1832),
.B(n_480),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1846),
.B(n_481),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1886),
.B(n_82),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1723),
.Y(n_2004)
);

NOR2xp67_ASAP7_75t_L g2005 ( 
.A(n_1759),
.B(n_485),
.Y(n_2005)
);

OAI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1858),
.A2(n_83),
.B(n_84),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1781),
.A2(n_488),
.B(n_487),
.Y(n_2007)
);

AOI21xp5_ASAP7_75t_L g2008 ( 
.A1(n_1812),
.A2(n_490),
.B(n_489),
.Y(n_2008)
);

OR2x6_ASAP7_75t_L g2009 ( 
.A(n_1775),
.B(n_492),
.Y(n_2009)
);

OAI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1882),
.A2(n_83),
.B(n_84),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1713),
.B(n_1825),
.Y(n_2011)
);

AOI21xp5_ASAP7_75t_L g2012 ( 
.A1(n_1812),
.A2(n_629),
.B(n_494),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1806),
.B(n_493),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1817),
.B(n_495),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1838),
.B(n_85),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1710),
.Y(n_2016)
);

AOI21xp5_ASAP7_75t_L g2017 ( 
.A1(n_1744),
.A2(n_627),
.B(n_498),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1839),
.B(n_85),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1770),
.B(n_496),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_1823),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1726),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1842),
.B(n_86),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1716),
.Y(n_2023)
);

BUFx3_ASAP7_75t_L g2024 ( 
.A(n_1786),
.Y(n_2024)
);

AOI21xp5_ASAP7_75t_L g2025 ( 
.A1(n_1884),
.A2(n_501),
.B(n_500),
.Y(n_2025)
);

BUFx6f_ASAP7_75t_L g2026 ( 
.A(n_1823),
.Y(n_2026)
);

O2A1O1Ixp33_ASAP7_75t_SL g2027 ( 
.A1(n_1789),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1889),
.B(n_502),
.Y(n_2028)
);

AOI21xp5_ASAP7_75t_L g2029 ( 
.A1(n_1884),
.A2(n_504),
.B(n_503),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_SL g2030 ( 
.A(n_1784),
.B(n_88),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1892),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1722),
.A2(n_619),
.B(n_506),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_SL g2033 ( 
.A(n_1755),
.B(n_505),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1888),
.B(n_91),
.Y(n_2034)
);

OAI21xp5_ASAP7_75t_L g2035 ( 
.A1(n_1767),
.A2(n_92),
.B(n_93),
.Y(n_2035)
);

AOI33xp33_ASAP7_75t_L g2036 ( 
.A1(n_1885),
.A2(n_95),
.A3(n_97),
.B1(n_92),
.B2(n_94),
.B3(n_96),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1718),
.B(n_94),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1720),
.B(n_95),
.Y(n_2038)
);

AOI22xp5_ASAP7_75t_L g2039 ( 
.A1(n_1837),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1727),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1847),
.A2(n_99),
.B(n_100),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1729),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1750),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1751),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1743),
.Y(n_2045)
);

NOR2xp33_ASAP7_75t_L g2046 ( 
.A(n_1717),
.B(n_507),
.Y(n_2046)
);

AOI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1745),
.A2(n_1748),
.B(n_1747),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1753),
.B(n_100),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1768),
.B(n_508),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1851),
.B(n_102),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1864),
.B(n_103),
.Y(n_2051)
);

OAI22xp5_ASAP7_75t_L g2052 ( 
.A1(n_1758),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_2052)
);

OAI21x1_ASAP7_75t_L g2053 ( 
.A1(n_1764),
.A2(n_511),
.B(n_509),
.Y(n_2053)
);

AOI21x1_ASAP7_75t_L g2054 ( 
.A1(n_1765),
.A2(n_513),
.B(n_512),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1850),
.B(n_104),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1859),
.B(n_105),
.Y(n_2056)
);

A2O1A1Ixp33_ASAP7_75t_L g2057 ( 
.A1(n_1827),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1769),
.A2(n_616),
.B(n_515),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1773),
.A2(n_615),
.B(n_516),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1869),
.B(n_514),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_1872),
.B(n_110),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_1874),
.B(n_111),
.Y(n_2062)
);

NAND2x1p5_ASAP7_75t_L g2063 ( 
.A(n_1823),
.B(n_517),
.Y(n_2063)
);

NOR3xp33_ASAP7_75t_L g2064 ( 
.A(n_1875),
.B(n_1783),
.C(n_1782),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1788),
.B(n_111),
.Y(n_2065)
);

AOI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1797),
.A2(n_611),
.B(n_519),
.Y(n_2066)
);

BUFx6f_ASAP7_75t_L g2067 ( 
.A(n_1841),
.Y(n_2067)
);

AOI221x1_ASAP7_75t_L g2068 ( 
.A1(n_1948),
.A2(n_1814),
.B1(n_1808),
.B2(n_1794),
.C(n_1779),
.Y(n_2068)
);

AOI21xp5_ASAP7_75t_L g2069 ( 
.A1(n_1921),
.A2(n_1841),
.B(n_1796),
.Y(n_2069)
);

OAI21x1_ASAP7_75t_L g2070 ( 
.A1(n_1895),
.A2(n_1830),
.B(n_1880),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1901),
.Y(n_2071)
);

AND3x4_ASAP7_75t_L g2072 ( 
.A(n_1944),
.B(n_1818),
.C(n_1856),
.Y(n_2072)
);

OAI21xp5_ASAP7_75t_L g2073 ( 
.A1(n_1907),
.A2(n_1880),
.B(n_1730),
.Y(n_2073)
);

OAI21xp5_ASAP7_75t_L g2074 ( 
.A1(n_1903),
.A2(n_1880),
.B(n_1730),
.Y(n_2074)
);

BUFx2_ASAP7_75t_L g2075 ( 
.A(n_1994),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1909),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1964),
.B(n_1844),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1929),
.A2(n_1880),
.B(n_1730),
.Y(n_2078)
);

OA21x2_ASAP7_75t_L g2079 ( 
.A1(n_1935),
.A2(n_1927),
.B(n_1922),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1943),
.B(n_1819),
.Y(n_2080)
);

AND2x4_ASAP7_75t_L g2081 ( 
.A(n_2004),
.B(n_1841),
.Y(n_2081)
);

OAI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1972),
.A2(n_1730),
.B(n_1701),
.Y(n_2082)
);

AOI21x1_ASAP7_75t_L g2083 ( 
.A1(n_1947),
.A2(n_1766),
.B(n_1826),
.Y(n_2083)
);

INVx3_ASAP7_75t_L g2084 ( 
.A(n_1978),
.Y(n_2084)
);

OAI21xp5_ASAP7_75t_SL g2085 ( 
.A1(n_2039),
.A2(n_1779),
.B(n_1778),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1908),
.B(n_1778),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1962),
.Y(n_2087)
);

OAI21xp5_ASAP7_75t_L g2088 ( 
.A1(n_2010),
.A2(n_1701),
.B(n_1857),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1899),
.A2(n_1824),
.B(n_1701),
.Y(n_2089)
);

INVx8_ASAP7_75t_L g2090 ( 
.A(n_1978),
.Y(n_2090)
);

OAI21x1_ASAP7_75t_L g2091 ( 
.A1(n_2053),
.A2(n_1883),
.B(n_1855),
.Y(n_2091)
);

AOI21x1_ASAP7_75t_L g2092 ( 
.A1(n_1919),
.A2(n_1877),
.B(n_1868),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1904),
.B(n_1778),
.Y(n_2093)
);

AOI21xp5_ASAP7_75t_L g2094 ( 
.A1(n_1905),
.A2(n_1824),
.B(n_1855),
.Y(n_2094)
);

OAI21x1_ASAP7_75t_L g2095 ( 
.A1(n_2054),
.A2(n_1883),
.B(n_1802),
.Y(n_2095)
);

OAI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_1911),
.A2(n_1794),
.B1(n_1779),
.B2(n_1802),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1910),
.B(n_1918),
.Y(n_2097)
);

OAI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1902),
.A2(n_1794),
.B(n_1802),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1920),
.B(n_112),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1960),
.A2(n_520),
.B(n_518),
.Y(n_2100)
);

AOI21xp5_ASAP7_75t_SL g2101 ( 
.A1(n_2001),
.A2(n_524),
.B(n_522),
.Y(n_2101)
);

OAI21x1_ASAP7_75t_L g2102 ( 
.A1(n_1931),
.A2(n_527),
.B(n_525),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_1928),
.A2(n_530),
.B(n_529),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1917),
.B(n_112),
.Y(n_2104)
);

AOI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_1978),
.A2(n_532),
.B(n_531),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_1912),
.B(n_533),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1913),
.Y(n_2107)
);

OAI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_1900),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_2108)
);

BUFx2_ASAP7_75t_L g2109 ( 
.A(n_2024),
.Y(n_2109)
);

OAI21x1_ASAP7_75t_L g2110 ( 
.A1(n_2047),
.A2(n_535),
.B(n_534),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_1968),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1953),
.A2(n_537),
.B(n_536),
.Y(n_2112)
);

AOI21xp5_ASAP7_75t_L g2113 ( 
.A1(n_1914),
.A2(n_542),
.B(n_538),
.Y(n_2113)
);

INVx4_ASAP7_75t_L g2114 ( 
.A(n_1989),
.Y(n_2114)
);

O2A1O1Ixp5_ASAP7_75t_L g2115 ( 
.A1(n_1982),
.A2(n_116),
.B(n_114),
.C(n_115),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_SL g2116 ( 
.A(n_2001),
.B(n_117),
.Y(n_2116)
);

AOI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_1930),
.A2(n_544),
.B(n_543),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_1938),
.A2(n_546),
.B(n_545),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_1906),
.Y(n_2119)
);

AND2x4_ASAP7_75t_L g2120 ( 
.A(n_2064),
.B(n_548),
.Y(n_2120)
);

AOI21xp5_ASAP7_75t_L g2121 ( 
.A1(n_1966),
.A2(n_554),
.B(n_549),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_SL g2122 ( 
.A(n_2035),
.B(n_118),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1916),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_L g2124 ( 
.A1(n_1934),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1915),
.B(n_121),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1973),
.B(n_122),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1969),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2023),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1980),
.B(n_122),
.Y(n_2129)
);

AOI221xp5_ASAP7_75t_L g2130 ( 
.A1(n_1977),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_2130)
);

AOI21xp33_ASAP7_75t_L g2131 ( 
.A1(n_1963),
.A2(n_123),
.B(n_125),
.Y(n_2131)
);

OAI21x1_ASAP7_75t_L g2132 ( 
.A1(n_2025),
.A2(n_557),
.B(n_555),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2016),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2036),
.B(n_126),
.Y(n_2134)
);

NOR2xp67_ASAP7_75t_L g2135 ( 
.A(n_1896),
.B(n_558),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_2029),
.A2(n_1992),
.B(n_1985),
.Y(n_2136)
);

A2O1A1Ixp33_ASAP7_75t_L g2137 ( 
.A1(n_2041),
.A2(n_1997),
.B(n_2006),
.C(n_1981),
.Y(n_2137)
);

OAI22x1_ASAP7_75t_L g2138 ( 
.A1(n_1933),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2048),
.B(n_559),
.Y(n_2139)
);

OAI21xp5_ASAP7_75t_L g2140 ( 
.A1(n_1932),
.A2(n_128),
.B(n_130),
.Y(n_2140)
);

INVx3_ASAP7_75t_L g2141 ( 
.A(n_1989),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1942),
.B(n_1955),
.Y(n_2142)
);

AOI21x1_ASAP7_75t_SL g2143 ( 
.A1(n_1970),
.A2(n_130),
.B(n_131),
.Y(n_2143)
);

AOI21xp5_ASAP7_75t_SL g2144 ( 
.A1(n_2009),
.A2(n_566),
.B(n_561),
.Y(n_2144)
);

OAI21x1_ASAP7_75t_L g2145 ( 
.A1(n_1993),
.A2(n_568),
.B(n_567),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1940),
.A2(n_571),
.B(n_569),
.Y(n_2146)
);

BUFx3_ASAP7_75t_L g2147 ( 
.A(n_1897),
.Y(n_2147)
);

OAI21x1_ASAP7_75t_SL g2148 ( 
.A1(n_1949),
.A2(n_131),
.B(n_132),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_SL g2149 ( 
.A(n_1923),
.B(n_573),
.Y(n_2149)
);

OAI21xp5_ASAP7_75t_L g2150 ( 
.A1(n_2057),
.A2(n_132),
.B(n_134),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_1996),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.C(n_137),
.Y(n_2151)
);

AOI21x1_ASAP7_75t_L g2152 ( 
.A1(n_1941),
.A2(n_579),
.B(n_578),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2011),
.B(n_135),
.Y(n_2153)
);

OAI21x1_ASAP7_75t_L g2154 ( 
.A1(n_2007),
.A2(n_582),
.B(n_581),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_SL g2155 ( 
.A(n_1998),
.B(n_583),
.Y(n_2155)
);

BUFx3_ASAP7_75t_L g2156 ( 
.A(n_1951),
.Y(n_2156)
);

AOI21xp5_ASAP7_75t_L g2157 ( 
.A1(n_2058),
.A2(n_585),
.B(n_584),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2040),
.B(n_136),
.Y(n_2158)
);

AOI21xp5_ASAP7_75t_L g2159 ( 
.A1(n_2059),
.A2(n_587),
.B(n_586),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2042),
.B(n_138),
.Y(n_2160)
);

AOI21xp5_ASAP7_75t_L g2161 ( 
.A1(n_2066),
.A2(n_590),
.B(n_589),
.Y(n_2161)
);

AOI21xp5_ASAP7_75t_L g2162 ( 
.A1(n_1952),
.A2(n_595),
.B(n_593),
.Y(n_2162)
);

AND2x4_ASAP7_75t_L g2163 ( 
.A(n_1950),
.B(n_596),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1925),
.B(n_597),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_2021),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2043),
.B(n_138),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_2044),
.B(n_1990),
.Y(n_2167)
);

OAI21x1_ASAP7_75t_SL g2168 ( 
.A1(n_1976),
.A2(n_140),
.B(n_141),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_1926),
.A2(n_599),
.B(n_598),
.Y(n_2169)
);

A2O1A1Ixp33_ASAP7_75t_L g2170 ( 
.A1(n_1946),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_2170)
);

AO21x2_ASAP7_75t_L g2171 ( 
.A1(n_2045),
.A2(n_142),
.B(n_143),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_2008),
.A2(n_604),
.B(n_600),
.Y(n_2172)
);

INVx2_ASAP7_75t_SL g2173 ( 
.A(n_1898),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2015),
.Y(n_2174)
);

NAND2x1_ASAP7_75t_L g2175 ( 
.A(n_1926),
.B(n_2009),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2018),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2034),
.Y(n_2177)
);

INVx1_ASAP7_75t_SL g2178 ( 
.A(n_2003),
.Y(n_2178)
);

OAI21xp5_ASAP7_75t_L g2179 ( 
.A1(n_1961),
.A2(n_143),
.B(n_144),
.Y(n_2179)
);

OAI21xp5_ASAP7_75t_L g2180 ( 
.A1(n_1967),
.A2(n_145),
.B(n_146),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2022),
.Y(n_2181)
);

OAI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_1999),
.A2(n_145),
.B(n_146),
.Y(n_2182)
);

AO31x2_ASAP7_75t_L g2183 ( 
.A1(n_1975),
.A2(n_608),
.A3(n_609),
.B(n_605),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_1954),
.B(n_147),
.Y(n_2184)
);

BUFx2_ASAP7_75t_R g2185 ( 
.A(n_2156),
.Y(n_2185)
);

INVx2_ASAP7_75t_L g2186 ( 
.A(n_2076),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2087),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2127),
.Y(n_2188)
);

BUFx6f_ASAP7_75t_L g2189 ( 
.A(n_2123),
.Y(n_2189)
);

INVx2_ASAP7_75t_SL g2190 ( 
.A(n_2147),
.Y(n_2190)
);

BUFx3_ASAP7_75t_L g2191 ( 
.A(n_2109),
.Y(n_2191)
);

INVx5_ASAP7_75t_L g2192 ( 
.A(n_2090),
.Y(n_2192)
);

AOI22xp33_ASAP7_75t_L g2193 ( 
.A1(n_2122),
.A2(n_1936),
.B1(n_2030),
.B2(n_1971),
.Y(n_2193)
);

INVx5_ASAP7_75t_L g2194 ( 
.A(n_2090),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_2081),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_2133),
.Y(n_2196)
);

INVx1_ASAP7_75t_SL g2197 ( 
.A(n_2119),
.Y(n_2197)
);

BUFx12f_ASAP7_75t_L g2198 ( 
.A(n_2123),
.Y(n_2198)
);

NOR2x1_ASAP7_75t_SL g2199 ( 
.A(n_2083),
.B(n_1989),
.Y(n_2199)
);

AND2x2_ASAP7_75t_L g2200 ( 
.A(n_2142),
.B(n_1979),
.Y(n_2200)
);

BUFx4f_ASAP7_75t_L g2201 ( 
.A(n_2123),
.Y(n_2201)
);

BUFx12f_ASAP7_75t_L g2202 ( 
.A(n_2173),
.Y(n_2202)
);

BUFx3_ASAP7_75t_L g2203 ( 
.A(n_2075),
.Y(n_2203)
);

BUFx2_ASAP7_75t_SL g2204 ( 
.A(n_2081),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2165),
.Y(n_2205)
);

BUFx6f_ASAP7_75t_L g2206 ( 
.A(n_2090),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2097),
.B(n_1965),
.Y(n_2207)
);

INVxp67_ASAP7_75t_SL g2208 ( 
.A(n_2079),
.Y(n_2208)
);

INVx4_ASAP7_75t_L g2209 ( 
.A(n_2084),
.Y(n_2209)
);

OAI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_2137),
.A2(n_1958),
.B1(n_1984),
.B2(n_2000),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2178),
.B(n_1995),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_2178),
.B(n_2065),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2071),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2107),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_2141),
.Y(n_2215)
);

BUFx12f_ASAP7_75t_L g2216 ( 
.A(n_2114),
.Y(n_2216)
);

INVx2_ASAP7_75t_L g2217 ( 
.A(n_2111),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2077),
.Y(n_2218)
);

BUFx6f_ASAP7_75t_L g2219 ( 
.A(n_2175),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_2141),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_2114),
.Y(n_2221)
);

BUFx6f_ASAP7_75t_L g2222 ( 
.A(n_2084),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2174),
.B(n_2055),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2080),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2128),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2171),
.Y(n_2226)
);

BUFx12f_ASAP7_75t_L g2227 ( 
.A(n_2163),
.Y(n_2227)
);

BUFx6f_ASAP7_75t_L g2228 ( 
.A(n_2086),
.Y(n_2228)
);

BUFx2_ASAP7_75t_L g2229 ( 
.A(n_2093),
.Y(n_2229)
);

BUFx12f_ASAP7_75t_L g2230 ( 
.A(n_2163),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_2092),
.Y(n_2231)
);

INVx1_ASAP7_75t_SL g2232 ( 
.A(n_2167),
.Y(n_2232)
);

CKINVDCx20_ASAP7_75t_R g2233 ( 
.A(n_2106),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2171),
.Y(n_2234)
);

BUFx2_ASAP7_75t_L g2235 ( 
.A(n_2098),
.Y(n_2235)
);

INVx5_ASAP7_75t_L g2236 ( 
.A(n_2120),
.Y(n_2236)
);

BUFx6f_ASAP7_75t_L g2237 ( 
.A(n_2070),
.Y(n_2237)
);

INVxp67_ASAP7_75t_SL g2238 ( 
.A(n_2079),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2176),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_2091),
.Y(n_2240)
);

OAI22xp5_ASAP7_75t_L g2241 ( 
.A1(n_2150),
.A2(n_2031),
.B1(n_1959),
.B2(n_1986),
.Y(n_2241)
);

BUFx3_ASAP7_75t_L g2242 ( 
.A(n_2177),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2181),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2095),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_2104),
.B(n_2061),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_2120),
.Y(n_2246)
);

BUFx3_ASAP7_75t_L g2247 ( 
.A(n_2072),
.Y(n_2247)
);

BUFx8_ASAP7_75t_SL g2248 ( 
.A(n_2184),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_2078),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2125),
.B(n_2037),
.Y(n_2250)
);

BUFx3_ASAP7_75t_L g2251 ( 
.A(n_2158),
.Y(n_2251)
);

INVx2_ASAP7_75t_L g2252 ( 
.A(n_2110),
.Y(n_2252)
);

INVx8_ASAP7_75t_L g2253 ( 
.A(n_2139),
.Y(n_2253)
);

NAND2x1p5_ASAP7_75t_L g2254 ( 
.A(n_2192),
.B(n_2194),
.Y(n_2254)
);

OAI21x1_ASAP7_75t_L g2255 ( 
.A1(n_2244),
.A2(n_2136),
.B(n_2069),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2186),
.B(n_2183),
.Y(n_2256)
);

OR2x6_ASAP7_75t_L g2257 ( 
.A(n_2204),
.B(n_2074),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2186),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2205),
.Y(n_2259)
);

CKINVDCx20_ASAP7_75t_R g2260 ( 
.A(n_2233),
.Y(n_2260)
);

AOI22xp33_ASAP7_75t_L g2261 ( 
.A1(n_2241),
.A2(n_2122),
.B1(n_2140),
.B2(n_2130),
.Y(n_2261)
);

OA21x2_ASAP7_75t_L g2262 ( 
.A1(n_2208),
.A2(n_2068),
.B(n_2115),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2205),
.B(n_2187),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2188),
.Y(n_2264)
);

OAI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2244),
.A2(n_2102),
.B(n_2074),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2208),
.A2(n_2073),
.B(n_2132),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2236),
.B(n_2116),
.Y(n_2267)
);

INVx5_ASAP7_75t_L g2268 ( 
.A(n_2237),
.Y(n_2268)
);

AO21x2_ASAP7_75t_L g2269 ( 
.A1(n_2226),
.A2(n_2179),
.B(n_2148),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2238),
.A2(n_2089),
.B(n_2145),
.Y(n_2270)
);

CKINVDCx11_ASAP7_75t_R g2271 ( 
.A(n_2202),
.Y(n_2271)
);

CKINVDCx16_ASAP7_75t_R g2272 ( 
.A(n_2202),
.Y(n_2272)
);

AOI22xp33_ASAP7_75t_L g2273 ( 
.A1(n_2246),
.A2(n_2180),
.B1(n_2179),
.B2(n_2116),
.Y(n_2273)
);

OAI21x1_ASAP7_75t_SL g2274 ( 
.A1(n_2199),
.A2(n_2168),
.B(n_2082),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2196),
.Y(n_2275)
);

OR2x2_ASAP7_75t_L g2276 ( 
.A(n_2229),
.B(n_2153),
.Y(n_2276)
);

INVx2_ASAP7_75t_L g2277 ( 
.A(n_2213),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2213),
.Y(n_2278)
);

A2O1A1Ixp33_ASAP7_75t_L g2279 ( 
.A1(n_2193),
.A2(n_2162),
.B(n_2182),
.C(n_2131),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2217),
.Y(n_2280)
);

BUFx6f_ASAP7_75t_L g2281 ( 
.A(n_2206),
.Y(n_2281)
);

INVx2_ASAP7_75t_L g2282 ( 
.A(n_2217),
.Y(n_2282)
);

BUFx12f_ASAP7_75t_L g2283 ( 
.A(n_2216),
.Y(n_2283)
);

AOI22xp33_ASAP7_75t_L g2284 ( 
.A1(n_2246),
.A2(n_2124),
.B1(n_2099),
.B2(n_2151),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2193),
.A2(n_2170),
.B1(n_2085),
.B2(n_2134),
.Y(n_2285)
);

BUFx3_ASAP7_75t_L g2286 ( 
.A(n_2216),
.Y(n_2286)
);

INVx4_ASAP7_75t_L g2287 ( 
.A(n_2192),
.Y(n_2287)
);

AOI221xp5_ASAP7_75t_L g2288 ( 
.A1(n_2210),
.A2(n_2108),
.B1(n_2138),
.B2(n_1957),
.C(n_2052),
.Y(n_2288)
);

OAI21x1_ASAP7_75t_L g2289 ( 
.A1(n_2249),
.A2(n_2252),
.B(n_2231),
.Y(n_2289)
);

OAI211xp5_ASAP7_75t_SL g2290 ( 
.A1(n_2245),
.A2(n_2129),
.B(n_2126),
.C(n_1983),
.Y(n_2290)
);

AOI22xp33_ASAP7_75t_L g2291 ( 
.A1(n_2246),
.A2(n_2164),
.B1(n_2155),
.B2(n_2149),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2239),
.Y(n_2292)
);

NAND2xp5_ASAP7_75t_L g2293 ( 
.A(n_2232),
.B(n_2160),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2243),
.Y(n_2294)
);

NOR2xp33_ASAP7_75t_SL g2295 ( 
.A(n_2185),
.B(n_1924),
.Y(n_2295)
);

OAI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2233),
.A2(n_2085),
.B1(n_2169),
.B2(n_2101),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2243),
.Y(n_2297)
);

AOI22xp33_ASAP7_75t_SL g2298 ( 
.A1(n_2285),
.A2(n_2236),
.B1(n_2246),
.B2(n_2235),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_2261),
.A2(n_2236),
.B1(n_2251),
.B2(n_2248),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2264),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_2287),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2264),
.Y(n_2302)
);

AOI21x1_ASAP7_75t_L g2303 ( 
.A1(n_2267),
.A2(n_2234),
.B(n_2249),
.Y(n_2303)
);

BUFx10_ASAP7_75t_L g2304 ( 
.A(n_2281),
.Y(n_2304)
);

NAND2x1p5_ASAP7_75t_L g2305 ( 
.A(n_2268),
.B(n_2192),
.Y(n_2305)
);

NAND2x1p5_ASAP7_75t_L g2306 ( 
.A(n_2268),
.B(n_2192),
.Y(n_2306)
);

AOI21xp33_ASAP7_75t_SL g2307 ( 
.A1(n_2272),
.A2(n_2253),
.B(n_2207),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_2276),
.Y(n_2308)
);

OAI22xp33_ASAP7_75t_L g2309 ( 
.A1(n_2267),
.A2(n_2236),
.B1(n_2296),
.B2(n_2257),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2273),
.A2(n_2247),
.B1(n_2251),
.B2(n_2250),
.Y(n_2310)
);

INVxp33_ASAP7_75t_L g2311 ( 
.A(n_2271),
.Y(n_2311)
);

BUFx2_ASAP7_75t_L g2312 ( 
.A(n_2287),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2275),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2294),
.B(n_2218),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2275),
.Y(n_2315)
);

INVxp67_ASAP7_75t_SL g2316 ( 
.A(n_2277),
.Y(n_2316)
);

AOI21x1_ASAP7_75t_L g2317 ( 
.A1(n_2289),
.A2(n_2212),
.B(n_2240),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2277),
.Y(n_2318)
);

AOI22xp33_ASAP7_75t_SL g2319 ( 
.A1(n_2269),
.A2(n_2230),
.B1(n_2227),
.B2(n_2247),
.Y(n_2319)
);

AOI22xp33_ASAP7_75t_SL g2320 ( 
.A1(n_2269),
.A2(n_2230),
.B1(n_2227),
.B2(n_2219),
.Y(n_2320)
);

INVx3_ASAP7_75t_L g2321 ( 
.A(n_2268),
.Y(n_2321)
);

INVx3_ASAP7_75t_L g2322 ( 
.A(n_2268),
.Y(n_2322)
);

INVx3_ASAP7_75t_L g2323 ( 
.A(n_2268),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2308),
.B(n_2297),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2300),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_2318),
.Y(n_2326)
);

INVx3_ASAP7_75t_L g2327 ( 
.A(n_2321),
.Y(n_2327)
);

BUFx2_ASAP7_75t_L g2328 ( 
.A(n_2301),
.Y(n_2328)
);

INVx2_ASAP7_75t_SL g2329 ( 
.A(n_2304),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2299),
.A2(n_2279),
.B1(n_2284),
.B2(n_2291),
.Y(n_2330)
);

HB1xp67_ASAP7_75t_L g2331 ( 
.A(n_2308),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2300),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2317),
.A2(n_2289),
.B(n_2255),
.Y(n_2333)
);

OAI21x1_ASAP7_75t_L g2334 ( 
.A1(n_2327),
.A2(n_2303),
.B(n_2317),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2331),
.Y(n_2335)
);

OR2x2_ASAP7_75t_L g2336 ( 
.A(n_2324),
.B(n_2314),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2329),
.B(n_2311),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2328),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2328),
.Y(n_2339)
);

HB1xp67_ASAP7_75t_L g2340 ( 
.A(n_2325),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_2335),
.B(n_2310),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_2337),
.B(n_2283),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_2338),
.Y(n_2343)
);

AOI33xp33_ASAP7_75t_L g2344 ( 
.A1(n_2339),
.A2(n_2298),
.A3(n_2319),
.B1(n_2320),
.B2(n_2309),
.B3(n_2288),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2335),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2336),
.B(n_2329),
.Y(n_2346)
);

INVx3_ASAP7_75t_L g2347 ( 
.A(n_2338),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2334),
.Y(n_2348)
);

BUFx2_ASAP7_75t_L g2349 ( 
.A(n_2340),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2340),
.B(n_2327),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2342),
.B(n_2327),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2347),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2347),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2347),
.Y(n_2354)
);

AND2x2_ASAP7_75t_L g2355 ( 
.A(n_2342),
.B(n_2286),
.Y(n_2355)
);

INVx2_ASAP7_75t_SL g2356 ( 
.A(n_2342),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_2346),
.B(n_2286),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2345),
.B(n_2271),
.Y(n_2358)
);

AO21x2_ASAP7_75t_L g2359 ( 
.A1(n_2343),
.A2(n_2348),
.B(n_2350),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2343),
.B(n_2326),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2349),
.B(n_2326),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2352),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2352),
.Y(n_2363)
);

OA21x2_ASAP7_75t_L g2364 ( 
.A1(n_2353),
.A2(n_2348),
.B(n_2350),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2356),
.A2(n_2341),
.B(n_2330),
.Y(n_2365)
);

INVx2_ASAP7_75t_L g2366 ( 
.A(n_2359),
.Y(n_2366)
);

AOI21x1_ASAP7_75t_L g2367 ( 
.A1(n_2354),
.A2(n_2312),
.B(n_2301),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2359),
.Y(n_2368)
);

BUFx6f_ASAP7_75t_L g2369 ( 
.A(n_2358),
.Y(n_2369)
);

AND2x4_ASAP7_75t_L g2370 ( 
.A(n_2355),
.B(n_2312),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2369),
.A2(n_2351),
.B1(n_2357),
.B2(n_2361),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2365),
.B(n_2361),
.Y(n_2372)
);

OAI21xp5_ASAP7_75t_L g2373 ( 
.A1(n_2370),
.A2(n_2344),
.B(n_2279),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2366),
.Y(n_2374)
);

INVx2_ASAP7_75t_L g2375 ( 
.A(n_2374),
.Y(n_2375)
);

INVx2_ASAP7_75t_L g2376 ( 
.A(n_2372),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2371),
.B(n_2369),
.Y(n_2377)
);

OAI33xp33_ASAP7_75t_L g2378 ( 
.A1(n_2373),
.A2(n_2362),
.A3(n_2363),
.B1(n_2368),
.B2(n_2366),
.B3(n_2360),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2377),
.Y(n_2379)
);

INVx3_ASAP7_75t_L g2380 ( 
.A(n_2375),
.Y(n_2380)
);

INVx1_ASAP7_75t_L g2381 ( 
.A(n_2376),
.Y(n_2381)
);

NOR2x1p5_ASAP7_75t_L g2382 ( 
.A(n_2378),
.B(n_2369),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2376),
.B(n_2369),
.Y(n_2383)
);

AND2x2_ASAP7_75t_L g2384 ( 
.A(n_2376),
.B(n_2370),
.Y(n_2384)
);

A2O1A1Ixp33_ASAP7_75t_L g2385 ( 
.A1(n_2382),
.A2(n_2344),
.B(n_2368),
.C(n_2370),
.Y(n_2385)
);

AOI22xp5_ASAP7_75t_L g2386 ( 
.A1(n_2379),
.A2(n_2364),
.B1(n_2360),
.B2(n_2295),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2383),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2384),
.Y(n_2388)
);

INVxp67_ASAP7_75t_L g2389 ( 
.A(n_2380),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2381),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2381),
.B(n_2260),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2380),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2383),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2383),
.Y(n_2394)
);

NAND2xp5_ASAP7_75t_L g2395 ( 
.A(n_2387),
.B(n_2364),
.Y(n_2395)
);

HB1xp67_ASAP7_75t_L g2396 ( 
.A(n_2389),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2388),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2391),
.B(n_2364),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2394),
.B(n_2367),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2393),
.B(n_2367),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2392),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_2389),
.B(n_2260),
.Y(n_2402)
);

AND2x2_ASAP7_75t_L g2403 ( 
.A(n_2390),
.B(n_2190),
.Y(n_2403)
);

HB1xp67_ASAP7_75t_L g2404 ( 
.A(n_2386),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2385),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2388),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2391),
.B(n_2248),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2395),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2402),
.B(n_1956),
.Y(n_2409)
);

OAI222xp33_ASAP7_75t_L g2410 ( 
.A1(n_2405),
.A2(n_2322),
.B1(n_2323),
.B2(n_2321),
.C1(n_2303),
.C2(n_2305),
.Y(n_2410)
);

O2A1O1Ixp33_ASAP7_75t_L g2411 ( 
.A1(n_2395),
.A2(n_2033),
.B(n_1991),
.C(n_2002),
.Y(n_2411)
);

NAND2xp5_ASAP7_75t_L g2412 ( 
.A(n_2400),
.B(n_2325),
.Y(n_2412)
);

OR2x2_ASAP7_75t_L g2413 ( 
.A(n_2402),
.B(n_2203),
.Y(n_2413)
);

OAI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_2407),
.A2(n_2283),
.B1(n_2322),
.B2(n_2321),
.Y(n_2414)
);

OR2x2_ASAP7_75t_L g2415 ( 
.A(n_2397),
.B(n_2406),
.Y(n_2415)
);

AOI32xp33_ASAP7_75t_L g2416 ( 
.A1(n_2399),
.A2(n_2290),
.A3(n_2211),
.B1(n_2203),
.B2(n_1987),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2398),
.B(n_2332),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2404),
.A2(n_2191),
.B1(n_2322),
.B2(n_2321),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2396),
.Y(n_2419)
);

OAI21xp33_ASAP7_75t_L g2420 ( 
.A1(n_2401),
.A2(n_2293),
.B(n_2191),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2403),
.B(n_2200),
.Y(n_2421)
);

OAI322xp33_ASAP7_75t_L g2422 ( 
.A1(n_2405),
.A2(n_1937),
.A3(n_2113),
.B1(n_2062),
.B2(n_2056),
.C1(n_2223),
.C2(n_2166),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_2419),
.B(n_2307),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_2415),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2421),
.B(n_2332),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2409),
.B(n_2224),
.Y(n_2426)
);

INVx1_ASAP7_75t_L g2427 ( 
.A(n_2408),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2413),
.Y(n_2428)
);

NOR2xp33_ASAP7_75t_L g2429 ( 
.A(n_2420),
.B(n_2414),
.Y(n_2429)
);

AOI22xp33_ASAP7_75t_L g2430 ( 
.A1(n_2418),
.A2(n_2219),
.B1(n_2281),
.B2(n_2322),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2412),
.B(n_2307),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2416),
.B(n_2197),
.Y(n_2432)
);

OAI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2411),
.A2(n_2005),
.B(n_2144),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2417),
.Y(n_2434)
);

AOI22xp33_ASAP7_75t_SL g2435 ( 
.A1(n_2410),
.A2(n_1945),
.B1(n_1916),
.B2(n_2323),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2422),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_2423),
.B(n_2242),
.Y(n_2437)
);

HB1xp67_ASAP7_75t_L g2438 ( 
.A(n_2424),
.Y(n_2438)
);

OR2x2_ASAP7_75t_L g2439 ( 
.A(n_2428),
.B(n_147),
.Y(n_2439)
);

OR2x2_ASAP7_75t_L g2440 ( 
.A(n_2432),
.B(n_148),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2427),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2431),
.B(n_2436),
.Y(n_2442)
);

INVxp67_ASAP7_75t_L g2443 ( 
.A(n_2429),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2426),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2434),
.B(n_2242),
.Y(n_2445)
);

AND2x2_ASAP7_75t_L g2446 ( 
.A(n_2435),
.B(n_2219),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2425),
.Y(n_2447)
);

INVxp67_ASAP7_75t_L g2448 ( 
.A(n_2433),
.Y(n_2448)
);

AOI22xp33_ASAP7_75t_L g2449 ( 
.A1(n_2430),
.A2(n_2219),
.B1(n_2323),
.B2(n_2281),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2433),
.B(n_2323),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2424),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2423),
.B(n_2304),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2424),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_2424),
.B(n_148),
.Y(n_2454)
);

NOR2xp33_ASAP7_75t_L g2455 ( 
.A(n_2424),
.B(n_149),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2423),
.B(n_2333),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2423),
.B(n_2333),
.Y(n_2457)
);

AND2x4_ASAP7_75t_SL g2458 ( 
.A(n_2424),
.B(n_1916),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2438),
.B(n_149),
.Y(n_2459)
);

NOR2xp33_ASAP7_75t_L g2460 ( 
.A(n_2453),
.B(n_150),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2451),
.B(n_151),
.Y(n_2461)
);

NAND4xp25_ASAP7_75t_L g2462 ( 
.A(n_2443),
.B(n_1939),
.C(n_2046),
.D(n_2105),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2439),
.B(n_152),
.Y(n_2463)
);

OAI211xp5_ASAP7_75t_L g2464 ( 
.A1(n_2441),
.A2(n_1945),
.B(n_2027),
.C(n_2038),
.Y(n_2464)
);

INVx1_ASAP7_75t_SL g2465 ( 
.A(n_2454),
.Y(n_2465)
);

OAI21xp5_ASAP7_75t_SL g2466 ( 
.A1(n_2442),
.A2(n_1945),
.B(n_1988),
.Y(n_2466)
);

NOR2xp33_ASAP7_75t_L g2467 ( 
.A(n_2455),
.B(n_2440),
.Y(n_2467)
);

OAI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_2449),
.A2(n_2305),
.B1(n_2306),
.B2(n_2281),
.Y(n_2468)
);

BUFx2_ASAP7_75t_L g2469 ( 
.A(n_2441),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2452),
.B(n_152),
.Y(n_2470)
);

NAND4xp25_ASAP7_75t_L g2471 ( 
.A(n_2444),
.B(n_2014),
.C(n_2019),
.D(n_1974),
.Y(n_2471)
);

OAI211xp5_ASAP7_75t_L g2472 ( 
.A1(n_2448),
.A2(n_2051),
.B(n_2050),
.C(n_2026),
.Y(n_2472)
);

NAND2x1_ASAP7_75t_L g2473 ( 
.A(n_2446),
.B(n_2020),
.Y(n_2473)
);

INVxp67_ASAP7_75t_SL g2474 ( 
.A(n_2458),
.Y(n_2474)
);

NAND3xp33_ASAP7_75t_L g2475 ( 
.A(n_2447),
.B(n_2019),
.C(n_2014),
.Y(n_2475)
);

NOR3x1_ASAP7_75t_L g2476 ( 
.A(n_2445),
.B(n_153),
.C(n_154),
.Y(n_2476)
);

NOR2x1_ASAP7_75t_L g2477 ( 
.A(n_2450),
.B(n_153),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2437),
.B(n_2304),
.Y(n_2478)
);

NOR3xp33_ASAP7_75t_L g2479 ( 
.A(n_2456),
.B(n_2117),
.C(n_2028),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2457),
.B(n_155),
.Y(n_2480)
);

NAND2x1_ASAP7_75t_L g2481 ( 
.A(n_2453),
.B(n_2020),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_L g2482 ( 
.A(n_2454),
.B(n_156),
.Y(n_2482)
);

NAND3xp33_ASAP7_75t_L g2483 ( 
.A(n_2438),
.B(n_2026),
.C(n_2020),
.Y(n_2483)
);

NOR2xp67_ASAP7_75t_L g2484 ( 
.A(n_2438),
.B(n_156),
.Y(n_2484)
);

INVxp33_ASAP7_75t_SL g2485 ( 
.A(n_2438),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2438),
.B(n_157),
.Y(n_2486)
);

NAND4xp25_ASAP7_75t_L g2487 ( 
.A(n_2443),
.B(n_2060),
.C(n_2032),
.D(n_2103),
.Y(n_2487)
);

AOI221xp5_ASAP7_75t_L g2488 ( 
.A1(n_2443),
.A2(n_2121),
.B1(n_2157),
.B2(n_2161),
.C(n_2159),
.Y(n_2488)
);

NOR2xp33_ASAP7_75t_L g2489 ( 
.A(n_2438),
.B(n_157),
.Y(n_2489)
);

AOI21xp5_ASAP7_75t_L g2490 ( 
.A1(n_2438),
.A2(n_2100),
.B(n_2146),
.Y(n_2490)
);

AOI211x1_ASAP7_75t_L g2491 ( 
.A1(n_2451),
.A2(n_2152),
.B(n_2094),
.C(n_2012),
.Y(n_2491)
);

NAND3xp33_ASAP7_75t_SL g2492 ( 
.A(n_2438),
.B(n_2063),
.C(n_2013),
.Y(n_2492)
);

INVx1_ASAP7_75t_L g2493 ( 
.A(n_2438),
.Y(n_2493)
);

NAND3xp33_ASAP7_75t_SL g2494 ( 
.A(n_2438),
.B(n_2306),
.C(n_2305),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2454),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2484),
.B(n_158),
.Y(n_2496)
);

AOI211xp5_ASAP7_75t_L g2497 ( 
.A1(n_2459),
.A2(n_2067),
.B(n_2026),
.C(n_160),
.Y(n_2497)
);

NAND4xp25_ASAP7_75t_SL g2498 ( 
.A(n_2493),
.B(n_2017),
.C(n_2088),
.D(n_160),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2486),
.B(n_158),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2485),
.A2(n_2469),
.B(n_2474),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2482),
.Y(n_2501)
);

NAND4xp75_ASAP7_75t_L g2502 ( 
.A(n_2477),
.B(n_162),
.C(n_159),
.D(n_161),
.Y(n_2502)
);

AND4x1_ASAP7_75t_L g2503 ( 
.A(n_2489),
.B(n_163),
.C(n_159),
.D(n_161),
.Y(n_2503)
);

AOI211xp5_ASAP7_75t_SL g2504 ( 
.A1(n_2470),
.A2(n_2467),
.B(n_2480),
.C(n_2463),
.Y(n_2504)
);

OAI22xp5_ASAP7_75t_L g2505 ( 
.A1(n_2483),
.A2(n_2306),
.B1(n_2067),
.B2(n_2221),
.Y(n_2505)
);

NAND3xp33_ASAP7_75t_L g2506 ( 
.A(n_2495),
.B(n_2067),
.C(n_163),
.Y(n_2506)
);

INVxp67_ASAP7_75t_L g2507 ( 
.A(n_2461),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_L g2508 ( 
.A(n_2460),
.B(n_164),
.Y(n_2508)
);

NOR4xp75_ASAP7_75t_L g2509 ( 
.A(n_2473),
.B(n_167),
.C(n_165),
.D(n_166),
.Y(n_2509)
);

NAND4xp25_ASAP7_75t_L g2510 ( 
.A(n_2476),
.B(n_2049),
.C(n_167),
.D(n_165),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_2478),
.B(n_2304),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_2481),
.Y(n_2512)
);

AND2x2_ASAP7_75t_L g2513 ( 
.A(n_2465),
.B(n_2316),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2475),
.B(n_166),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_L g2515 ( 
.A(n_2466),
.B(n_168),
.C(n_169),
.Y(n_2515)
);

INVxp67_ASAP7_75t_L g2516 ( 
.A(n_2472),
.Y(n_2516)
);

NOR4xp25_ASAP7_75t_L g2517 ( 
.A(n_2494),
.B(n_170),
.C(n_168),
.D(n_169),
.Y(n_2517)
);

NAND2xp33_ASAP7_75t_SL g2518 ( 
.A(n_2468),
.B(n_2189),
.Y(n_2518)
);

NOR3xp33_ASAP7_75t_SL g2519 ( 
.A(n_2490),
.B(n_2464),
.C(n_2492),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2487),
.B(n_170),
.C(n_171),
.Y(n_2520)
);

NOR3xp33_ASAP7_75t_L g2521 ( 
.A(n_2462),
.B(n_171),
.C(n_172),
.Y(n_2521)
);

OR2x2_ASAP7_75t_L g2522 ( 
.A(n_2479),
.B(n_172),
.Y(n_2522)
);

AOI21xp5_ASAP7_75t_L g2523 ( 
.A1(n_2488),
.A2(n_2471),
.B(n_2491),
.Y(n_2523)
);

NOR2xp67_ASAP7_75t_SL g2524 ( 
.A(n_2493),
.B(n_2198),
.Y(n_2524)
);

A2O1A1Ixp33_ASAP7_75t_L g2525 ( 
.A1(n_2484),
.A2(n_2135),
.B(n_2201),
.C(n_175),
.Y(n_2525)
);

NOR2xp33_ASAP7_75t_SL g2526 ( 
.A(n_2485),
.B(n_2198),
.Y(n_2526)
);

AND4x1_ASAP7_75t_L g2527 ( 
.A(n_2459),
.B(n_176),
.C(n_173),
.D(n_174),
.Y(n_2527)
);

AOI22xp33_ASAP7_75t_L g2528 ( 
.A1(n_2485),
.A2(n_2221),
.B1(n_2287),
.B2(n_2189),
.Y(n_2528)
);

NAND4xp25_ASAP7_75t_L g2529 ( 
.A(n_2485),
.B(n_177),
.C(n_174),
.D(n_176),
.Y(n_2529)
);

INVx1_ASAP7_75t_SL g2530 ( 
.A(n_2469),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2493),
.B(n_177),
.Y(n_2531)
);

NOR4xp75_ASAP7_75t_L g2532 ( 
.A(n_2480),
.B(n_180),
.C(n_178),
.D(n_179),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2484),
.B(n_178),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2530),
.B(n_180),
.Y(n_2534)
);

INVx1_ASAP7_75t_L g2535 ( 
.A(n_2531),
.Y(n_2535)
);

AOI32xp33_ASAP7_75t_L g2536 ( 
.A1(n_2526),
.A2(n_2096),
.A3(n_2118),
.B1(n_2231),
.B2(n_2112),
.Y(n_2536)
);

OAI211xp5_ASAP7_75t_SL g2537 ( 
.A1(n_2500),
.A2(n_183),
.B(n_181),
.C(n_182),
.Y(n_2537)
);

NAND2x1_ASAP7_75t_L g2538 ( 
.A(n_2501),
.B(n_2524),
.Y(n_2538)
);

OAI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2496),
.A2(n_2201),
.B1(n_2194),
.B2(n_2135),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2502),
.Y(n_2540)
);

NOR2x1_ASAP7_75t_L g2541 ( 
.A(n_2529),
.B(n_181),
.Y(n_2541)
);

O2A1O1Ixp33_ASAP7_75t_L g2542 ( 
.A1(n_2533),
.A2(n_2512),
.B(n_2499),
.C(n_2516),
.Y(n_2542)
);

INVxp67_ASAP7_75t_SL g2543 ( 
.A(n_2503),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2527),
.Y(n_2544)
);

OAI211xp5_ASAP7_75t_SL g2545 ( 
.A1(n_2504),
.A2(n_184),
.B(n_182),
.C(n_183),
.Y(n_2545)
);

NAND3xp33_ASAP7_75t_L g2546 ( 
.A(n_2506),
.B(n_184),
.C(n_185),
.Y(n_2546)
);

OR2x2_ASAP7_75t_L g2547 ( 
.A(n_2517),
.B(n_185),
.Y(n_2547)
);

NOR2x1_ASAP7_75t_L g2548 ( 
.A(n_2508),
.B(n_186),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2511),
.B(n_186),
.Y(n_2549)
);

AOI22xp5_ASAP7_75t_L g2550 ( 
.A1(n_2513),
.A2(n_2521),
.B1(n_2510),
.B2(n_2498),
.Y(n_2550)
);

NOR2xp67_ASAP7_75t_L g2551 ( 
.A(n_2515),
.B(n_187),
.Y(n_2551)
);

XNOR2xp5_ASAP7_75t_L g2552 ( 
.A(n_2532),
.B(n_2509),
.Y(n_2552)
);

AOI32xp33_ASAP7_75t_L g2553 ( 
.A1(n_2518),
.A2(n_2172),
.A3(n_2154),
.B1(n_2215),
.B2(n_189),
.Y(n_2553)
);

OAI332xp33_ASAP7_75t_L g2554 ( 
.A1(n_2514),
.A2(n_187),
.A3(n_188),
.B1(n_190),
.B2(n_191),
.B3(n_192),
.C1(n_193),
.C2(n_194),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2507),
.B(n_2302),
.Y(n_2555)
);

INVx1_ASAP7_75t_SL g2556 ( 
.A(n_2522),
.Y(n_2556)
);

AOI31xp33_ASAP7_75t_L g2557 ( 
.A1(n_2497),
.A2(n_2254),
.A3(n_192),
.B(n_188),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2520),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2525),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2519),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2523),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2528),
.Y(n_2562)
);

OR2x2_ASAP7_75t_L g2563 ( 
.A(n_2505),
.B(n_190),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2531),
.Y(n_2564)
);

INVxp67_ASAP7_75t_L g2565 ( 
.A(n_2526),
.Y(n_2565)
);

OR2x2_ASAP7_75t_L g2566 ( 
.A(n_2517),
.B(n_193),
.Y(n_2566)
);

XNOR2x2_ASAP7_75t_L g2567 ( 
.A(n_2530),
.B(n_194),
.Y(n_2567)
);

AOI22xp5_ASAP7_75t_L g2568 ( 
.A1(n_2526),
.A2(n_2206),
.B1(n_2189),
.B2(n_2253),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2531),
.Y(n_2569)
);

INVxp67_ASAP7_75t_L g2570 ( 
.A(n_2526),
.Y(n_2570)
);

NAND4xp25_ASAP7_75t_L g2571 ( 
.A(n_2500),
.B(n_197),
.C(n_195),
.D(n_196),
.Y(n_2571)
);

AOI221xp5_ASAP7_75t_L g2572 ( 
.A1(n_2517),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.C(n_198),
.Y(n_2572)
);

A2O1A1Ixp33_ASAP7_75t_L g2573 ( 
.A1(n_2500),
.A2(n_202),
.B(n_199),
.C(n_201),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2531),
.Y(n_2574)
);

XNOR2x2_ASAP7_75t_L g2575 ( 
.A(n_2530),
.B(n_202),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2531),
.Y(n_2576)
);

OAI21xp5_ASAP7_75t_L g2577 ( 
.A1(n_2500),
.A2(n_2270),
.B(n_2265),
.Y(n_2577)
);

AOI322xp5_ASAP7_75t_L g2578 ( 
.A1(n_2530),
.A2(n_2220),
.A3(n_2253),
.B1(n_2143),
.B2(n_2302),
.C1(n_2313),
.C2(n_2315),
.Y(n_2578)
);

NOR2xp33_ASAP7_75t_L g2579 ( 
.A(n_2529),
.B(n_203),
.Y(n_2579)
);

AOI221xp5_ASAP7_75t_L g2580 ( 
.A1(n_2517),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.C(n_207),
.Y(n_2580)
);

OAI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2500),
.A2(n_2270),
.B(n_2265),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2530),
.B(n_204),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2509),
.Y(n_2583)
);

NOR2x1_ASAP7_75t_L g2584 ( 
.A(n_2502),
.B(n_206),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2531),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2530),
.B(n_2189),
.Y(n_2586)
);

AOI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2500),
.A2(n_207),
.B(n_208),
.Y(n_2587)
);

OA22x2_ASAP7_75t_L g2588 ( 
.A1(n_2530),
.A2(n_2274),
.B1(n_2209),
.B2(n_2318),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2501),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2531),
.Y(n_2590)
);

XNOR2x1_ASAP7_75t_L g2591 ( 
.A(n_2532),
.B(n_208),
.Y(n_2591)
);

AOI21xp5_ASAP7_75t_L g2592 ( 
.A1(n_2500),
.A2(n_209),
.B(n_210),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2531),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_2530),
.B(n_209),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2531),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_SL g2596 ( 
.A(n_2530),
.B(n_2206),
.Y(n_2596)
);

OAI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2528),
.A2(n_2254),
.B1(n_2194),
.B2(n_2206),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2547),
.Y(n_2598)
);

NOR4xp25_ASAP7_75t_L g2599 ( 
.A(n_2542),
.B(n_213),
.C(n_211),
.D(n_212),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2566),
.Y(n_2600)
);

NOR2x1_ASAP7_75t_L g2601 ( 
.A(n_2571),
.B(n_211),
.Y(n_2601)
);

INVx1_ASAP7_75t_L g2602 ( 
.A(n_2591),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_SL g2603 ( 
.A(n_2572),
.B(n_2194),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2583),
.B(n_212),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2580),
.B(n_213),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2567),
.Y(n_2606)
);

AO211x2_ASAP7_75t_L g2607 ( 
.A1(n_2546),
.A2(n_216),
.B(n_214),
.C(n_215),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2552),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2575),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_2587),
.B(n_214),
.Y(n_2610)
);

AOI22xp5_ASAP7_75t_L g2611 ( 
.A1(n_2579),
.A2(n_2215),
.B1(n_2222),
.B2(n_2257),
.Y(n_2611)
);

NOR2x1_ASAP7_75t_L g2612 ( 
.A(n_2548),
.B(n_2584),
.Y(n_2612)
);

AOI221xp5_ASAP7_75t_L g2613 ( 
.A1(n_2557),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.C(n_220),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2589),
.Y(n_2614)
);

AOI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2560),
.A2(n_2222),
.B1(n_2257),
.B2(n_2292),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2534),
.Y(n_2616)
);

AOI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2543),
.A2(n_2222),
.B1(n_2257),
.B2(n_2313),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2582),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_2565),
.A2(n_2222),
.B1(n_2315),
.B2(n_2209),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_SL g2620 ( 
.A(n_2551),
.B(n_2594),
.Y(n_2620)
);

NOR4xp25_ASAP7_75t_L g2621 ( 
.A(n_2570),
.B(n_221),
.C(n_217),
.D(n_220),
.Y(n_2621)
);

NOR2xp33_ASAP7_75t_L g2622 ( 
.A(n_2537),
.B(n_222),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2549),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2592),
.B(n_222),
.Y(n_2624)
);

AO22x2_ASAP7_75t_L g2625 ( 
.A1(n_2540),
.A2(n_225),
.B1(n_223),
.B2(n_224),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2541),
.Y(n_2626)
);

AOI22xp33_ASAP7_75t_SL g2627 ( 
.A1(n_2561),
.A2(n_2209),
.B1(n_2237),
.B2(n_227),
.Y(n_2627)
);

OA22x2_ASAP7_75t_L g2628 ( 
.A1(n_2550),
.A2(n_228),
.B1(n_223),
.B2(n_225),
.Y(n_2628)
);

AOI221xp5_ASAP7_75t_L g2629 ( 
.A1(n_2596),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.C(n_231),
.Y(n_2629)
);

NOR2x1_ASAP7_75t_L g2630 ( 
.A(n_2545),
.B(n_230),
.Y(n_2630)
);

NOR2x1_ASAP7_75t_L g2631 ( 
.A(n_2573),
.B(n_232),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2544),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2554),
.B(n_232),
.Y(n_2633)
);

AOI31xp33_ASAP7_75t_L g2634 ( 
.A1(n_2535),
.A2(n_235),
.A3(n_233),
.B(n_234),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2569),
.Y(n_2635)
);

AOI22xp5_ASAP7_75t_L g2636 ( 
.A1(n_2586),
.A2(n_2195),
.B1(n_2240),
.B2(n_2228),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2538),
.Y(n_2637)
);

AO22x1_ASAP7_75t_L g2638 ( 
.A1(n_2559),
.A2(n_237),
.B1(n_233),
.B2(n_236),
.Y(n_2638)
);

AOI22xp5_ASAP7_75t_L g2639 ( 
.A1(n_2551),
.A2(n_2195),
.B1(n_2228),
.B2(n_2256),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2563),
.Y(n_2640)
);

NOR2xp33_ASAP7_75t_L g2641 ( 
.A(n_2564),
.B(n_238),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2574),
.Y(n_2642)
);

NOR2x1_ASAP7_75t_L g2643 ( 
.A(n_2576),
.B(n_238),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2585),
.Y(n_2644)
);

AO22x2_ASAP7_75t_L g2645 ( 
.A1(n_2590),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2593),
.Y(n_2646)
);

NOR3xp33_ASAP7_75t_L g2647 ( 
.A(n_2558),
.B(n_239),
.C(n_240),
.Y(n_2647)
);

NOR2x1_ASAP7_75t_L g2648 ( 
.A(n_2595),
.B(n_2562),
.Y(n_2648)
);

NOR2x1_ASAP7_75t_L g2649 ( 
.A(n_2556),
.B(n_242),
.Y(n_2649)
);

BUFx3_ASAP7_75t_L g2650 ( 
.A(n_2555),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2568),
.B(n_243),
.Y(n_2651)
);

AO22x2_ASAP7_75t_L g2652 ( 
.A1(n_2597),
.A2(n_246),
.B1(n_243),
.B2(n_244),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2588),
.Y(n_2653)
);

AOI22xp5_ASAP7_75t_L g2654 ( 
.A1(n_2539),
.A2(n_2581),
.B1(n_2577),
.B2(n_2553),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2578),
.Y(n_2655)
);

AOI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_2536),
.A2(n_2228),
.B1(n_2256),
.B2(n_2237),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2547),
.Y(n_2657)
);

NOR2x1_ASAP7_75t_L g2658 ( 
.A(n_2571),
.B(n_244),
.Y(n_2658)
);

NOR2x1_ASAP7_75t_L g2659 ( 
.A(n_2571),
.B(n_246),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2572),
.B(n_247),
.Y(n_2660)
);

AOI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2579),
.A2(n_2228),
.B1(n_2237),
.B2(n_2262),
.Y(n_2661)
);

AOI22xp5_ASAP7_75t_L g2662 ( 
.A1(n_2579),
.A2(n_2262),
.B1(n_2280),
.B2(n_2278),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2547),
.Y(n_2663)
);

AOI221xp5_ASAP7_75t_L g2664 ( 
.A1(n_2557),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.C(n_251),
.Y(n_2664)
);

AOI221xp5_ASAP7_75t_L g2665 ( 
.A1(n_2557),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.C(n_253),
.Y(n_2665)
);

OA22x2_ASAP7_75t_L g2666 ( 
.A1(n_2550),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_SL g2667 ( 
.A(n_2572),
.B(n_254),
.Y(n_2667)
);

OAI22x1_ASAP7_75t_L g2668 ( 
.A1(n_2552),
.A2(n_257),
.B1(n_255),
.B2(n_256),
.Y(n_2668)
);

AOI22xp5_ASAP7_75t_L g2669 ( 
.A1(n_2579),
.A2(n_2262),
.B1(n_2088),
.B2(n_2225),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2614),
.B(n_2263),
.Y(n_2670)
);

NOR2x1_ASAP7_75t_L g2671 ( 
.A(n_2643),
.B(n_255),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2599),
.B(n_256),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2621),
.B(n_258),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2604),
.B(n_258),
.Y(n_2674)
);

NOR4xp75_ASAP7_75t_L g2675 ( 
.A(n_2633),
.B(n_261),
.C(n_259),
.D(n_260),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2649),
.B(n_259),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2647),
.B(n_260),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2637),
.B(n_261),
.Y(n_2678)
);

AND2x2_ASAP7_75t_L g2679 ( 
.A(n_2630),
.B(n_2263),
.Y(n_2679)
);

CKINVDCx20_ASAP7_75t_R g2680 ( 
.A(n_2608),
.Y(n_2680)
);

NOR3xp33_ASAP7_75t_L g2681 ( 
.A(n_2648),
.B(n_262),
.C(n_263),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2628),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2666),
.Y(n_2683)
);

OR2x2_ASAP7_75t_L g2684 ( 
.A(n_2610),
.B(n_262),
.Y(n_2684)
);

INVx2_ASAP7_75t_L g2685 ( 
.A(n_2645),
.Y(n_2685)
);

AOI22xp33_ASAP7_75t_L g2686 ( 
.A1(n_2606),
.A2(n_2214),
.B1(n_2282),
.B2(n_2252),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2624),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2607),
.Y(n_2688)
);

OAI21xp5_ASAP7_75t_L g2689 ( 
.A1(n_2622),
.A2(n_2266),
.B(n_263),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2613),
.B(n_264),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2601),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2658),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2664),
.B(n_264),
.Y(n_2693)
);

NAND3xp33_ASAP7_75t_L g2694 ( 
.A(n_2665),
.B(n_265),
.C(n_266),
.Y(n_2694)
);

NAND3xp33_ASAP7_75t_L g2695 ( 
.A(n_2629),
.B(n_265),
.C(n_266),
.Y(n_2695)
);

NOR2x1p5_ASAP7_75t_L g2696 ( 
.A(n_2635),
.B(n_2602),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2638),
.B(n_267),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_L g2698 ( 
.A(n_2609),
.B(n_267),
.Y(n_2698)
);

OAI22xp5_ASAP7_75t_L g2699 ( 
.A1(n_2639),
.A2(n_2259),
.B1(n_2258),
.B2(n_2282),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_SL g2700 ( 
.A(n_2642),
.B(n_268),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2620),
.A2(n_268),
.B(n_269),
.Y(n_2701)
);

NOR3x1_ASAP7_75t_L g2702 ( 
.A(n_2605),
.B(n_269),
.C(n_270),
.Y(n_2702)
);

NOR3xp33_ASAP7_75t_SL g2703 ( 
.A(n_2644),
.B(n_271),
.C(n_272),
.Y(n_2703)
);

INVxp67_ASAP7_75t_L g2704 ( 
.A(n_2641),
.Y(n_2704)
);

INVx1_ASAP7_75t_SL g2705 ( 
.A(n_2668),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2634),
.B(n_271),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2659),
.B(n_273),
.Y(n_2707)
);

NAND3xp33_ASAP7_75t_L g2708 ( 
.A(n_2612),
.B(n_273),
.C(n_274),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2625),
.Y(n_2709)
);

OAI21xp5_ASAP7_75t_SL g2710 ( 
.A1(n_2627),
.A2(n_274),
.B(n_275),
.Y(n_2710)
);

NAND3xp33_ASAP7_75t_SL g2711 ( 
.A(n_2626),
.B(n_275),
.C(n_276),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2646),
.B(n_276),
.Y(n_2712)
);

NAND3xp33_ASAP7_75t_L g2713 ( 
.A(n_2632),
.B(n_277),
.C(n_278),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2598),
.B(n_278),
.Y(n_2714)
);

AOI211xp5_ASAP7_75t_SL g2715 ( 
.A1(n_2600),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2625),
.Y(n_2716)
);

INVx1_ASAP7_75t_L g2717 ( 
.A(n_2631),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2645),
.Y(n_2718)
);

NAND3xp33_ASAP7_75t_L g2719 ( 
.A(n_2653),
.B(n_279),
.C(n_280),
.Y(n_2719)
);

OR2x2_ASAP7_75t_L g2720 ( 
.A(n_2651),
.B(n_283),
.Y(n_2720)
);

OAI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2611),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2657),
.B(n_284),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2663),
.B(n_285),
.Y(n_2723)
);

NOR2x1_ASAP7_75t_L g2724 ( 
.A(n_2650),
.B(n_2640),
.Y(n_2724)
);

AOI221xp5_ASAP7_75t_L g2725 ( 
.A1(n_2652),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.C(n_292),
.Y(n_2725)
);

INVxp67_ASAP7_75t_L g2726 ( 
.A(n_2652),
.Y(n_2726)
);

NOR3xp33_ASAP7_75t_L g2727 ( 
.A(n_2616),
.B(n_289),
.C(n_290),
.Y(n_2727)
);

NOR3xp33_ASAP7_75t_L g2728 ( 
.A(n_2618),
.B(n_291),
.C(n_293),
.Y(n_2728)
);

INVxp67_ASAP7_75t_L g2729 ( 
.A(n_2660),
.Y(n_2729)
);

OAI22xp5_ASAP7_75t_L g2730 ( 
.A1(n_2619),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_2730)
);

NAND3xp33_ASAP7_75t_L g2731 ( 
.A(n_2655),
.B(n_294),
.C(n_297),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2623),
.B(n_297),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2603),
.B(n_298),
.Y(n_2733)
);

OR2x2_ASAP7_75t_L g2734 ( 
.A(n_2667),
.B(n_298),
.Y(n_2734)
);

NAND2xp33_ASAP7_75t_SL g2735 ( 
.A(n_2654),
.B(n_2656),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2712),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2671),
.Y(n_2737)
);

NOR3xp33_ASAP7_75t_L g2738 ( 
.A(n_2724),
.B(n_2661),
.C(n_2662),
.Y(n_2738)
);

NAND4xp75_ASAP7_75t_L g2739 ( 
.A(n_2698),
.B(n_2669),
.C(n_2636),
.D(n_2615),
.Y(n_2739)
);

NOR3xp33_ASAP7_75t_L g2740 ( 
.A(n_2735),
.B(n_2617),
.C(n_299),
.Y(n_2740)
);

OAI211xp5_ASAP7_75t_L g2741 ( 
.A1(n_2697),
.A2(n_300),
.B(n_301),
.C(n_302),
.Y(n_2741)
);

NOR2x1p5_ASAP7_75t_L g2742 ( 
.A(n_2711),
.B(n_301),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2696),
.Y(n_2743)
);

OR2x2_ASAP7_75t_L g2744 ( 
.A(n_2673),
.B(n_302),
.Y(n_2744)
);

NAND3xp33_ASAP7_75t_SL g2745 ( 
.A(n_2680),
.B(n_303),
.C(n_304),
.Y(n_2745)
);

OAI211xp5_ASAP7_75t_L g2746 ( 
.A1(n_2672),
.A2(n_303),
.B(n_304),
.C(n_306),
.Y(n_2746)
);

NAND3xp33_ASAP7_75t_SL g2747 ( 
.A(n_2681),
.B(n_306),
.C(n_307),
.Y(n_2747)
);

INVx2_ASAP7_75t_SL g2748 ( 
.A(n_2674),
.Y(n_2748)
);

NAND4xp75_ASAP7_75t_L g2749 ( 
.A(n_2702),
.B(n_309),
.C(n_311),
.D(n_312),
.Y(n_2749)
);

NAND3xp33_ASAP7_75t_SL g2750 ( 
.A(n_2675),
.B(n_309),
.C(n_311),
.Y(n_2750)
);

NOR2xp33_ASAP7_75t_L g2751 ( 
.A(n_2706),
.B(n_312),
.Y(n_2751)
);

OAI211xp5_ASAP7_75t_L g2752 ( 
.A1(n_2710),
.A2(n_313),
.B(n_314),
.C(n_315),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2727),
.B(n_313),
.Y(n_2753)
);

NOR5xp2_ASAP7_75t_L g2754 ( 
.A(n_2726),
.B(n_314),
.C(n_315),
.D(n_316),
.E(n_317),
.Y(n_2754)
);

INVx4_ASAP7_75t_L g2755 ( 
.A(n_2707),
.Y(n_2755)
);

NOR3xp33_ASAP7_75t_L g2756 ( 
.A(n_2717),
.B(n_317),
.C(n_318),
.Y(n_2756)
);

AND2x4_ASAP7_75t_L g2757 ( 
.A(n_2679),
.B(n_318),
.Y(n_2757)
);

NOR2x1_ASAP7_75t_L g2758 ( 
.A(n_2708),
.B(n_319),
.Y(n_2758)
);

AOI22xp5_ASAP7_75t_SL g2759 ( 
.A1(n_2688),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_2759)
);

AND4x1_ASAP7_75t_L g2760 ( 
.A(n_2731),
.B(n_2703),
.C(n_2719),
.D(n_2715),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2728),
.B(n_320),
.Y(n_2761)
);

NAND3xp33_ASAP7_75t_L g2762 ( 
.A(n_2725),
.B(n_2733),
.C(n_2701),
.Y(n_2762)
);

NOR2x1_ASAP7_75t_L g2763 ( 
.A(n_2708),
.B(n_321),
.Y(n_2763)
);

NAND4xp25_ASAP7_75t_L g2764 ( 
.A(n_2694),
.B(n_322),
.C(n_323),
.D(n_324),
.Y(n_2764)
);

NOR2x1_ASAP7_75t_L g2765 ( 
.A(n_2718),
.B(n_322),
.Y(n_2765)
);

NOR3xp33_ASAP7_75t_L g2766 ( 
.A(n_2691),
.B(n_323),
.C(n_325),
.Y(n_2766)
);

NOR2x1p5_ASAP7_75t_L g2767 ( 
.A(n_2676),
.B(n_325),
.Y(n_2767)
);

NOR2xp33_ASAP7_75t_L g2768 ( 
.A(n_2720),
.B(n_326),
.Y(n_2768)
);

NAND2xp5_ASAP7_75t_L g2769 ( 
.A(n_2678),
.B(n_326),
.Y(n_2769)
);

NOR4xp25_ASAP7_75t_L g2770 ( 
.A(n_2705),
.B(n_327),
.C(n_328),
.D(n_329),
.Y(n_2770)
);

INVx4_ASAP7_75t_L g2771 ( 
.A(n_2692),
.Y(n_2771)
);

NAND4xp25_ASAP7_75t_L g2772 ( 
.A(n_2695),
.B(n_327),
.C(n_328),
.D(n_329),
.Y(n_2772)
);

AOI21xp5_ASAP7_75t_L g2773 ( 
.A1(n_2690),
.A2(n_330),
.B(n_331),
.Y(n_2773)
);

OAI22xp5_ASAP7_75t_L g2774 ( 
.A1(n_2682),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_2774)
);

NOR3xp33_ASAP7_75t_L g2775 ( 
.A(n_2729),
.B(n_332),
.C(n_333),
.Y(n_2775)
);

NOR4xp25_ASAP7_75t_L g2776 ( 
.A(n_2709),
.B(n_333),
.C(n_334),
.D(n_335),
.Y(n_2776)
);

NOR2xp33_ASAP7_75t_L g2777 ( 
.A(n_2684),
.B(n_335),
.Y(n_2777)
);

OR2x2_ASAP7_75t_L g2778 ( 
.A(n_2677),
.B(n_336),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2723),
.Y(n_2779)
);

NAND3xp33_ASAP7_75t_L g2780 ( 
.A(n_2683),
.B(n_337),
.C(n_338),
.Y(n_2780)
);

NOR3xp33_ASAP7_75t_L g2781 ( 
.A(n_2704),
.B(n_338),
.C(n_339),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2685),
.B(n_2716),
.Y(n_2782)
);

HB1xp67_ASAP7_75t_L g2783 ( 
.A(n_2700),
.Y(n_2783)
);

NOR2xp33_ASAP7_75t_L g2784 ( 
.A(n_2746),
.B(n_2693),
.Y(n_2784)
);

AOI221xp5_ASAP7_75t_SL g2785 ( 
.A1(n_2782),
.A2(n_2773),
.B1(n_2737),
.B2(n_2721),
.C(n_2772),
.Y(n_2785)
);

NAND4xp75_ASAP7_75t_L g2786 ( 
.A(n_2765),
.B(n_2687),
.C(n_2732),
.D(n_2722),
.Y(n_2786)
);

NAND3xp33_ASAP7_75t_SL g2787 ( 
.A(n_2770),
.B(n_2734),
.C(n_2713),
.Y(n_2787)
);

OAI21xp33_ASAP7_75t_SL g2788 ( 
.A1(n_2749),
.A2(n_2670),
.B(n_2689),
.Y(n_2788)
);

NOR2xp67_ASAP7_75t_L g2789 ( 
.A(n_2750),
.B(n_2730),
.Y(n_2789)
);

INVxp67_ASAP7_75t_SL g2790 ( 
.A(n_2754),
.Y(n_2790)
);

A2O1A1Ixp33_ASAP7_75t_SL g2791 ( 
.A1(n_2736),
.A2(n_2714),
.B(n_2686),
.C(n_2699),
.Y(n_2791)
);

AND2x4_ASAP7_75t_L g2792 ( 
.A(n_2757),
.B(n_339),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2757),
.Y(n_2793)
);

NAND5xp2_ASAP7_75t_L g2794 ( 
.A(n_2740),
.B(n_340),
.C(n_341),
.D(n_342),
.E(n_343),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2767),
.Y(n_2795)
);

NOR2x1p5_ASAP7_75t_L g2796 ( 
.A(n_2745),
.B(n_341),
.Y(n_2796)
);

AND3x4_ASAP7_75t_L g2797 ( 
.A(n_2760),
.B(n_344),
.C(n_345),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_L g2798 ( 
.A(n_2764),
.B(n_344),
.Y(n_2798)
);

NOR4xp75_ASAP7_75t_SL g2799 ( 
.A(n_2753),
.B(n_345),
.C(n_346),
.D(n_347),
.Y(n_2799)
);

AOI221xp5_ASAP7_75t_L g2800 ( 
.A1(n_2747),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.C(n_349),
.Y(n_2800)
);

NAND3xp33_ASAP7_75t_L g2801 ( 
.A(n_2751),
.B(n_348),
.C(n_350),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2743),
.A2(n_350),
.B1(n_351),
.B2(n_352),
.Y(n_2802)
);

OAI221xp5_ASAP7_75t_L g2803 ( 
.A1(n_2752),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.C(n_355),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2744),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_SL g2805 ( 
.A(n_2755),
.B(n_353),
.Y(n_2805)
);

NOR3xp33_ASAP7_75t_SL g2806 ( 
.A(n_2762),
.B(n_354),
.C(n_355),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2769),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2768),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2741),
.B(n_356),
.Y(n_2809)
);

NOR2x1_ASAP7_75t_L g2810 ( 
.A(n_2780),
.B(n_356),
.Y(n_2810)
);

AND2x2_ASAP7_75t_L g2811 ( 
.A(n_2776),
.B(n_357),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2778),
.Y(n_2812)
);

OR2x2_ASAP7_75t_L g2813 ( 
.A(n_2761),
.B(n_357),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2758),
.Y(n_2814)
);

OAI21xp33_ASAP7_75t_L g2815 ( 
.A1(n_2748),
.A2(n_358),
.B(n_359),
.Y(n_2815)
);

NOR2xp33_ASAP7_75t_R g2816 ( 
.A(n_2777),
.B(n_358),
.Y(n_2816)
);

AOI221xp5_ASAP7_75t_L g2817 ( 
.A1(n_2738),
.A2(n_359),
.B1(n_360),
.B2(n_361),
.C(n_363),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2756),
.B(n_360),
.Y(n_2818)
);

INVx2_ASAP7_75t_SL g2819 ( 
.A(n_2742),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2771),
.B(n_361),
.Y(n_2820)
);

NOR2x1p5_ASAP7_75t_L g2821 ( 
.A(n_2771),
.B(n_363),
.Y(n_2821)
);

NOR2x1_ASAP7_75t_L g2822 ( 
.A(n_2763),
.B(n_364),
.Y(n_2822)
);

OR2x2_ASAP7_75t_L g2823 ( 
.A(n_2783),
.B(n_364),
.Y(n_2823)
);

AND3x2_ASAP7_75t_L g2824 ( 
.A(n_2766),
.B(n_365),
.C(n_366),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2775),
.B(n_365),
.Y(n_2825)
);

OR2x2_ASAP7_75t_L g2826 ( 
.A(n_2779),
.B(n_366),
.Y(n_2826)
);

AND2x4_ASAP7_75t_L g2827 ( 
.A(n_2793),
.B(n_2781),
.Y(n_2827)
);

NAND4xp75_ASAP7_75t_L g2828 ( 
.A(n_2785),
.B(n_2822),
.C(n_2810),
.D(n_2789),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2792),
.B(n_2759),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2806),
.B(n_2739),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_2826),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_2821),
.Y(n_2832)
);

XOR2x2_ASAP7_75t_L g2833 ( 
.A(n_2797),
.B(n_2824),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2792),
.B(n_2774),
.Y(n_2834)
);

OR2x2_ASAP7_75t_L g2835 ( 
.A(n_2794),
.B(n_367),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2805),
.B(n_367),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2823),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2813),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2811),
.B(n_368),
.Y(n_2839)
);

NOR2x1_ASAP7_75t_L g2840 ( 
.A(n_2786),
.B(n_368),
.Y(n_2840)
);

NAND2x1p5_ASAP7_75t_L g2841 ( 
.A(n_2795),
.B(n_369),
.Y(n_2841)
);

NAND3xp33_ASAP7_75t_L g2842 ( 
.A(n_2800),
.B(n_2798),
.C(n_2801),
.Y(n_2842)
);

HB1xp67_ASAP7_75t_L g2843 ( 
.A(n_2816),
.Y(n_2843)
);

AND4x1_ASAP7_75t_L g2844 ( 
.A(n_2784),
.B(n_369),
.C(n_370),
.D(n_371),
.Y(n_2844)
);

AND2x4_ASAP7_75t_SL g2845 ( 
.A(n_2814),
.B(n_370),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2815),
.B(n_372),
.Y(n_2846)
);

NAND3x1_ASAP7_75t_L g2847 ( 
.A(n_2818),
.B(n_373),
.C(n_374),
.Y(n_2847)
);

INVxp67_ASAP7_75t_L g2848 ( 
.A(n_2820),
.Y(n_2848)
);

OR4x2_ASAP7_75t_L g2849 ( 
.A(n_2787),
.B(n_373),
.C(n_374),
.D(n_375),
.Y(n_2849)
);

NAND2xp5_ASAP7_75t_SL g2850 ( 
.A(n_2799),
.B(n_375),
.Y(n_2850)
);

OR3x1_ASAP7_75t_L g2851 ( 
.A(n_2809),
.B(n_376),
.C(n_377),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2790),
.B(n_377),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2796),
.B(n_378),
.Y(n_2853)
);

NAND3xp33_ASAP7_75t_SL g2854 ( 
.A(n_2825),
.B(n_378),
.C(n_379),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2804),
.Y(n_2855)
);

AND2x2_ASAP7_75t_L g2856 ( 
.A(n_2839),
.B(n_2819),
.Y(n_2856)
);

CKINVDCx20_ASAP7_75t_R g2857 ( 
.A(n_2833),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2841),
.B(n_2812),
.Y(n_2858)
);

NAND3xp33_ASAP7_75t_L g2859 ( 
.A(n_2852),
.B(n_2807),
.C(n_2808),
.Y(n_2859)
);

NAND2xp33_ASAP7_75t_R g2860 ( 
.A(n_2830),
.B(n_2803),
.Y(n_2860)
);

NAND2x1p5_ASAP7_75t_L g2861 ( 
.A(n_2840),
.B(n_2788),
.Y(n_2861)
);

AND2x4_ASAP7_75t_L g2862 ( 
.A(n_2850),
.B(n_2802),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2851),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2835),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2847),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2849),
.Y(n_2866)
);

O2A1O1Ixp33_ASAP7_75t_L g2867 ( 
.A1(n_2853),
.A2(n_2791),
.B(n_2817),
.C(n_381),
.Y(n_2867)
);

XNOR2x1_ASAP7_75t_L g2868 ( 
.A(n_2828),
.B(n_379),
.Y(n_2868)
);

NAND4xp75_ASAP7_75t_L g2869 ( 
.A(n_2855),
.B(n_380),
.C(n_382),
.D(n_383),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2836),
.Y(n_2870)
);

INVx1_ASAP7_75t_SL g2871 ( 
.A(n_2845),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2846),
.Y(n_2872)
);

AOI221xp5_ASAP7_75t_L g2873 ( 
.A1(n_2854),
.A2(n_2827),
.B1(n_2829),
.B2(n_2842),
.C(n_2848),
.Y(n_2873)
);

AOI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_2837),
.A2(n_382),
.B1(n_384),
.B2(n_385),
.Y(n_2874)
);

AOI211xp5_ASAP7_75t_SL g2875 ( 
.A1(n_2843),
.A2(n_385),
.B(n_386),
.C(n_387),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2834),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2832),
.B(n_386),
.Y(n_2877)
);

NOR2xp33_ASAP7_75t_L g2878 ( 
.A(n_2831),
.B(n_387),
.Y(n_2878)
);

NOR2x1_ASAP7_75t_L g2879 ( 
.A(n_2838),
.B(n_388),
.Y(n_2879)
);

CKINVDCx20_ASAP7_75t_R g2880 ( 
.A(n_2844),
.Y(n_2880)
);

INVx1_ASAP7_75t_L g2881 ( 
.A(n_2850),
.Y(n_2881)
);

OAI211xp5_ASAP7_75t_L g2882 ( 
.A1(n_2852),
.A2(n_389),
.B(n_390),
.C(n_391),
.Y(n_2882)
);

OAI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2852),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_2883)
);

AOI22xp5_ASAP7_75t_L g2884 ( 
.A1(n_2852),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_2884)
);

AOI22xp5_ASAP7_75t_L g2885 ( 
.A1(n_2852),
.A2(n_392),
.B1(n_393),
.B2(n_395),
.Y(n_2885)
);

OAI22xp5_ASAP7_75t_L g2886 ( 
.A1(n_2852),
.A2(n_395),
.B1(n_396),
.B2(n_397),
.Y(n_2886)
);

XOR2xp5_ASAP7_75t_L g2887 ( 
.A(n_2857),
.B(n_396),
.Y(n_2887)
);

XOR2xp5_ASAP7_75t_L g2888 ( 
.A(n_2868),
.B(n_398),
.Y(n_2888)
);

AO22x1_ASAP7_75t_L g2889 ( 
.A1(n_2879),
.A2(n_398),
.B1(n_399),
.B2(n_401),
.Y(n_2889)
);

OA22x2_ASAP7_75t_L g2890 ( 
.A1(n_2881),
.A2(n_399),
.B1(n_401),
.B2(n_403),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2866),
.Y(n_2891)
);

AO22x2_ASAP7_75t_L g2892 ( 
.A1(n_2871),
.A2(n_404),
.B1(n_405),
.B2(n_406),
.Y(n_2892)
);

XNOR2x1_ASAP7_75t_L g2893 ( 
.A(n_2876),
.B(n_404),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2861),
.Y(n_2894)
);

INVx3_ASAP7_75t_L g2895 ( 
.A(n_2862),
.Y(n_2895)
);

OA22x2_ASAP7_75t_L g2896 ( 
.A1(n_2882),
.A2(n_407),
.B1(n_408),
.B2(n_409),
.Y(n_2896)
);

INVx1_ASAP7_75t_SL g2897 ( 
.A(n_2880),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2869),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2862),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2858),
.Y(n_2900)
);

AOI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_2860),
.A2(n_409),
.B1(n_410),
.B2(n_411),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2863),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2856),
.Y(n_2903)
);

AO211x2_ASAP7_75t_L g2904 ( 
.A1(n_2891),
.A2(n_2859),
.B(n_2865),
.C(n_2864),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2896),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2888),
.B(n_2867),
.Y(n_2906)
);

HB1xp67_ASAP7_75t_L g2907 ( 
.A(n_2889),
.Y(n_2907)
);

INVx1_ASAP7_75t_SL g2908 ( 
.A(n_2887),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2903),
.A2(n_2870),
.B1(n_2872),
.B2(n_2873),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2893),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2890),
.Y(n_2911)
);

XNOR2xp5_ASAP7_75t_L g2912 ( 
.A(n_2897),
.B(n_2884),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2907),
.Y(n_2913)
);

INVx2_ASAP7_75t_L g2914 ( 
.A(n_2904),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2911),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2905),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2912),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2910),
.Y(n_2918)
);

XOR2xp5_ASAP7_75t_L g2919 ( 
.A(n_2917),
.B(n_2899),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2914),
.B(n_2895),
.Y(n_2920)
);

NAND2xp33_ASAP7_75t_SL g2921 ( 
.A(n_2913),
.B(n_2898),
.Y(n_2921)
);

OAI21xp5_ASAP7_75t_SL g2922 ( 
.A1(n_2915),
.A2(n_2909),
.B(n_2894),
.Y(n_2922)
);

NOR3xp33_ASAP7_75t_L g2923 ( 
.A(n_2922),
.B(n_2916),
.C(n_2900),
.Y(n_2923)
);

XNOR2x1_ASAP7_75t_L g2924 ( 
.A(n_2919),
.B(n_2902),
.Y(n_2924)
);

OAI21x1_ASAP7_75t_SL g2925 ( 
.A1(n_2920),
.A2(n_2918),
.B(n_2901),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_2921),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2926),
.Y(n_2927)
);

INVxp33_ASAP7_75t_SL g2928 ( 
.A(n_2923),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2924),
.Y(n_2929)
);

NOR2xp33_ASAP7_75t_L g2930 ( 
.A(n_2928),
.B(n_2908),
.Y(n_2930)
);

AOI22xp33_ASAP7_75t_L g2931 ( 
.A1(n_2930),
.A2(n_2927),
.B1(n_2929),
.B2(n_2925),
.Y(n_2931)
);

AOI21xp5_ASAP7_75t_L g2932 ( 
.A1(n_2931),
.A2(n_2906),
.B(n_2883),
.Y(n_2932)
);

AOI22xp5_ASAP7_75t_L g2933 ( 
.A1(n_2932),
.A2(n_2892),
.B1(n_2886),
.B2(n_2878),
.Y(n_2933)
);

OAI221xp5_ASAP7_75t_R g2934 ( 
.A1(n_2933),
.A2(n_2885),
.B1(n_2874),
.B2(n_2875),
.C(n_2877),
.Y(n_2934)
);

A2O1A1Ixp33_ASAP7_75t_L g2935 ( 
.A1(n_2934),
.A2(n_410),
.B(n_411),
.C(n_412),
.Y(n_2935)
);

AOI211xp5_ASAP7_75t_L g2936 ( 
.A1(n_2935),
.A2(n_413),
.B(n_414),
.C(n_415),
.Y(n_2936)
);


endmodule