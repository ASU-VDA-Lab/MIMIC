module fake_jpeg_28730_n_111 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_111);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_111;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_1),
.Y(n_50)
);

INVx3_ASAP7_75t_SL g51 ( 
.A(n_47),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_54),
.Y(n_60)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_2),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_63),
.Y(n_75)
);

CKINVDCx6p67_ASAP7_75t_R g57 ( 
.A(n_54),
.Y(n_57)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_38),
.B1(n_48),
.B2(n_41),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_58),
.A2(n_36),
.B1(n_35),
.B2(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_49),
.B(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g64 ( 
.A(n_55),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_49),
.B(n_45),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_45),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_60),
.A2(n_44),
.B(n_42),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_70),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_73),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_14),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_57),
.B(n_59),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_65),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_74),
.B(n_76),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_62),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_19),
.Y(n_78)
);

XNOR2x1_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_79),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_32),
.B(n_17),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_57),
.B(n_3),
.C(n_4),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_21),
.B(n_22),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_86),
.B(n_88),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_87),
.B(n_94),
.C(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_16),
.B(n_18),
.C(n_20),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_99),
.Y(n_104)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_100),
.A2(n_92),
.B(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_89),
.C(n_95),
.Y(n_103)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_104),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g107 ( 
.A1(n_105),
.A2(n_97),
.B(n_84),
.C(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_106),
.C(n_100),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_110),
.Y(n_111)
);


endmodule