module real_jpeg_17322_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_61;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_206;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

AND2x2_ASAP7_75t_L g32 ( 
.A(n_0),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_0),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_0),
.B(n_39),
.Y(n_82)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_0),
.B(n_91),
.Y(n_90)
);

AND2x4_ASAP7_75t_SL g127 ( 
.A(n_0),
.B(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_0),
.Y(n_145)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_2),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_3),
.B(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_4),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_4),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_5),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_5),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_5),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_5),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_5),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_5),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_5),
.B(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_6),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_8),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_9),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_9),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_9),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_9),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_9),
.B(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_10),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_12),
.Y(n_152)
);

BUFx4f_ASAP7_75t_L g227 ( 
.A(n_12),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_13),
.Y(n_102)
);

AOI22x1_ASAP7_75t_SL g110 ( 
.A1(n_13),
.A2(n_14),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_14),
.B(n_60),
.Y(n_59)
);

AOI31xp33_ASAP7_75t_L g100 ( 
.A1(n_14),
.A2(n_101),
.A3(n_104),
.B(n_110),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_14),
.B(n_174),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_14),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_14),
.B(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_160),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_158),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NOR2xp67_ASAP7_75t_SL g159 ( 
.A(n_18),
.B(n_96),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.C(n_83),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_19),
.A2(n_20),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_47),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_22),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_28),
.C(n_31),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_23),
.A2(n_31),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_23),
.Y(n_183)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

XOR2x1_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_32),
.Y(n_182)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_36),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_37),
.B(n_42),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_41),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_47),
.B(n_133),
.C(n_134),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_48),
.B(n_53),
.C(n_59),
.Y(n_157)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_51),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_53),
.A2(n_64),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_53),
.B(n_210),
.C(n_214),
.Y(n_234)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_65),
.A2(n_83),
.B1(n_84),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_74),
.C(n_78),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_66),
.B(n_74),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_67),
.B(n_70),
.Y(n_85)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_70),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_70),
.A2(n_205),
.B1(n_206),
.B2(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_78),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g197 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_82),
.Y(n_198)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_86)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_90),
.Y(n_95)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_131),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_117),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_127),
.B2(n_130),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_171),
.C(n_173),
.Y(n_170)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2x1_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

XNOR2x1_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_155),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_143),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_148),
.B1(n_153),
.B2(n_154),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_144),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_148),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_150),
.Y(n_193)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_184),
.B(n_237),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_163),
.B(n_167),
.Y(n_237)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_179),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_173),
.Y(n_188)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21x1_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_201),
.B(n_236),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_199),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_186),
.B(n_199),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_189),
.C(n_197),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_187),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_190),
.B1(n_197),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_191),
.B(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_197),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_224),
.Y(n_223)
);

AOI21x1_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_230),
.B(n_235),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_217),
.B(n_229),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_209),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_223),
.B(n_228),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_219),
.B(n_221),
.Y(n_228)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2x1_ASAP7_75t_SL g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);


endmodule