module real_aes_2753_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_791;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_505;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g556 ( .A(n_0), .B(n_179), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_1), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g140 ( .A(n_2), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_3), .B(n_479), .Y(n_511) );
NAND2xp33_ASAP7_75t_SL g505 ( .A(n_4), .B(n_161), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_5), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_6), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g498 ( .A(n_7), .Y(n_498) );
INVx1_ASAP7_75t_L g238 ( .A(n_8), .Y(n_238) );
CKINVDCx16_ASAP7_75t_R g804 ( .A(n_9), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_10), .Y(n_230) );
AND2x2_ASAP7_75t_L g509 ( .A(n_11), .B(n_130), .Y(n_509) );
INVx2_ASAP7_75t_L g131 ( .A(n_12), .Y(n_131) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_13), .Y(n_113) );
NOR3xp33_ASAP7_75t_L g802 ( .A(n_13), .B(n_803), .C(n_805), .Y(n_802) );
INVx1_ASAP7_75t_L g180 ( .A(n_14), .Y(n_180) );
AOI221x1_ASAP7_75t_L g501 ( .A1(n_15), .A2(n_163), .B1(n_478), .B2(n_502), .C(n_504), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_16), .B(n_479), .Y(n_487) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
INVx1_ASAP7_75t_L g177 ( .A(n_18), .Y(n_177) );
INVx1_ASAP7_75t_SL g152 ( .A(n_19), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_20), .B(n_155), .Y(n_194) );
AOI33xp33_ASAP7_75t_L g247 ( .A1(n_21), .A2(n_52), .A3(n_137), .B1(n_148), .B2(n_248), .B3(n_249), .Y(n_247) );
AOI221xp5_ASAP7_75t_SL g477 ( .A1(n_22), .A2(n_40), .B1(n_478), .B2(n_479), .C(n_480), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_23), .A2(n_478), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_24), .B(n_179), .Y(n_514) );
INVx1_ASAP7_75t_L g223 ( .A(n_25), .Y(n_223) );
OR2x2_ASAP7_75t_L g132 ( .A(n_26), .B(n_92), .Y(n_132) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_26), .A2(n_92), .B(n_131), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_27), .B(n_182), .Y(n_491) );
INVxp67_ASAP7_75t_L g500 ( .A(n_28), .Y(n_500) );
AND2x2_ASAP7_75t_L g545 ( .A(n_29), .B(n_129), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_30), .B(n_135), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_31), .A2(n_478), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_32), .B(n_182), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g759 ( .A1(n_33), .A2(n_43), .B1(n_760), .B2(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_33), .Y(n_760) );
AND2x2_ASAP7_75t_L g142 ( .A(n_34), .B(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g147 ( .A(n_34), .Y(n_147) );
AND2x2_ASAP7_75t_L g161 ( .A(n_34), .B(n_140), .Y(n_161) );
OR2x6_ASAP7_75t_L g114 ( .A(n_35), .B(n_115), .Y(n_114) );
INVxp67_ASAP7_75t_L g805 ( .A(n_35), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_36), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_37), .B(n_135), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_38), .A2(n_164), .B1(n_170), .B2(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_39), .B(n_196), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_41), .A2(n_83), .B1(n_145), .B2(n_478), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_42), .B(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g761 ( .A(n_43), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_44), .B(n_179), .Y(n_543) );
OAI22xp5_ASAP7_75t_SL g782 ( .A1(n_45), .A2(n_79), .B1(n_783), .B2(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_45), .Y(n_784) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_46), .B(n_198), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_47), .B(n_155), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_48), .Y(n_191) );
AND2x2_ASAP7_75t_L g559 ( .A(n_49), .B(n_129), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_50), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_51), .B(n_129), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_53), .B(n_155), .Y(n_269) );
INVx1_ASAP7_75t_L g138 ( .A(n_54), .Y(n_138) );
INVx1_ASAP7_75t_L g157 ( .A(n_54), .Y(n_157) );
AND2x2_ASAP7_75t_L g270 ( .A(n_55), .B(n_129), .Y(n_270) );
AOI221xp5_ASAP7_75t_L g236 ( .A1(n_56), .A2(n_74), .B1(n_135), .B2(n_145), .C(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_57), .B(n_135), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g544 ( .A(n_58), .B(n_479), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_59), .B(n_164), .Y(n_232) );
AOI21xp5_ASAP7_75t_SL g203 ( .A1(n_60), .A2(n_145), .B(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g524 ( .A(n_61), .B(n_129), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_62), .B(n_182), .Y(n_557) );
INVx1_ASAP7_75t_L g173 ( .A(n_63), .Y(n_173) );
AND2x2_ASAP7_75t_SL g492 ( .A(n_64), .B(n_130), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_65), .B(n_179), .Y(n_522) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_66), .A2(n_478), .B(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g268 ( .A(n_67), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_68), .B(n_182), .Y(n_515) );
AND2x2_ASAP7_75t_SL g530 ( .A(n_69), .B(n_198), .Y(n_530) );
OAI22xp5_ASAP7_75t_SL g790 ( .A1(n_70), .A2(n_91), .B1(n_791), .B2(n_792), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_70), .Y(n_791) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_71), .A2(n_145), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g143 ( .A(n_72), .Y(n_143) );
INVx1_ASAP7_75t_L g159 ( .A(n_72), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_73), .B(n_135), .Y(n_250) );
AND2x2_ASAP7_75t_L g162 ( .A(n_75), .B(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g174 ( .A(n_76), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_77), .A2(n_145), .B(n_151), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_78), .Y(n_808) );
INVx1_ASAP7_75t_L g783 ( .A(n_79), .Y(n_783) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_80), .A2(n_145), .B(n_193), .C(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_81), .B(n_479), .Y(n_523) );
AOI22xp5_ASAP7_75t_L g528 ( .A1(n_82), .A2(n_86), .B1(n_135), .B2(n_479), .Y(n_528) );
INVx1_ASAP7_75t_L g117 ( .A(n_84), .Y(n_117) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_85), .B(n_163), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_87), .A2(n_145), .B1(n_245), .B2(n_246), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_88), .B(n_179), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_89), .B(n_179), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_90), .A2(n_478), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_91), .B(n_412), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g464 ( .A1(n_91), .A2(n_465), .B(n_466), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g467 ( .A1(n_91), .A2(n_412), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g792 ( .A(n_91), .Y(n_792) );
INVx1_ASAP7_75t_L g205 ( .A(n_93), .Y(n_205) );
XNOR2xp5_ASAP7_75t_L g758 ( .A(n_94), .B(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_95), .B(n_182), .Y(n_521) );
AND2x2_ASAP7_75t_L g251 ( .A(n_96), .B(n_163), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_97), .A2(n_221), .B(n_222), .C(n_224), .Y(n_220) );
INVxp67_ASAP7_75t_L g503 ( .A(n_98), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_99), .B(n_479), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_100), .B(n_182), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_101), .A2(n_478), .B(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g772 ( .A(n_102), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_103), .B(n_155), .Y(n_206) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_798), .B(n_807), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_769), .B1(n_777), .B2(n_794), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_758), .B(n_762), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OAI21x1_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_118), .B(n_469), .Y(n_108) );
OAI22xp5_ASAP7_75t_SL g763 ( .A1(n_109), .A2(n_119), .B1(n_470), .B2(n_764), .Y(n_763) );
CKINVDCx6p67_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
INVx3_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
AND2x6_ASAP7_75t_SL g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OR2x6_ASAP7_75t_SL g756 ( .A(n_113), .B(n_757), .Y(n_756) );
OR2x2_ASAP7_75t_L g768 ( .A(n_113), .B(n_114), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_113), .B(n_757), .Y(n_776) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_114), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_116), .B(n_117), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_116), .B(n_117), .Y(n_806) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_464), .C(n_467), .Y(n_119) );
NAND4xp25_ASAP7_75t_L g120 ( .A(n_121), .B(n_351), .C(n_411), .D(n_439), .Y(n_120) );
INVx1_ASAP7_75t_L g468 ( .A(n_121), .Y(n_468) );
NAND3x1_ASAP7_75t_L g786 ( .A(n_121), .B(n_351), .C(n_787), .Y(n_786) );
AND3x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_290), .C(n_318), .Y(n_121) );
AOI221x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_213), .B1(n_252), .B2(n_256), .C(n_276), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AOI21xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_184), .B(n_208), .Y(n_124) );
AND2x4_ASAP7_75t_L g360 ( .A(n_125), .B(n_210), .Y(n_360) );
AND2x4_ASAP7_75t_SL g125 ( .A(n_126), .B(n_166), .Y(n_125) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_126), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_126), .B(n_342), .Y(n_459) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g209 ( .A(n_127), .B(n_168), .Y(n_209) );
INVx2_ASAP7_75t_L g283 ( .A(n_127), .Y(n_283) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_127), .Y(n_343) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_127), .Y(n_350) );
AND2x2_ASAP7_75t_L g355 ( .A(n_127), .B(n_167), .Y(n_355) );
INVx1_ASAP7_75t_L g385 ( .A(n_127), .Y(n_385) );
OR2x2_ASAP7_75t_L g438 ( .A(n_127), .B(n_200), .Y(n_438) );
AO21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_133), .B(n_162), .Y(n_127) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_128), .A2(n_518), .B(n_524), .Y(n_517) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_128), .A2(n_539), .B(n_545), .Y(n_538) );
AO21x2_ASAP7_75t_L g602 ( .A1(n_128), .A2(n_539), .B(n_545), .Y(n_602) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_129), .A2(n_477), .B(n_483), .Y(n_476) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_SL g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x4_ASAP7_75t_L g170 ( .A(n_131), .B(n_132), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_134), .B(n_144), .Y(n_133) );
INVx1_ASAP7_75t_L g233 ( .A(n_135), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_135), .A2(n_145), .B1(n_497), .B2(n_499), .Y(n_496) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_141), .Y(n_135) );
INVx1_ASAP7_75t_L g189 ( .A(n_136), .Y(n_189) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
OR2x6_ASAP7_75t_L g153 ( .A(n_137), .B(n_149), .Y(n_153) );
INVxp33_ASAP7_75t_L g248 ( .A(n_137), .Y(n_248) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g150 ( .A(n_138), .B(n_140), .Y(n_150) );
AND2x4_ASAP7_75t_L g182 ( .A(n_138), .B(n_158), .Y(n_182) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g190 ( .A(n_141), .Y(n_190) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g478 ( .A(n_142), .B(n_150), .Y(n_478) );
INVx2_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
AND2x6_ASAP7_75t_L g179 ( .A(n_143), .B(n_156), .Y(n_179) );
INVxp67_ASAP7_75t_L g231 ( .A(n_145), .Y(n_231) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NOR2x1p5_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx1_ASAP7_75t_L g249 ( .A(n_148), .Y(n_249) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_SL g151 ( .A1(n_152), .A2(n_153), .B(n_154), .C(n_160), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_173), .B1(n_174), .B2(n_175), .Y(n_172) );
INVx2_ASAP7_75t_L g196 ( .A(n_153), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g204 ( .A1(n_153), .A2(n_160), .B(n_205), .C(n_206), .Y(n_204) );
INVxp67_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
O2A1O1Ixp33_ASAP7_75t_SL g237 ( .A1(n_153), .A2(n_160), .B(n_238), .C(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g267 ( .A1(n_153), .A2(n_160), .B(n_268), .C(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g175 ( .A(n_155), .Y(n_175) );
AND2x4_ASAP7_75t_L g479 ( .A(n_155), .B(n_161), .Y(n_479) );
AND2x4_ASAP7_75t_L g155 ( .A(n_156), .B(n_158), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_160), .B(n_170), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_160), .A2(n_194), .B(n_195), .Y(n_193) );
INVx1_ASAP7_75t_L g245 ( .A(n_160), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_160), .A2(n_481), .B(n_482), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_160), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_160), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_160), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_160), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g555 ( .A1(n_160), .A2(n_556), .B(n_557), .Y(n_555) );
INVx5_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_161), .Y(n_224) );
OAI22xp5_ASAP7_75t_L g219 ( .A1(n_163), .A2(n_220), .B1(n_225), .B2(n_226), .Y(n_219) );
INVx3_ASAP7_75t_L g226 ( .A(n_163), .Y(n_226) );
INVx4_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_164), .B(n_229), .Y(n_228) );
AOI21x1_ASAP7_75t_L g552 ( .A1(n_164), .A2(n_553), .B(n_559), .Y(n_552) );
INVx3_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx4f_ASAP7_75t_L g198 ( .A(n_165), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_166), .B(n_200), .Y(n_365) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g255 ( .A(n_167), .B(n_186), .Y(n_255) );
AND2x2_ASAP7_75t_L g342 ( .A(n_167), .B(n_212), .Y(n_342) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g313 ( .A(n_168), .Y(n_313) );
NOR2x1_ASAP7_75t_SL g374 ( .A(n_168), .B(n_200), .Y(n_374) );
AND2x2_ASAP7_75t_L g395 ( .A(n_168), .B(n_186), .Y(n_395) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_171), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_170), .A2(n_203), .B(n_207), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_170), .B(n_498), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_170), .B(n_500), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_170), .B(n_503), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_170), .B(n_175), .C(n_505), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_170), .A2(n_511), .B(n_512), .Y(n_510) );
OAI21xp5_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_176), .B(n_183), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_175), .B(n_223), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B1(n_180), .B2(n_181), .Y(n_176) );
INVxp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVxp67_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g391 ( .A(n_184), .B(n_281), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_184), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_SL g184 ( .A(n_185), .B(n_199), .Y(n_184) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g212 ( .A(n_186), .Y(n_212) );
INVx1_ASAP7_75t_L g280 ( .A(n_186), .Y(n_280) );
AND2x2_ASAP7_75t_L g338 ( .A(n_186), .B(n_200), .Y(n_338) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_192), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .C(n_191), .Y(n_188) );
AO21x2_ASAP7_75t_L g242 ( .A1(n_197), .A2(n_243), .B(n_251), .Y(n_242) );
AO21x2_ASAP7_75t_L g289 ( .A1(n_197), .A2(n_243), .B(n_251), .Y(n_289) );
AOI21x1_ASAP7_75t_L g526 ( .A1(n_197), .A2(n_527), .B(n_530), .Y(n_526) );
INVx2_ASAP7_75t_SL g197 ( .A(n_198), .Y(n_197) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_198), .A2(n_236), .B(n_240), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_198), .A2(n_487), .B(n_488), .Y(n_486) );
NOR2x1_ASAP7_75t_L g253 ( .A(n_199), .B(n_254), .Y(n_253) );
AND2x4_ASAP7_75t_L g279 ( .A(n_199), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g317 ( .A(n_199), .B(n_209), .Y(n_317) );
INVx4_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g298 ( .A(n_200), .Y(n_298) );
AND2x4_ASAP7_75t_L g327 ( .A(n_200), .B(n_280), .Y(n_327) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_200), .Y(n_363) );
AND2x2_ASAP7_75t_L g462 ( .A(n_200), .B(n_313), .Y(n_462) );
OR2x6_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
OAI21xp33_ASAP7_75t_SL g460 ( .A1(n_208), .A2(n_461), .B(n_463), .Y(n_460) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_210), .Y(n_208) );
NOR2xp33_ASAP7_75t_SL g335 ( .A(n_209), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_SL g417 ( .A(n_210), .Y(n_417) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g381 ( .A1(n_215), .A2(n_285), .B1(n_326), .B2(n_342), .Y(n_381) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_234), .Y(n_215) );
INVx1_ASAP7_75t_L g436 ( .A(n_216), .Y(n_436) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g378 ( .A(n_217), .B(n_371), .Y(n_378) );
AND2x2_ASAP7_75t_L g416 ( .A(n_217), .B(n_234), .Y(n_416) );
INVx1_ASAP7_75t_L g430 ( .A(n_217), .Y(n_430) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g260 ( .A(n_218), .Y(n_260) );
AND2x4_ASAP7_75t_L g294 ( .A(n_218), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g303 ( .A(n_218), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_218), .B(n_263), .Y(n_333) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_227), .Y(n_218) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_226), .A2(n_264), .B(n_270), .Y(n_263) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_226), .A2(n_264), .B(n_270), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_231), .B1(n_232), .B2(n_233), .Y(n_227) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g274 ( .A(n_234), .B(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g314 ( .A(n_234), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g357 ( .A(n_234), .B(n_358), .Y(n_357) );
AND2x4_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
INVx1_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
INVx2_ASAP7_75t_L g295 ( .A(n_235), .Y(n_295) );
INVx1_ASAP7_75t_L g310 ( .A(n_235), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_235), .B(n_289), .Y(n_334) );
INVxp67_ASAP7_75t_L g390 ( .A(n_235), .Y(n_390) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g259 ( .A(n_242), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
AND2x4_ASAP7_75t_L g409 ( .A(n_242), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_244), .B(n_250), .Y(n_243) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
BUFx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_254), .A2(n_448), .B(n_449), .Y(n_447) );
INVx4_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g297 ( .A(n_255), .B(n_298), .Y(n_297) );
NAND2xp33_ASAP7_75t_SL g256 ( .A(n_257), .B(n_273), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g463 ( .A(n_259), .B(n_308), .Y(n_463) );
AND2x2_ASAP7_75t_L g286 ( .A(n_260), .B(n_272), .Y(n_286) );
AND2x2_ASAP7_75t_L g331 ( .A(n_260), .B(n_309), .Y(n_331) );
NOR2xp67_ASAP7_75t_L g358 ( .A(n_260), .B(n_309), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_262), .B(n_271), .Y(n_261) );
INVx3_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
AND2x4_ASAP7_75t_L g287 ( .A(n_262), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_262), .B(n_303), .Y(n_323) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_263), .B(n_289), .Y(n_305) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_263), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_271), .B(n_322), .Y(n_321) );
INVx3_ASAP7_75t_L g367 ( .A(n_271), .Y(n_367) );
BUFx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_275), .B(n_286), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_275), .B(n_343), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_284), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_278), .A2(n_428), .B(n_429), .Y(n_427) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
AND2x2_ASAP7_75t_L g311 ( .A(n_279), .B(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
AND2x2_ASAP7_75t_L g433 ( .A(n_279), .B(n_434), .Y(n_433) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_281), .B(n_321), .C(n_323), .Y(n_320) );
INVx1_ASAP7_75t_L g445 ( .A(n_281), .Y(n_445) );
INVx1_ASAP7_75t_L g455 ( .A(n_281), .Y(n_455) );
AND2x2_ASAP7_75t_L g461 ( .A(n_281), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_282), .Y(n_434) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_285), .B(n_363), .Y(n_441) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g345 ( .A(n_286), .Y(n_345) );
INVx1_ASAP7_75t_L g344 ( .A(n_287), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_287), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g322 ( .A(n_288), .Y(n_322) );
AND2x2_ASAP7_75t_L g371 ( .A(n_288), .B(n_309), .Y(n_371) );
AND2x2_ASAP7_75t_L g389 ( .A(n_288), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI222xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_297), .B1(n_299), .B2(n_311), .C1(n_314), .C2(n_317), .Y(n_290) );
NAND2xp33_ASAP7_75t_SL g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVx2_ASAP7_75t_SL g379 ( .A(n_292), .Y(n_379) );
NAND2x1_ASAP7_75t_SL g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g362 ( .A(n_293), .B(n_345), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_293), .B(n_307), .Y(n_448) );
INVx3_ASAP7_75t_L g398 ( .A(n_294), .Y(n_398) );
AND2x2_ASAP7_75t_L g408 ( .A(n_294), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_297), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g387 ( .A(n_298), .Y(n_387) );
NAND2xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_306), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OAI21xp33_ASAP7_75t_SL g442 ( .A1(n_301), .A2(n_443), .B(n_446), .Y(n_442) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g401 ( .A(n_302), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g307 ( .A(n_303), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2x1_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
INVx2_ASAP7_75t_L g410 ( .A(n_309), .Y(n_410) );
AND2x2_ASAP7_75t_L g326 ( .A(n_312), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NOR2x1_ASAP7_75t_L g386 ( .A(n_313), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_324), .C(n_339), .Y(n_318) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_322), .B(n_331), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B1(n_332), .B2(n_335), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g428 ( .A(n_327), .B(n_420), .Y(n_428) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_329), .A2(n_384), .B1(n_388), .B2(n_391), .Y(n_383) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g366 ( .A(n_330), .B(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g388 ( .A(n_331), .B(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_SL g400 ( .A(n_333), .Y(n_400) );
INVx2_ASAP7_75t_L g431 ( .A(n_334), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
AND2x2_ASAP7_75t_L g347 ( .A(n_338), .B(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_338), .A2(n_373), .B1(n_397), .B2(n_401), .Y(n_396) );
AND2x2_ASAP7_75t_L g422 ( .A(n_338), .B(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_344), .B1(n_345), .B2(n_346), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AND2x2_ASAP7_75t_SL g380 ( .A(n_342), .B(n_363), .Y(n_380) );
INVx2_ASAP7_75t_L g406 ( .A(n_342), .Y(n_406) );
BUFx2_ASAP7_75t_L g420 ( .A(n_343), .Y(n_420) );
NOR2xp33_ASAP7_75t_SL g435 ( .A(n_344), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g373 ( .A(n_348), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g465 ( .A(n_351), .Y(n_465) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_375), .Y(n_351) );
AOI21xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_363), .B(n_364), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_359), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_355), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_355), .A2(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_357), .A2(n_433), .B1(n_435), .B2(n_437), .Y(n_432) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_360), .A2(n_378), .B1(n_379), .B2(n_380), .Y(n_377) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g393 ( .A(n_363), .B(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g405 ( .A(n_363), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g407 ( .A(n_363), .B(n_395), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_368), .B2(n_372), .Y(n_364) );
NOR2xp67_ASAP7_75t_SL g369 ( .A(n_367), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g452 ( .A(n_367), .Y(n_452) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g424 ( .A(n_374), .Y(n_424) );
NOR2xp67_ASAP7_75t_L g375 ( .A(n_376), .B(n_382), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_381), .Y(n_376) );
NAND4xp25_ASAP7_75t_L g382 ( .A(n_383), .B(n_392), .C(n_396), .D(n_403), .Y(n_382) );
AND2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AND2x2_ASAP7_75t_L g394 ( .A(n_385), .B(n_395), .Y(n_394) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_389), .B(n_400), .Y(n_425) );
NAND2xp33_ASAP7_75t_SL g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g415 ( .A(n_402), .Y(n_415) );
OAI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_407), .B(n_408), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g454 ( .A(n_409), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g787 ( .A(n_413), .B(n_788), .Y(n_787) );
AOI211x1_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_417), .B(n_418), .C(n_426), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_417), .B(n_445), .Y(n_446) );
AOI31xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .A3(n_424), .B(n_425), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .Y(n_426) );
AND2x2_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_431), .B(n_457), .Y(n_456) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_434), .Y(n_450) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g466 ( .A(n_439), .Y(n_466) );
AOI21xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_447), .B(n_451), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g788 ( .A1(n_440), .A2(n_447), .B(n_451), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVxp33_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_456), .C(n_460), .Y(n_451) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NAND2x1_ASAP7_75t_SL g469 ( .A(n_470), .B(n_752), .Y(n_469) );
INVx4_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
OR2x6_ASAP7_75t_L g471 ( .A(n_472), .B(n_665), .Y(n_471) );
NAND3xp33_ASAP7_75t_SL g472 ( .A(n_473), .B(n_575), .C(n_615), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_493), .B(n_506), .C(n_531), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_474), .B(n_580), .Y(n_614) );
NOR2x1p5_ASAP7_75t_L g474 ( .A(n_475), .B(n_484), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g550 ( .A(n_476), .Y(n_550) );
INVx2_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
OR2x2_ASAP7_75t_L g578 ( .A(n_476), .B(n_485), .Y(n_578) );
AND2x2_ASAP7_75t_L g592 ( .A(n_476), .B(n_551), .Y(n_592) );
INVx1_ASAP7_75t_L g620 ( .A(n_476), .Y(n_620) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_476), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_476), .B(n_485), .Y(n_726) );
OR2x2_ASAP7_75t_L g547 ( .A(n_484), .B(n_548), .Y(n_547) );
HB1xp67_ASAP7_75t_L g682 ( .A(n_484), .Y(n_682) );
AND2x2_ASAP7_75t_L g687 ( .A(n_484), .B(n_549), .Y(n_687) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AND2x4_ASAP7_75t_L g493 ( .A(n_485), .B(n_494), .Y(n_493) );
OR2x2_ASAP7_75t_L g546 ( .A(n_485), .B(n_495), .Y(n_546) );
OR2x2_ASAP7_75t_L g565 ( .A(n_485), .B(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g594 ( .A(n_485), .Y(n_594) );
AND2x4_ASAP7_75t_SL g633 ( .A(n_485), .B(n_495), .Y(n_633) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_485), .Y(n_637) );
OR2x2_ASAP7_75t_L g654 ( .A(n_485), .B(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g664 ( .A(n_485), .B(n_571), .Y(n_664) );
INVx1_ASAP7_75t_L g693 ( .A(n_485), .Y(n_693) );
OR2x6_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_493), .B(n_622), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_494), .B(n_551), .Y(n_568) );
AND2x2_ASAP7_75t_L g580 ( .A(n_494), .B(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g598 ( .A(n_494), .B(n_565), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_494), .B(n_619), .Y(n_618) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_L g571 ( .A(n_495), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g593 ( .A(n_495), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g628 ( .A(n_495), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_495), .B(n_551), .Y(n_652) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_501), .Y(n_495) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_516), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_507), .B(n_584), .Y(n_583) );
AND2x4_ASAP7_75t_L g601 ( .A(n_507), .B(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_507), .B(n_517), .Y(n_606) );
NAND3xp33_ASAP7_75t_L g621 ( .A(n_507), .B(n_622), .C(n_623), .Y(n_621) );
AND2x2_ASAP7_75t_L g669 ( .A(n_507), .B(n_574), .Y(n_669) );
INVx5_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g536 ( .A(n_508), .B(n_537), .Y(n_536) );
AND2x4_ASAP7_75t_SL g573 ( .A(n_508), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g589 ( .A(n_508), .Y(n_589) );
OR2x2_ASAP7_75t_L g612 ( .A(n_508), .B(n_602), .Y(n_612) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_508), .Y(n_629) );
AND2x2_ASAP7_75t_SL g647 ( .A(n_508), .B(n_535), .Y(n_647) );
AND2x4_ASAP7_75t_L g662 ( .A(n_508), .B(n_538), .Y(n_662) );
AND2x2_ASAP7_75t_L g676 ( .A(n_508), .B(n_517), .Y(n_676) );
OR2x2_ASAP7_75t_L g697 ( .A(n_508), .B(n_525), .Y(n_697) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
AND2x2_ASAP7_75t_L g751 ( .A(n_516), .B(n_629), .Y(n_751) );
AND2x2_ASAP7_75t_L g516 ( .A(n_517), .B(n_525), .Y(n_516) );
AND2x4_ASAP7_75t_L g574 ( .A(n_517), .B(n_537), .Y(n_574) );
INVx2_ASAP7_75t_L g585 ( .A(n_517), .Y(n_585) );
AND2x2_ASAP7_75t_L g590 ( .A(n_517), .B(n_535), .Y(n_590) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_517), .Y(n_623) );
OR2x2_ASAP7_75t_L g646 ( .A(n_517), .B(n_538), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_517), .B(n_538), .Y(n_649) );
INVx1_ASAP7_75t_L g658 ( .A(n_517), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AND2x2_ASAP7_75t_L g561 ( .A(n_525), .B(n_538), .Y(n_561) );
BUFx2_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
AND2x2_ASAP7_75t_L g705 ( .A(n_525), .B(n_585), .Y(n_705) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_526), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_546), .B1(n_547), .B2(n_560), .C(n_562), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_534), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_534), .B(n_601), .Y(n_641) );
OR2x2_ASAP7_75t_L g653 ( .A(n_534), .B(n_649), .Y(n_653) );
OR2x2_ASAP7_75t_L g656 ( .A(n_534), .B(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g745 ( .A(n_534), .B(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g584 ( .A(n_535), .B(n_585), .Y(n_584) );
OA33x2_ASAP7_75t_L g617 ( .A1(n_535), .A2(n_578), .A3(n_618), .B1(n_621), .B2(n_624), .B3(n_627), .Y(n_617) );
OR2x2_ASAP7_75t_L g648 ( .A(n_535), .B(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g672 ( .A(n_535), .B(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g680 ( .A(n_535), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g700 ( .A(n_535), .B(n_574), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_535), .B(n_589), .Y(n_738) );
INVx2_ASAP7_75t_L g608 ( .A(n_536), .Y(n_608) );
AOI322xp5_ASAP7_75t_L g678 ( .A1(n_536), .A2(n_591), .A3(n_679), .B1(n_682), .B2(n_683), .C1(n_685), .C2(n_687), .Y(n_678) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_538), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
OR2x2_ASAP7_75t_L g660 ( .A(n_546), .B(n_639), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g712 ( .A(n_546), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g733 ( .A(n_546), .Y(n_733) );
INVx1_ASAP7_75t_SL g599 ( .A(n_547), .Y(n_599) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g632 ( .A(n_549), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_L g572 ( .A(n_551), .Y(n_572) );
INVx1_ASAP7_75t_L g581 ( .A(n_551), .Y(n_581) );
INVx1_ASAP7_75t_L g622 ( .A(n_551), .Y(n_622) );
OR2x2_ASAP7_75t_L g639 ( .A(n_551), .B(n_566), .Y(n_639) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_551), .Y(n_714) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_558), .Y(n_553) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_SL g683 ( .A(n_561), .B(n_684), .Y(n_683) );
OAI21xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_569), .B(n_573), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_563), .A2(n_637), .B(n_638), .C(n_640), .Y(n_636) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g701 ( .A(n_565), .B(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_566), .Y(n_570) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g725 ( .A(n_568), .B(n_726), .Y(n_725) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
AND2x2_ASAP7_75t_SL g694 ( .A(n_571), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g702 ( .A(n_571), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_571), .B(n_693), .Y(n_710) );
INVx3_ASAP7_75t_SL g635 ( .A(n_574), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_576), .A2(n_582), .B1(n_586), .B2(n_591), .C(n_595), .Y(n_575) );
INVx1_ASAP7_75t_SL g576 ( .A(n_577), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
INVx1_ASAP7_75t_SL g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_581), .Y(n_626) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_584), .A2(n_611), .B(n_683), .Y(n_689) );
AND2x2_ASAP7_75t_L g715 ( .A(n_584), .B(n_662), .Y(n_715) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_585), .Y(n_603) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_589), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g724 ( .A(n_589), .B(n_646), .Y(n_724) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
INVx2_ASAP7_75t_L g673 ( .A(n_592), .Y(n_673) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_600), .B(n_604), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx2_ASAP7_75t_L g746 ( .A(n_601), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_602), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g675 ( .A(n_602), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_603), .B(n_625), .Y(n_624) );
OAI31xp33_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .A3(n_609), .B(n_613), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_608), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
OR2x2_ASAP7_75t_L g686 ( .A(n_610), .B(n_612), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_610), .B(n_662), .Y(n_741) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR5xp2_ASAP7_75t_L g615 ( .A(n_616), .B(n_630), .C(n_642), .D(n_651), .E(n_659), .Y(n_615) );
INVxp67_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_620), .B(n_622), .Y(n_655) );
INVx1_ASAP7_75t_L g695 ( .A(n_620), .Y(n_695) );
INVxp67_ASAP7_75t_SL g732 ( .A(n_620), .Y(n_732) );
INVx1_ASAP7_75t_L g684 ( .A(n_623), .Y(n_684) );
INVxp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp33_ASAP7_75t_SL g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OAI321xp33_ASAP7_75t_L g667 ( .A1(n_628), .A2(n_668), .A3(n_670), .B1(n_674), .B2(n_677), .C(n_678), .Y(n_667) );
INVx1_ASAP7_75t_L g721 ( .A(n_629), .Y(n_721) );
OAI21xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_636), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_632), .A2(n_705), .B1(n_712), .B2(n_715), .Y(n_711) );
AND2x2_ASAP7_75t_L g740 ( .A(n_633), .B(n_714), .Y(n_740) );
INVx1_ASAP7_75t_L g650 ( .A(n_638), .Y(n_650) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_648), .B(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_649), .A2(n_660), .B1(n_661), .B2(n_663), .Y(n_659) );
INVx1_ASAP7_75t_L g722 ( .A(n_649), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_654), .B2(n_656), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_658), .B(n_662), .Y(n_661) );
OAI221xp5_ASAP7_75t_L g736 ( .A1(n_660), .A2(n_737), .B1(n_739), .B2(n_741), .C(n_742), .Y(n_736) );
INVx1_ASAP7_75t_L g743 ( .A(n_660), .Y(n_743) );
OAI221xp5_ASAP7_75t_L g717 ( .A1(n_661), .A2(n_718), .B1(n_725), .B2(n_727), .C(n_728), .Y(n_717) );
OAI21xp5_ASAP7_75t_L g688 ( .A1(n_663), .A2(n_689), .B(n_690), .Y(n_688) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_716), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_688), .C(n_706), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_669), .Y(n_735) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g734 ( .A(n_677), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_679), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g727 ( .A(n_687), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_696), .B(n_698), .Y(n_690) );
INVxp67_ASAP7_75t_L g748 ( .A(n_691), .Y(n_748) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g703 ( .A(n_694), .Y(n_703) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_703), .B2(n_704), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B(n_711), .Y(n_706) );
INVx1_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g749 ( .A(n_712), .Y(n_749) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_736), .C(n_747), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_734), .B(n_735), .Y(n_728) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g742 ( .A1(n_740), .A2(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
AOI21xp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_750), .Y(n_747) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
BUFx4f_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g764 ( .A(n_755), .Y(n_764) );
CKINVDCx11_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
AOI21xp33_ASAP7_75t_SL g762 ( .A1(n_758), .A2(n_763), .B(n_765), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
BUFx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_770), .B(n_773), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_772), .Y(n_771) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_772), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g777 ( .A1(n_773), .A2(n_778), .B(n_780), .Y(n_777) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
BUFx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx2_ASAP7_75t_R g779 ( .A(n_776), .Y(n_779) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
OAI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_782), .B1(n_785), .B2(n_793), .Y(n_780) );
CKINVDCx20_ASAP7_75t_R g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g793 ( .A(n_785), .Y(n_793) );
XOR2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_789), .Y(n_785) );
CKINVDCx5p33_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g794 ( .A(n_795), .Y(n_794) );
BUFx3_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_797), .Y(n_796) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_799), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_800), .Y(n_799) );
INVx3_ASAP7_75t_SL g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g809 ( .A(n_801), .Y(n_809) );
NAND2xp5_ASAP7_75t_SL g801 ( .A(n_802), .B(n_806), .Y(n_801) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
endmodule