module fake_aes_6722_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_33;
wire n_26;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_3), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_2), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_11), .B(n_0), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_17), .B(n_0), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
NAND2x1p5_ASAP7_75t_L g21 ( .A(n_13), .B(n_9), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_14), .Y(n_22) );
NOR3xp33_ASAP7_75t_SL g23 ( .A(n_13), .B(n_2), .C(n_3), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_14), .Y(n_24) );
INVxp67_ASAP7_75t_SL g25 ( .A(n_20), .Y(n_25) );
NAND2xp33_ASAP7_75t_R g26 ( .A(n_23), .B(n_15), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_22), .B(n_16), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_18), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
INVx2_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
NAND4xp25_ASAP7_75t_L g33 ( .A(n_30), .B(n_28), .C(n_19), .D(n_16), .Y(n_33) );
NOR2xp67_ASAP7_75t_L g34 ( .A(n_33), .B(n_30), .Y(n_34) );
AOI222xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_24), .B1(n_26), .B2(n_21), .C1(n_7), .C2(n_6), .Y(n_35) );
OAI21xp33_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_24), .B(n_5), .Y(n_36) );
AOI22xp33_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_34), .B1(n_24), .B2(n_4), .Y(n_37) );
endmodule