module real_aes_17045_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_1404;
wire n_602;
wire n_402;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1605;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_1292;
wire n_518;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_892;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1647;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_0), .A2(n_93), .B1(n_1450), .B2(n_1451), .Y(n_1473) );
AND2x2_ASAP7_75t_L g375 ( .A(n_1), .B(n_218), .Y(n_375) );
AND2x2_ASAP7_75t_L g394 ( .A(n_1), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g420 ( .A(n_1), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g1013 ( .A(n_1), .B(n_419), .Y(n_1013) );
AOI22xp33_ASAP7_75t_SL g704 ( .A1(n_2), .A2(n_274), .B1(n_384), .B2(n_649), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_2), .A2(n_3), .B1(n_417), .B2(n_725), .C(n_726), .Y(n_724) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_3), .A2(n_8), .B1(n_593), .B2(n_648), .Y(n_711) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_4), .A2(n_271), .B1(n_646), .B2(n_649), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g669 ( .A1(n_4), .A2(n_229), .B1(n_552), .B2(n_670), .C(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g837 ( .A(n_5), .Y(n_837) );
INVx1_ASAP7_75t_L g1284 ( .A(n_6), .Y(n_1284) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_6), .A2(n_301), .B1(n_456), .B2(n_759), .Y(n_1302) );
CKINVDCx5p33_ASAP7_75t_R g1320 ( .A(n_7), .Y(n_1320) );
A2O1A1Ixp33_ASAP7_75t_L g737 ( .A1(n_8), .A2(n_738), .B(n_739), .C(n_745), .Y(n_737) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_9), .A2(n_193), .B1(n_353), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g1192 ( .A1(n_10), .A2(n_195), .B1(n_652), .B2(n_829), .Y(n_1192) );
INVxp67_ASAP7_75t_SL g1218 ( .A(n_10), .Y(n_1218) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_11), .Y(n_754) );
AND4x1_ASAP7_75t_L g805 ( .A(n_11), .B(n_756), .C(n_760), .D(n_786), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_12), .A2(n_286), .B1(n_557), .B2(n_615), .Y(n_1408) );
INVx1_ASAP7_75t_L g1424 ( .A(n_12), .Y(n_1424) );
INVx2_ASAP7_75t_L g335 ( .A(n_13), .Y(n_335) );
OAI22xp5_ASAP7_75t_SL g539 ( .A1(n_14), .A2(n_249), .B1(n_540), .B2(n_542), .Y(n_539) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_14), .A2(n_249), .B1(n_392), .B2(n_428), .C(n_562), .Y(n_561) );
XNOR2x1_ASAP7_75t_L g508 ( .A(n_15), .B(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g1096 ( .A(n_16), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1330 ( .A1(n_17), .A2(n_120), .B1(n_1331), .B2(n_1333), .Y(n_1330) );
AOI22xp33_ASAP7_75t_L g1346 ( .A1(n_17), .A2(n_152), .B1(n_548), .B2(n_683), .Y(n_1346) );
INVx1_ASAP7_75t_L g1092 ( .A(n_18), .Y(n_1092) );
INVx1_ASAP7_75t_L g891 ( .A(n_19), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g1079 ( .A1(n_20), .A2(n_88), .B1(n_526), .B2(n_600), .C(n_949), .Y(n_1079) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_20), .A2(n_41), .B1(n_684), .B2(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g889 ( .A(n_21), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_21), .A2(n_64), .B1(n_903), .B2(n_904), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g758 ( .A1(n_22), .A2(n_149), .B1(n_456), .B2(n_759), .Y(n_758) );
OAI211xp5_ASAP7_75t_L g761 ( .A1(n_22), .A2(n_446), .B(n_762), .C(n_765), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_23), .A2(n_186), .B1(n_503), .B2(n_839), .Y(n_1341) );
INVx1_ASAP7_75t_L g1348 ( .A(n_23), .Y(n_1348) );
AOI22xp33_ASAP7_75t_SL g1337 ( .A1(n_24), .A2(n_84), .B1(n_593), .B2(n_1329), .Y(n_1337) );
AOI22xp33_ASAP7_75t_SL g1356 ( .A1(n_24), .A2(n_209), .B1(n_847), .B2(n_1357), .Y(n_1356) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_25), .A2(n_87), .B1(n_684), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_25), .A2(n_32), .B1(n_794), .B2(n_796), .Y(n_797) );
INVx1_ASAP7_75t_L g560 ( .A(n_26), .Y(n_560) );
HB1xp67_ASAP7_75t_L g1072 ( .A(n_27), .Y(n_1072) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_27), .B(n_1074), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_28), .Y(n_1178) );
INVx1_ASAP7_75t_L g338 ( .A(n_29), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g389 ( .A1(n_29), .A2(n_390), .B(n_398), .C(n_421), .Y(n_389) );
INVxp67_ASAP7_75t_L g636 ( .A(n_30), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g757 ( .A(n_31), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g784 ( .A1(n_32), .A2(n_292), .B1(n_412), .B2(n_624), .C(n_785), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g1251 ( .A1(n_33), .A2(n_48), .B1(n_528), .B2(n_800), .Y(n_1251) );
INVx1_ASAP7_75t_L g1262 ( .A(n_33), .Y(n_1262) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_34), .A2(n_63), .B1(n_1445), .B2(n_1458), .Y(n_1472) );
INVx1_ASAP7_75t_L g1022 ( .A(n_35), .Y(n_1022) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_36), .A2(n_45), .B1(n_988), .B2(n_989), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1041 ( .A1(n_36), .A2(n_147), .B1(n_597), .B2(n_799), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_37), .A2(n_96), .B1(n_642), .B2(n_706), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g740 ( .A1(n_37), .A2(n_176), .B1(n_575), .B2(n_673), .C(n_741), .Y(n_740) );
AOI221xp5_ASAP7_75t_L g437 ( .A1(n_38), .A2(n_268), .B1(n_412), .B2(n_438), .C(n_439), .Y(n_437) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_38), .Y(n_468) );
INVx1_ASAP7_75t_L g382 ( .A(n_39), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_39), .A2(n_187), .B1(n_443), .B2(n_446), .Y(n_442) );
AOI221xp5_ASAP7_75t_L g1241 ( .A1(n_40), .A2(n_303), .B1(n_349), .B2(n_1242), .C(n_1243), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1260 ( .A1(n_40), .A2(n_118), .B1(n_623), .B2(n_845), .C(n_1261), .Y(n_1260) );
AOI221xp5_ASAP7_75t_L g1080 ( .A1(n_41), .A2(n_67), .B1(n_526), .B2(n_949), .C(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_42), .A2(n_248), .B1(n_598), .B2(n_655), .Y(n_1190) );
INVx1_ASAP7_75t_L g1209 ( .A(n_42), .Y(n_1209) );
INVx1_ASAP7_75t_L g1411 ( .A(n_43), .Y(n_1411) );
NAND5xp2_ASAP7_75t_L g920 ( .A(n_44), .B(n_921), .C(n_943), .D(n_956), .E(n_964), .Y(n_920) );
INVx1_ASAP7_75t_L g972 ( .A(n_44), .Y(n_972) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_45), .A2(n_155), .B1(n_826), .B2(n_1035), .Y(n_1034) );
INVx1_ASAP7_75t_L g1410 ( .A(n_46), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g1289 ( .A1(n_47), .A2(n_166), .B1(n_677), .B2(n_683), .Y(n_1289) );
AOI22xp33_ASAP7_75t_SL g1309 ( .A1(n_47), .A2(n_280), .B1(n_792), .B2(n_946), .Y(n_1309) );
INVx1_ASAP7_75t_L g1256 ( .A(n_48), .Y(n_1256) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_49), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_49), .A2(n_132), .B1(n_500), .B2(n_501), .Y(n_499) );
INVxp67_ASAP7_75t_L g1318 ( .A(n_50), .Y(n_1318) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_51), .Y(n_380) );
INVx1_ASAP7_75t_L g763 ( .A(n_52), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g788 ( .A1(n_52), .A2(n_102), .B1(n_713), .B2(n_789), .Y(n_788) );
INVx1_ASAP7_75t_L g1084 ( .A(n_53), .Y(n_1084) );
AOI22xp33_ASAP7_75t_SL g1144 ( .A1(n_53), .A2(n_223), .B1(n_615), .B2(n_617), .Y(n_1144) );
XOR2x2_ASAP7_75t_L g1276 ( .A(n_54), .B(n_1277), .Y(n_1276) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_54), .A2(n_113), .B1(n_1445), .B2(n_1458), .Y(n_1457) );
AOI22xp5_ASAP7_75t_L g1478 ( .A1(n_55), .A2(n_222), .B1(n_1445), .B2(n_1458), .Y(n_1478) );
INVx1_ASAP7_75t_L g1186 ( .A(n_56), .Y(n_1186) );
INVx1_ASAP7_75t_L g559 ( .A(n_57), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_58), .A2(n_154), .B1(n_396), .B2(n_412), .C(n_439), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_58), .A2(n_205), .B1(n_597), .B2(n_949), .Y(n_948) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_59), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_60), .A2(n_205), .B1(n_557), .B2(n_771), .Y(n_927) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_60), .A2(n_154), .B1(n_597), .B2(n_598), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_61), .A2(n_146), .B1(n_641), .B2(n_655), .Y(n_654) );
AOI21xp33_ASAP7_75t_L g685 ( .A1(n_61), .A2(n_624), .B(n_686), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_62), .A2(n_291), .B1(n_686), .B2(n_767), .C(n_769), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g798 ( .A1(n_62), .A2(n_263), .B1(n_799), .B2(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g879 ( .A(n_64), .Y(n_879) );
INVx1_ASAP7_75t_L g701 ( .A(n_65), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_66), .A2(n_288), .B1(n_991), .B2(n_994), .C(n_996), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_66), .A2(n_257), .B1(n_538), .B2(n_1038), .C(n_1040), .Y(n_1037) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_67), .A2(n_88), .B1(n_551), .B2(n_623), .Y(n_1145) );
AOI22xp33_ASAP7_75t_SL g1188 ( .A1(n_68), .A2(n_156), .B1(n_538), .B2(n_646), .Y(n_1188) );
INVxp67_ASAP7_75t_SL g1215 ( .A(n_68), .Y(n_1215) );
OAI211xp5_ASAP7_75t_SL g1232 ( .A1(n_69), .A2(n_1050), .B(n_1057), .C(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1267 ( .A(n_69), .Y(n_1267) );
CKINVDCx5p33_ASAP7_75t_R g659 ( .A(n_70), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g692 ( .A1(n_71), .A2(n_456), .B(n_693), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g934 ( .A(n_72), .Y(n_934) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_73), .A2(n_203), .B1(n_822), .B2(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_SL g862 ( .A1(n_73), .A2(n_256), .B1(n_615), .B2(n_684), .Y(n_862) );
INVxp67_ASAP7_75t_SL g1028 ( .A(n_74), .Y(n_1028) );
OAI22xp5_ASAP7_75t_L g1042 ( .A1(n_74), .A2(n_298), .B1(n_1043), .B2(n_1046), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1485 ( .A1(n_75), .A2(n_213), .B1(n_1445), .B2(n_1458), .Y(n_1485) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_76), .A2(n_229), .B1(n_648), .B2(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_76), .A2(n_271), .B1(n_683), .B2(n_684), .Y(n_682) );
OR2x2_ASAP7_75t_L g364 ( .A(n_77), .B(n_365), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_78), .A2(n_185), .B1(n_424), .B2(n_428), .C(n_433), .Y(n_423) );
OAI322xp33_ASAP7_75t_L g466 ( .A1(n_78), .A2(n_467), .A3(n_475), .B1(n_478), .B2(n_486), .C1(n_492), .C2(n_503), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g1466 ( .A1(n_79), .A2(n_217), .B1(n_1450), .B2(n_1451), .Y(n_1466) );
AOI22xp33_ASAP7_75t_SL g596 ( .A1(n_80), .A2(n_181), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_80), .A2(n_92), .B1(n_615), .B2(n_617), .Y(n_614) );
AOI22xp33_ASAP7_75t_SL g827 ( .A1(n_81), .A2(n_197), .B1(n_824), .B2(n_826), .Y(n_827) );
INVx1_ASAP7_75t_L g854 ( .A(n_81), .Y(n_854) );
INVx1_ASAP7_75t_L g512 ( .A(n_82), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_83), .A2(n_253), .B1(n_523), .B2(n_524), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g550 ( .A1(n_83), .A2(n_95), .B1(n_416), .B2(n_551), .C(n_552), .Y(n_550) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_84), .A2(n_276), .B1(n_412), .B2(n_417), .C(n_1296), .Y(n_1345) );
INVx1_ASAP7_75t_L g1220 ( .A(n_85), .Y(n_1220) );
AOI22xp5_ASAP7_75t_L g1467 ( .A1(n_85), .A2(n_106), .B1(n_1445), .B2(n_1468), .Y(n_1467) );
AO22x1_ASAP7_75t_L g1449 ( .A1(n_86), .A2(n_224), .B1(n_1450), .B2(n_1451), .Y(n_1449) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_87), .A2(n_292), .B1(n_794), .B2(n_796), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_89), .A2(n_240), .B1(n_524), .B2(n_946), .Y(n_1383) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_89), .A2(n_235), .B1(n_417), .B2(n_613), .C(n_845), .Y(n_1388) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_90), .A2(n_172), .B1(n_1087), .B2(n_1088), .Y(n_1086) );
INVx1_ASAP7_75t_L g1114 ( .A(n_90), .Y(n_1114) );
INVx1_ASAP7_75t_L g515 ( .A(n_91), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g604 ( .A1(n_92), .A2(n_255), .B1(n_597), .B2(n_598), .Y(n_604) );
INVx1_ASAP7_75t_L g1375 ( .A(n_94), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1389 ( .A1(n_94), .A2(n_261), .B1(n_617), .B2(n_683), .Y(n_1389) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_95), .A2(n_169), .B1(n_500), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_96), .A2(n_130), .B1(n_615), .B2(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g888 ( .A(n_97), .Y(n_888) );
AOI221xp5_ASAP7_75t_L g897 ( .A1(n_97), .A2(n_198), .B1(n_438), .B2(n_624), .C(n_670), .Y(n_897) );
INVx1_ASAP7_75t_L g1100 ( .A(n_98), .Y(n_1100) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_99), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_100), .Y(n_667) );
XNOR2xp5_ASAP7_75t_L g1400 ( .A(n_101), .B(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g764 ( .A(n_102), .Y(n_764) );
OAI211xp5_ASAP7_75t_L g930 ( .A1(n_103), .A2(n_855), .B(n_931), .C(n_933), .Y(n_930) );
INVx1_ASAP7_75t_L g968 ( .A(n_103), .Y(n_968) );
INVx1_ASAP7_75t_L g434 ( .A(n_104), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_105), .Y(n_662) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_105), .A2(n_121), .B1(n_689), .B2(n_690), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g1415 ( .A1(n_107), .A2(n_845), .B(n_1416), .Y(n_1415) );
INVx1_ASAP7_75t_L g1423 ( .A(n_107), .Y(n_1423) );
INVx1_ASAP7_75t_L g1365 ( .A(n_108), .Y(n_1365) );
OAI221xp5_ASAP7_75t_L g772 ( .A1(n_109), .A2(n_237), .B1(n_773), .B2(n_774), .C(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g804 ( .A(n_109), .Y(n_804) );
INVx1_ASAP7_75t_L g1074 ( .A(n_110), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g1405 ( .A1(n_111), .A2(n_221), .B1(n_417), .B2(n_623), .C(n_1406), .Y(n_1405) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_111), .A2(n_158), .B1(n_348), .B2(n_946), .Y(n_1425) );
INVx1_ASAP7_75t_L g585 ( .A(n_112), .Y(n_585) );
INVx1_ASAP7_75t_L g583 ( .A(n_114), .Y(n_583) );
AO221x2_ASAP7_75t_L g1539 ( .A1(n_115), .A2(n_289), .B1(n_1450), .B2(n_1451), .C(n_1540), .Y(n_1539) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_116), .A2(n_254), .B1(n_500), .B2(n_593), .C(n_594), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_116), .A2(n_201), .B1(n_552), .B2(n_573), .C(n_613), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_117), .A2(n_163), .B1(n_526), .B2(n_598), .Y(n_1189) );
INVx1_ASAP7_75t_L g1213 ( .A(n_117), .Y(n_1213) );
INVx1_ASAP7_75t_L g1248 ( .A(n_118), .Y(n_1248) );
OAI22xp33_ASAP7_75t_L g874 ( .A1(n_119), .A2(n_265), .B1(n_713), .B2(n_789), .Y(n_874) );
INVx1_ASAP7_75t_L g907 ( .A(n_119), .Y(n_907) );
AOI21xp33_ASAP7_75t_L g1355 ( .A1(n_120), .A2(n_439), .B(n_672), .Y(n_1355) );
CKINVDCx5p33_ASAP7_75t_R g661 ( .A(n_121), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_122), .Y(n_1380) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_123), .A2(n_153), .B1(n_1061), .B2(n_1064), .Y(n_1060) );
INVxp67_ASAP7_75t_SL g1067 ( .A(n_123), .Y(n_1067) );
INVx1_ASAP7_75t_L g880 ( .A(n_124), .Y(n_880) );
AOI221xp5_ASAP7_75t_L g900 ( .A1(n_124), .A2(n_246), .B1(n_438), .B2(n_741), .C(n_901), .Y(n_900) );
INVxp67_ASAP7_75t_SL g1292 ( .A(n_125), .Y(n_1292) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_125), .A2(n_226), .B1(n_1311), .B2(n_1312), .Y(n_1310) );
INVx1_ASAP7_75t_L g1371 ( .A(n_126), .Y(n_1371) );
AOI21xp33_ASAP7_75t_L g1396 ( .A1(n_126), .A2(n_624), .B(n_845), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_127), .A2(n_151), .B1(n_514), .B2(n_759), .Y(n_1366) );
OAI211xp5_ASAP7_75t_L g1386 ( .A1(n_127), .A2(n_842), .B(n_1387), .C(n_1390), .Y(n_1386) );
INVx1_ASAP7_75t_L g1182 ( .A(n_128), .Y(n_1182) );
OAI222xp33_ASAP7_75t_L g1207 ( .A1(n_128), .A2(n_184), .B1(n_390), .B2(n_774), .C1(n_1208), .C2(n_1214), .Y(n_1207) );
INVx1_ASAP7_75t_L g1283 ( .A(n_129), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g1315 ( .A1(n_129), .A2(n_157), .B1(n_789), .B2(n_839), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_130), .A2(n_176), .B1(n_642), .B2(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_SL g1287 ( .A(n_131), .Y(n_1287) );
AOI22xp33_ASAP7_75t_SL g1313 ( .A1(n_131), .A2(n_175), .B1(n_796), .B2(n_824), .Y(n_1313) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_132), .A2(n_194), .B1(n_412), .B2(n_416), .C(n_417), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g1231 ( .A1(n_133), .A2(n_309), .B1(n_1061), .B2(n_1064), .Y(n_1231) );
INVxp33_ASAP7_75t_SL g1271 ( .A(n_133), .Y(n_1271) );
AOI31xp33_ASAP7_75t_L g1076 ( .A1(n_134), .A2(n_1077), .A3(n_1085), .B(n_1112), .Y(n_1076) );
NAND2xp33_ASAP7_75t_SL g1140 ( .A(n_134), .B(n_1141), .Y(n_1140) );
INVxp67_ASAP7_75t_SL g1150 ( .A(n_134), .Y(n_1150) );
AO22x1_ASAP7_75t_L g1463 ( .A1(n_134), .A2(n_296), .B1(n_1450), .B2(n_1451), .Y(n_1463) );
INVx1_ASAP7_75t_L g813 ( .A(n_135), .Y(n_813) );
OAI221xp5_ASAP7_75t_L g851 ( .A1(n_135), .A2(n_136), .B1(n_775), .B2(n_852), .C(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g816 ( .A(n_136), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_137), .Y(n_1234) );
OA21x2_ASAP7_75t_L g510 ( .A1(n_138), .A2(n_365), .B(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g1238 ( .A(n_139), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g1254 ( .A1(n_139), .A2(n_214), .B1(n_623), .B2(n_845), .C(n_1255), .Y(n_1254) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_140), .A2(n_147), .B1(n_989), .B2(n_1008), .C(n_1009), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1036 ( .A1(n_140), .A2(n_288), .B1(n_595), .B2(n_822), .C(n_946), .Y(n_1036) );
INVx1_ASAP7_75t_L g1196 ( .A(n_141), .Y(n_1196) );
INVx1_ASAP7_75t_L g1323 ( .A(n_142), .Y(n_1323) );
OAI221xp5_ASAP7_75t_SL g1350 ( .A1(n_142), .A2(n_227), .B1(n_773), .B2(n_774), .C(n_1351), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g1412 ( .A1(n_143), .A2(n_299), .B1(n_775), .B2(n_852), .C(n_1413), .Y(n_1412) );
OAI22xp33_ASAP7_75t_L g1430 ( .A1(n_143), .A2(n_299), .B1(n_542), .B2(n_815), .Y(n_1430) );
AO22x1_ASAP7_75t_L g640 ( .A1(n_144), .A2(n_174), .B1(n_641), .B2(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_144), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g963 ( .A(n_145), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_146), .A2(n_174), .B1(n_676), .B2(n_677), .Y(n_675) );
AO22x1_ASAP7_75t_L g1444 ( .A1(n_148), .A2(n_297), .B1(n_1445), .B2(n_1447), .Y(n_1444) );
CKINVDCx16_ASAP7_75t_R g1541 ( .A(n_150), .Y(n_1541) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_152), .A2(n_269), .B1(n_1333), .B2(n_1335), .Y(n_1334) );
INVxp67_ASAP7_75t_SL g1018 ( .A(n_153), .Y(n_1018) );
INVx1_ASAP7_75t_L g1010 ( .A(n_155), .Y(n_1010) );
AOI221xp5_ASAP7_75t_L g1201 ( .A1(n_156), .A2(n_195), .B1(n_769), .B2(n_1202), .C(n_1203), .Y(n_1201) );
INVx1_ASAP7_75t_L g1281 ( .A(n_157), .Y(n_1281) );
AOI22xp33_ASAP7_75t_SL g1417 ( .A1(n_158), .A2(n_272), .B1(n_448), .B2(n_676), .Y(n_1417) );
OAI211xp5_ASAP7_75t_L g1403 ( .A1(n_159), .A2(n_842), .B(n_1404), .C(n_1409), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g1433 ( .A1(n_159), .A2(n_290), .B1(n_514), .B2(n_759), .Y(n_1433) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_160), .A2(n_258), .B1(n_824), .B2(n_826), .Y(n_823) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_160), .A2(n_197), .B1(n_617), .B2(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g520 ( .A(n_161), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_161), .A2(n_196), .B1(n_569), .B2(n_573), .C(n_575), .Y(n_568) );
OAI211xp5_ASAP7_75t_L g922 ( .A1(n_162), .A2(n_923), .B(n_924), .C(n_929), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g942 ( .A(n_162), .B(n_353), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1204 ( .A1(n_163), .A2(n_248), .B1(n_904), .B2(n_1205), .Y(n_1204) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_164), .A2(n_201), .B1(n_500), .B2(n_538), .C(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_164), .A2(n_254), .B1(n_617), .B2(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g1167 ( .A(n_165), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1448 ( .A(n_165), .B(n_262), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_165), .B(n_1168), .Y(n_1452) );
AOI22xp33_ASAP7_75t_SL g1314 ( .A1(n_166), .A2(n_307), .B1(n_801), .B2(n_946), .Y(n_1314) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_167), .Y(n_465) );
INVx1_ASAP7_75t_L g1392 ( .A(n_168), .Y(n_1392) );
INVx1_ASAP7_75t_L g567 ( .A(n_169), .Y(n_567) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_170), .A2(n_251), .B1(n_353), .B2(n_456), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g722 ( .A1(n_170), .A2(n_446), .B(n_723), .C(n_730), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g666 ( .A(n_171), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g1122 ( .A1(n_172), .A2(n_242), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
INVx1_ASAP7_75t_L g1340 ( .A(n_173), .Y(n_1340) );
INVxp67_ASAP7_75t_SL g1294 ( .A(n_175), .Y(n_1294) );
NOR2xp33_ASAP7_75t_L g1297 ( .A(n_177), .B(n_852), .Y(n_1297) );
INVx1_ASAP7_75t_L g1307 ( .A(n_177), .Y(n_1307) );
INVx1_ASAP7_75t_L g1195 ( .A(n_178), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_179), .A2(n_245), .B1(n_556), .B2(n_557), .Y(n_925) );
AOI22xp33_ASAP7_75t_SL g950 ( .A1(n_179), .A2(n_260), .B1(n_946), .B2(n_951), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_180), .A2(n_235), .B1(n_524), .B2(n_946), .Y(n_1376) );
AOI22xp33_ASAP7_75t_SL g1397 ( .A1(n_180), .A2(n_240), .B1(n_676), .B2(n_684), .Y(n_1397) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_181), .A2(n_255), .B1(n_573), .B2(n_623), .C(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g884 ( .A(n_182), .Y(n_884) );
INVx1_ASAP7_75t_L g536 ( .A(n_183), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_183), .A2(n_239), .B1(n_554), .B2(n_557), .Y(n_553) );
INVx1_ASAP7_75t_L g1183 ( .A(n_184), .Y(n_1183) );
INVx1_ASAP7_75t_L g324 ( .A(n_185), .Y(n_324) );
INVx1_ASAP7_75t_L g1349 ( .A(n_186), .Y(n_1349) );
INVx1_ASAP7_75t_L g351 ( .A(n_187), .Y(n_351) );
CKINVDCx5p33_ASAP7_75t_R g1414 ( .A(n_188), .Y(n_1414) );
OAI22xp5_ASAP7_75t_L g838 ( .A1(n_189), .A2(n_306), .B1(n_503), .B2(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g849 ( .A(n_189), .Y(n_849) );
INVx1_ASAP7_75t_L g506 ( .A(n_190), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g937 ( .A(n_191), .Y(n_937) );
INVx2_ASAP7_75t_L g337 ( .A(n_192), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_192), .B(n_335), .Y(n_372) );
INVx1_ASAP7_75t_L g491 ( .A(n_192), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g898 ( .A1(n_193), .A2(n_842), .B(n_899), .C(n_906), .Y(n_898) );
INVx1_ASAP7_75t_L g483 ( .A(n_194), .Y(n_483) );
INVx1_ASAP7_75t_L g535 ( .A(n_196), .Y(n_535) );
INVx1_ASAP7_75t_L g885 ( .A(n_198), .Y(n_885) );
INVx1_ASAP7_75t_L g410 ( .A(n_199), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g940 ( .A1(n_200), .A2(n_266), .B1(n_931), .B2(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g966 ( .A(n_200), .Y(n_966) );
BUFx3_ASAP7_75t_L g329 ( .A(n_202), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g844 ( .A1(n_203), .A2(n_211), .B1(n_417), .B2(n_613), .C(n_845), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1486 ( .A1(n_204), .A2(n_210), .B1(n_1450), .B2(n_1451), .Y(n_1486) );
INVx1_ASAP7_75t_L g610 ( .A(n_206), .Y(n_610) );
CKINVDCx5p33_ASAP7_75t_R g1235 ( .A(n_207), .Y(n_1235) );
OAI22xp5_ASAP7_75t_L g871 ( .A1(n_208), .A2(n_212), .B1(n_815), .B2(n_872), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g895 ( .A1(n_208), .A2(n_212), .B1(n_773), .B2(n_774), .C(n_896), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g1328 ( .A1(n_209), .A2(n_276), .B1(n_652), .B2(n_1329), .Y(n_1328) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_211), .A2(n_256), .B1(n_646), .B2(n_822), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_213), .A2(n_868), .B1(n_869), .B2(n_914), .Y(n_867) );
INVx1_ASAP7_75t_L g914 ( .A(n_213), .Y(n_914) );
AOI21xp33_ASAP7_75t_L g1250 ( .A1(n_214), .A2(n_495), .B(n_1040), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_215), .B(n_809), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_215), .A2(n_834), .B1(n_835), .B2(n_863), .Y(n_833) );
INVx1_ASAP7_75t_L g865 ( .A(n_215), .Y(n_865) );
OAI22xp33_ASAP7_75t_L g712 ( .A1(n_216), .A2(n_233), .B1(n_503), .B2(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g731 ( .A(n_216), .Y(n_731) );
INVx1_ASAP7_75t_L g395 ( .A(n_218), .Y(n_395) );
BUFx3_ASAP7_75t_L g419 ( .A(n_218), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g1543 ( .A(n_219), .Y(n_1543) );
AOI22xp5_ASAP7_75t_L g1477 ( .A1(n_220), .A2(n_234), .B1(n_1450), .B2(n_1451), .Y(n_1477) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_221), .A2(n_272), .B1(n_538), .B2(n_946), .Y(n_1429) );
XNOR2x1_ASAP7_75t_L g580 ( .A(n_222), .B(n_581), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g1078 ( .A1(n_223), .A2(n_252), .B1(n_500), .B2(n_792), .Y(n_1078) );
INVxp67_ASAP7_75t_SL g1326 ( .A(n_225), .Y(n_1326) );
OAI211xp5_ASAP7_75t_SL g1343 ( .A1(n_225), .A2(n_446), .B(n_1344), .C(n_1347), .Y(n_1343) );
AOI21xp5_ASAP7_75t_L g1290 ( .A1(n_226), .A2(n_439), .B(n_670), .Y(n_1290) );
INVx1_ASAP7_75t_L g1324 ( .A(n_227), .Y(n_1324) );
CKINVDCx5p33_ASAP7_75t_R g1240 ( .A(n_228), .Y(n_1240) );
INVx1_ASAP7_75t_L g609 ( .A(n_230), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_231), .Y(n_832) );
INVx1_ASAP7_75t_L g702 ( .A(n_232), .Y(n_702) );
INVx1_ASAP7_75t_L g734 ( .A(n_233), .Y(n_734) );
INVx1_ASAP7_75t_L g403 ( .A(n_236), .Y(n_403) );
INVx1_ASAP7_75t_L g803 ( .A(n_237), .Y(n_803) );
INVx1_ASAP7_75t_L g1391 ( .A(n_238), .Y(n_1391) );
NAND2xp33_ASAP7_75t_SL g525 ( .A(n_239), .B(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g1456 ( .A1(n_241), .A2(n_302), .B1(n_1450), .B2(n_1451), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1103 ( .A1(n_242), .A2(n_281), .B1(n_1104), .B2(n_1106), .Y(n_1103) );
AO22x1_ASAP7_75t_L g1462 ( .A1(n_243), .A2(n_250), .B1(n_1445), .B2(n_1458), .Y(n_1462) );
XNOR2x2_ASAP7_75t_L g696 ( .A(n_244), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_SL g945 ( .A1(n_245), .A2(n_311), .B1(n_524), .B2(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g892 ( .A(n_246), .Y(n_892) );
INVx1_ASAP7_75t_L g345 ( .A(n_247), .Y(n_345) );
INVx1_ASAP7_75t_L g359 ( .A(n_247), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_252), .A2(n_282), .B1(n_551), .B2(n_623), .Y(n_1146) );
INVx1_ASAP7_75t_L g564 ( .A(n_253), .Y(n_564) );
INVx1_ASAP7_75t_L g1011 ( .A(n_257), .Y(n_1011) );
AOI21xp33_ASAP7_75t_L g859 ( .A1(n_258), .A2(n_624), .B(n_860), .Y(n_859) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_259), .Y(n_588) );
AOI221xp5_ASAP7_75t_SL g928 ( .A1(n_260), .A2(n_311), .B1(n_396), .B2(n_552), .C(n_672), .Y(n_928) );
INVx1_ASAP7_75t_L g1382 ( .A(n_261), .Y(n_1382) );
INVx1_ASAP7_75t_L g1168 ( .A(n_262), .Y(n_1168) );
AND2x2_ASAP7_75t_L g1446 ( .A(n_262), .B(n_1167), .Y(n_1446) );
INVxp67_ASAP7_75t_SL g783 ( .A(n_263), .Y(n_783) );
OAI211xp5_ASAP7_75t_SL g1285 ( .A1(n_264), .A2(n_428), .B(n_1286), .C(n_1291), .Y(n_1285) );
INVx1_ASAP7_75t_L g1306 ( .A(n_264), .Y(n_1306) );
INVx1_ASAP7_75t_L g908 ( .A(n_265), .Y(n_908) );
INVx1_ASAP7_75t_L g955 ( .A(n_266), .Y(n_955) );
XNOR2xp5_ASAP7_75t_L g1223 ( .A(n_267), .B(n_1224), .Y(n_1223) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_268), .Y(n_496) );
INVx1_ASAP7_75t_L g1352 ( .A(n_269), .Y(n_1352) );
INVxp67_ASAP7_75t_SL g818 ( .A(n_270), .Y(n_818) );
OAI211xp5_ASAP7_75t_L g841 ( .A1(n_270), .A2(n_842), .B(n_843), .C(n_848), .Y(n_841) );
AOI22xp33_ASAP7_75t_SL g980 ( .A1(n_273), .A2(n_981), .B1(n_982), .B2(n_983), .Y(n_980) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_273), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_274), .B(n_743), .Y(n_742) );
OAI21xp33_ASAP7_75t_L g1193 ( .A1(n_275), .A2(n_456), .B(n_1194), .Y(n_1193) );
INVx1_ASAP7_75t_L g1226 ( .A(n_277), .Y(n_1226) );
OAI21xp5_ASAP7_75t_SL g627 ( .A1(n_278), .A2(n_514), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g1246 ( .A(n_279), .Y(n_1246) );
AOI221xp5_ASAP7_75t_L g1295 ( .A1(n_280), .A2(n_307), .B1(n_417), .B2(n_767), .C(n_1296), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1118 ( .A(n_281), .Y(n_1118) );
INVx1_ASAP7_75t_L g1083 ( .A(n_282), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g695 ( .A(n_283), .Y(n_695) );
INVxp67_ASAP7_75t_SL g779 ( .A(n_284), .Y(n_779) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_284), .A2(n_291), .B1(n_648), .B2(n_792), .Y(n_791) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_285), .Y(n_378) );
INVx1_ASAP7_75t_L g1428 ( .A(n_286), .Y(n_1428) );
INVx1_ASAP7_75t_L g1301 ( .A(n_287), .Y(n_1301) );
INVxp67_ASAP7_75t_SL g1026 ( .A(n_293), .Y(n_1026) );
OAI221xp5_ASAP7_75t_L g1052 ( .A1(n_293), .A2(n_295), .B1(n_1053), .B2(n_1055), .C(n_1057), .Y(n_1052) );
INVx1_ASAP7_75t_L g1432 ( .A(n_294), .Y(n_1432) );
OAI221xp5_ASAP7_75t_L g998 ( .A1(n_295), .A2(n_298), .B1(n_999), .B2(n_1004), .C(n_1005), .Y(n_998) );
INVx1_ASAP7_75t_L g332 ( .A(n_300), .Y(n_332) );
INVx1_ASAP7_75t_L g363 ( .A(n_300), .Y(n_363) );
INVx2_ASAP7_75t_L g453 ( .A(n_300), .Y(n_453) );
INVx1_ASAP7_75t_L g1257 ( .A(n_303), .Y(n_1257) );
CKINVDCx5p33_ASAP7_75t_R g911 ( .A(n_304), .Y(n_911) );
OAI22xp33_ASAP7_75t_SL g1384 ( .A1(n_305), .A2(n_310), .B1(n_542), .B2(n_815), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g1393 ( .A1(n_305), .A2(n_310), .B1(n_773), .B2(n_775), .C(n_1394), .Y(n_1393) );
INVx1_ASAP7_75t_L g850 ( .A(n_306), .Y(n_850) );
XNOR2xp5_ASAP7_75t_L g1362 ( .A(n_308), .B(n_1363), .Y(n_1362) );
INVxp67_ASAP7_75t_SL g1229 ( .A(n_309), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_1646), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_978), .Y(n_313) );
INVxp67_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AOI21xp33_ASAP7_75t_SL g1646 ( .A1(n_315), .A2(n_1647), .B(n_1649), .Y(n_1646) );
OAI22xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_915), .B1(n_976), .B2(n_977), .Y(n_315) );
INVx1_ASAP7_75t_L g976 ( .A(n_316), .Y(n_976) );
XOR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_751), .Y(n_316) );
XOR2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_633), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B1(n_507), .B2(n_632), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
XNOR2x1_ASAP7_75t_L g320 ( .A(n_321), .B(n_506), .Y(n_320) );
NOR2x1_ASAP7_75t_L g321 ( .A(n_322), .B(n_387), .Y(n_321) );
NAND5xp2_ASAP7_75t_L g322 ( .A(n_323), .B(n_346), .C(n_350), .D(n_364), .E(n_381), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_325), .B1(n_338), .B2(n_339), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_325), .A2(n_339), .B1(n_661), .B2(n_662), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_325), .A2(n_339), .B1(n_701), .B2(n_702), .Y(n_700) );
AO22x1_ASAP7_75t_L g1181 ( .A1(n_325), .A2(n_339), .B1(n_1182), .B2(n_1183), .Y(n_1181) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_330), .Y(n_325) );
AND2x2_ASAP7_75t_L g541 ( .A(n_326), .B(n_330), .Y(n_541) );
AND2x4_ASAP7_75t_SL g589 ( .A(n_326), .B(n_330), .Y(n_589) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_326), .B(n_330), .Y(n_815) );
AND2x6_ASAP7_75t_L g1054 ( .A(n_326), .B(n_333), .Y(n_1054) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_328), .B(n_464), .Y(n_463) );
AND2x4_ASAP7_75t_L g528 ( .A(n_328), .B(n_343), .Y(n_528) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_328), .Y(n_1099) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g349 ( .A(n_329), .B(n_344), .Y(n_349) );
INVx2_ASAP7_75t_L g356 ( .A(n_329), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_329), .B(n_345), .Y(n_369) );
OR2x2_ASAP7_75t_L g482 ( .A(n_329), .B(n_358), .Y(n_482) );
AND2x4_ASAP7_75t_L g339 ( .A(n_330), .B(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_L g347 ( .A(n_330), .B(n_348), .Y(n_347) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_330), .B(n_340), .Y(n_543) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
OR2x2_ASAP7_75t_L g373 ( .A(n_331), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g1016 ( .A(n_331), .Y(n_1016) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g490 ( .A(n_332), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g1021 ( .A(n_332), .B(n_394), .Y(n_1021) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_333), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g1056 ( .A(n_333), .B(n_342), .Y(n_1056) );
INVx1_ASAP7_75t_L g1059 ( .A(n_333), .Y(n_1059) );
AND2x4_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
NAND3x1_ASAP7_75t_L g489 ( .A(n_334), .B(n_490), .C(n_491), .Y(n_489) );
NAND2x1p5_ASAP7_75t_L g595 ( .A(n_334), .B(n_491), .Y(n_595) );
OR2x4_ASAP7_75t_L g1087 ( .A(n_334), .B(n_482), .Y(n_1087) );
INVx1_ASAP7_75t_L g1089 ( .A(n_334), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1094 ( .A(n_334), .B(n_349), .Y(n_1094) );
OR2x6_ASAP7_75t_L g1106 ( .A(n_334), .B(n_498), .Y(n_1106) );
INVx3_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp33_ASAP7_75t_SL g477 ( .A(n_335), .B(n_337), .Y(n_477) );
BUFx3_ASAP7_75t_L g602 ( .A(n_335), .Y(n_602) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND3x4_ASAP7_75t_L g601 ( .A(n_337), .B(n_602), .C(n_603), .Y(n_601) );
HB1xp67_ASAP7_75t_L g1109 ( .A(n_337), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_339), .A2(n_541), .B1(n_803), .B2(n_804), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g812 ( .A1(n_339), .A2(n_813), .B1(n_814), .B2(n_816), .Y(n_812) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_339), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_339), .A2(n_541), .B1(n_1306), .B2(n_1307), .Y(n_1305) );
AOI22xp5_ASAP7_75t_L g1322 ( .A1(n_339), .A2(n_541), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g464 ( .A(n_345), .Y(n_464) );
NAND3xp33_ASAP7_75t_SL g586 ( .A(n_346), .B(n_587), .C(n_591), .Y(n_586) );
AND4x1_ASAP7_75t_L g786 ( .A(n_346), .B(n_787), .C(n_790), .D(n_802), .Y(n_786) );
INVx2_ASAP7_75t_SL g893 ( .A(n_346), .Y(n_893) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR3xp33_ASAP7_75t_SL g516 ( .A(n_347), .B(n_517), .C(n_539), .Y(n_516) );
INVx3_ASAP7_75t_L g657 ( .A(n_347), .Y(n_657) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_347), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_347), .A2(n_543), .B1(n_589), .B2(n_934), .C(n_955), .Y(n_954) );
NOR3xp33_ASAP7_75t_L g1419 ( .A(n_347), .B(n_1420), .C(n_1430), .Y(n_1419) );
BUFx2_ASAP7_75t_L g649 ( .A(n_348), .Y(n_649) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g502 ( .A(n_349), .Y(n_502) );
BUFx2_ASAP7_75t_L g524 ( .A(n_349), .Y(n_524) );
BUFx2_ASAP7_75t_L g593 ( .A(n_349), .Y(n_593) );
BUFx2_ASAP7_75t_L g792 ( .A(n_349), .Y(n_792) );
BUFx3_ASAP7_75t_L g822 ( .A(n_349), .Y(n_822) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_349), .B(n_1045), .Y(n_1047) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_352), .A2(n_512), .B1(n_513), .B2(n_515), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g582 ( .A1(n_352), .A2(n_583), .B1(n_584), .B2(n_585), .C(n_586), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_352), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx5_ASAP7_75t_L g819 ( .A(n_353), .Y(n_819) );
OR2x6_ASAP7_75t_L g353 ( .A(n_354), .B(n_360), .Y(n_353) );
OR2x2_ASAP7_75t_L g759 ( .A(n_354), .B(n_360), .Y(n_759) );
INVx2_ASAP7_75t_L g1051 ( .A(n_354), .Y(n_1051) );
INVx8_ASAP7_75t_L g385 ( .A(n_355), .Y(n_385) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_355), .Y(n_523) );
BUFx3_ASAP7_75t_L g648 ( .A(n_355), .Y(n_648) );
BUFx3_ASAP7_75t_L g800 ( .A(n_355), .Y(n_800) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_355), .B(n_1045), .Y(n_1044) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
AND2x4_ASAP7_75t_L g471 ( .A(n_356), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVxp67_ASAP7_75t_L g472 ( .A(n_359), .Y(n_472) );
INVxp67_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g457 ( .A(n_361), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g961 ( .A(n_361), .Y(n_961) );
OR2x2_ASAP7_75t_L g1004 ( .A(n_361), .B(n_458), .Y(n_1004) );
INVx1_ASAP7_75t_L g1136 ( .A(n_361), .Y(n_1136) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g371 ( .A(n_362), .Y(n_371) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx8_ASAP7_75t_L g584 ( .A(n_365), .Y(n_584) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_373), .Y(n_365) );
INVx1_ASAP7_75t_L g967 ( .A(n_366), .Y(n_967) );
OR2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_370), .Y(n_366) );
BUFx3_ASAP7_75t_L g1239 ( .A(n_367), .Y(n_1239) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_368), .Y(n_474) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
BUFx2_ASAP7_75t_L g498 ( .A(n_369), .Y(n_498) );
INVx1_ASAP7_75t_L g386 ( .A(n_370), .Y(n_386) );
OR2x2_ASAP7_75t_L g461 ( .A(n_370), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g631 ( .A(n_370), .Y(n_631) );
OR2x2_ASAP7_75t_L g370 ( .A(n_371), .B(n_372), .Y(n_370) );
OR2x2_ASAP7_75t_L g476 ( .A(n_371), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_SL g997 ( .A(n_371), .B(n_418), .Y(n_997) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_371), .Y(n_1111) );
INVx1_ASAP7_75t_L g1265 ( .A(n_371), .Y(n_1265) );
INVx1_ASAP7_75t_L g1045 ( .A(n_372), .Y(n_1045) );
INVx1_ASAP7_75t_L g1063 ( .A(n_372), .Y(n_1063) );
INVx1_ASAP7_75t_L g1017 ( .A(n_374), .Y(n_1017) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
AND2x6_ASAP7_75t_L g422 ( .A(n_375), .B(n_396), .Y(n_422) );
INVx1_ASAP7_75t_L g432 ( .A(n_375), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_375), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g625 ( .A(n_375), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g1001 ( .A(n_375), .B(n_453), .Y(n_1001) );
AND2x2_ASAP7_75t_L g445 ( .A(n_376), .B(n_394), .Y(n_445) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_376), .Y(n_556) );
INVx3_ASAP7_75t_L g616 ( .A(n_376), .Y(n_616) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_377), .Y(n_936) );
OR2x2_ASAP7_75t_L g993 ( .A(n_377), .B(n_380), .Y(n_993) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x2_ASAP7_75t_L g397 ( .A(n_378), .B(n_380), .Y(n_397) );
OR2x2_ASAP7_75t_L g402 ( .A(n_378), .B(n_380), .Y(n_402) );
INVx2_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
AND2x2_ASAP7_75t_L g414 ( .A(n_378), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g460 ( .A(n_378), .Y(n_460) );
NAND2x1_ASAP7_75t_L g858 ( .A(n_378), .B(n_380), .Y(n_858) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_380), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g415 ( .A(n_380), .Y(n_415) );
BUFx2_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
AND2x2_ASAP7_75t_L g449 ( .A(n_380), .B(n_409), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_383), .A2(n_559), .B1(n_560), .B2(n_579), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_383), .A2(n_504), .B1(n_666), .B2(n_667), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_383), .A2(n_504), .B1(n_1195), .B2(n_1196), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1398 ( .A1(n_383), .A2(n_504), .B1(n_1391), .B2(n_1392), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1434 ( .A1(n_383), .A2(n_504), .B1(n_1410), .B2(n_1411), .Y(n_1434) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_386), .Y(n_383) );
AND2x4_ASAP7_75t_L g629 ( .A(n_384), .B(n_386), .Y(n_629) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g500 ( .A(n_385), .Y(n_500) );
INVx3_ASAP7_75t_L g829 ( .A(n_385), .Y(n_829) );
INVx8_ASAP7_75t_L g946 ( .A(n_385), .Y(n_946) );
CKINVDCx5p33_ASAP7_75t_R g1242 ( .A(n_385), .Y(n_1242) );
AND2x4_ASAP7_75t_L g504 ( .A(n_386), .B(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_454), .Y(n_387) );
OAI31xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_423), .A3(n_442), .B(n_450), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_391), .A2(n_429), .B1(n_701), .B2(n_702), .Y(n_745) );
INVx2_ASAP7_75t_L g773 ( .A(n_391), .Y(n_773) );
INVx2_ASAP7_75t_L g852 ( .A(n_391), .Y(n_852) );
INVx4_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
BUFx3_ASAP7_75t_L g619 ( .A(n_393), .Y(n_619) );
AND2x4_ASAP7_75t_SL g393 ( .A(n_394), .B(n_396), .Y(n_393) );
AND2x4_ASAP7_75t_L g426 ( .A(n_394), .B(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g447 ( .A(n_394), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g547 ( .A(n_394), .B(n_548), .Y(n_547) );
BUFx2_ASAP7_75t_L g939 ( .A(n_394), .Y(n_939) );
AND2x2_ASAP7_75t_L g962 ( .A(n_394), .B(n_427), .Y(n_962) );
HB1xp67_ASAP7_75t_L g1120 ( .A(n_395), .Y(n_1120) );
BUFx3_ASAP7_75t_L g416 ( .A(n_396), .Y(n_416) );
BUFx3_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_396), .Y(n_613) );
BUFx3_ASAP7_75t_L g623 ( .A(n_396), .Y(n_623) );
INVx1_ASAP7_75t_L g687 ( .A(n_396), .Y(n_687) );
BUFx3_ASAP7_75t_L g1296 ( .A(n_396), .Y(n_1296) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g572 ( .A(n_397), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_403), .B1(n_404), .B2(n_410), .C(n_411), .Y(n_398) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_399), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_437), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g896 ( .A1(n_399), .A2(n_780), .B1(n_884), .B2(n_891), .C(n_897), .Y(n_896) );
INVx1_ASAP7_75t_L g989 ( .A(n_399), .Y(n_989) );
OAI221xp5_ASAP7_75t_L g1291 ( .A1(n_399), .A2(n_1292), .B1(n_1293), .B2(n_1294), .C(n_1295), .Y(n_1291) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g563 ( .A(n_400), .Y(n_563) );
INVx2_ASAP7_75t_SL g778 ( .A(n_400), .Y(n_778) );
OR2x6_ASAP7_75t_L g1116 ( .A(n_400), .B(n_1117), .Y(n_1116) );
OAI22xp5_ASAP7_75t_L g1255 ( .A1(n_400), .A2(n_1256), .B1(n_1257), .B2(n_1258), .Y(n_1255) );
OAI22x1_ASAP7_75t_SL g1261 ( .A1(n_400), .A2(n_1240), .B1(n_1258), .B2(n_1262), .Y(n_1261) );
INVx3_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g744 ( .A(n_401), .Y(n_744) );
BUFx4f_ASAP7_75t_L g932 ( .A(n_401), .Y(n_932) );
INVx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_403), .A2(n_468), .B1(n_469), .B2(n_473), .Y(n_467) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_405), .Y(n_1293) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g566 ( .A(n_406), .Y(n_566) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_406), .Y(n_738) );
INVx2_ASAP7_75t_L g782 ( .A(n_406), .Y(n_782) );
INVx2_ASAP7_75t_L g1258 ( .A(n_406), .Y(n_1258) );
INVx8_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx2_ASAP7_75t_L g435 ( .A(n_407), .Y(n_435) );
OR2x2_ASAP7_75t_L g1124 ( .A(n_407), .B(n_1125), .Y(n_1124) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g492 ( .A1(n_410), .A2(n_493), .B1(n_496), .B2(n_497), .C(n_499), .Y(n_492) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g672 ( .A(n_413), .Y(n_672) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_414), .Y(n_427) );
BUFx3_ASAP7_75t_L g845 ( .A(n_414), .Y(n_845) );
AND2x4_ASAP7_75t_L g1119 ( .A(n_414), .B(n_1120), .Y(n_1119) );
HB1xp67_ASAP7_75t_SL g901 ( .A(n_417), .Y(n_901) );
INVx4_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx4_ASAP7_75t_L g552 ( .A(n_418), .Y(n_552) );
INVx1_ASAP7_75t_SL g769 ( .A(n_418), .Y(n_769) );
AND2x4_ASAP7_75t_L g1263 ( .A(n_418), .B(n_1264), .Y(n_1263) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx2_ASAP7_75t_L g441 ( .A(n_419), .Y(n_441) );
AND2x4_ASAP7_75t_L g1129 ( .A(n_419), .B(n_459), .Y(n_1129) );
AND2x4_ASAP7_75t_L g440 ( .A(n_420), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g1135 ( .A(n_420), .Y(n_1135) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_422), .A2(n_515), .B1(n_547), .B2(n_550), .C(n_553), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_422), .A2(n_547), .B1(n_583), .B2(n_612), .C(n_614), .Y(n_611) );
AOI221xp5_ASAP7_75t_SL g668 ( .A1(n_422), .A2(n_447), .B1(n_659), .B2(n_669), .C(n_675), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g723 ( .A1(n_422), .A2(n_724), .B(n_728), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_422), .A2(n_766), .B(n_770), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g843 ( .A1(n_422), .A2(n_844), .B(n_846), .Y(n_843) );
AOI21xp5_ASAP7_75t_L g899 ( .A1(n_422), .A2(n_900), .B(n_902), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g1200 ( .A1(n_422), .A2(n_1201), .B(n_1204), .Y(n_1200) );
AOI21xp5_ASAP7_75t_L g1280 ( .A1(n_422), .A2(n_425), .B(n_1281), .Y(n_1280) );
AOI21xp5_ASAP7_75t_L g1344 ( .A1(n_422), .A2(n_1345), .B(n_1346), .Y(n_1344) );
AOI21xp5_ASAP7_75t_L g1387 ( .A1(n_422), .A2(n_1388), .B(n_1389), .Y(n_1387) );
AOI21xp5_ASAP7_75t_L g1404 ( .A1(n_422), .A2(n_1405), .B(n_1408), .Y(n_1404) );
INVxp67_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_425), .A2(n_444), .B1(n_763), .B2(n_764), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g1347 ( .A1(n_425), .A2(n_444), .B1(n_1348), .B2(n_1349), .Y(n_1347) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI22xp5_ASAP7_75t_L g558 ( .A1(n_426), .A2(n_444), .B1(n_559), .B2(n_560), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_426), .A2(n_444), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_426), .A2(n_444), .B1(n_666), .B2(n_667), .Y(n_665) );
INVx1_ASAP7_75t_L g736 ( .A(n_426), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_426), .A2(n_444), .B1(n_849), .B2(n_850), .Y(n_848) );
HB1xp67_ASAP7_75t_L g909 ( .A(n_426), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_426), .A2(n_732), .B1(n_1195), .B2(n_1196), .Y(n_1199) );
AOI22xp33_ASAP7_75t_L g1390 ( .A1(n_426), .A2(n_444), .B1(n_1391), .B2(n_1392), .Y(n_1390) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_426), .A2(n_445), .B1(n_1410), .B2(n_1411), .Y(n_1409) );
BUFx6f_ASAP7_75t_L g551 ( .A(n_427), .Y(n_551) );
INVx2_ASAP7_75t_L g574 ( .A(n_427), .Y(n_574) );
INVx1_ASAP7_75t_L g1407 ( .A(n_427), .Y(n_1407) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g775 ( .A(n_429), .Y(n_775) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g626 ( .A(n_431), .Y(n_626) );
INVx1_ASAP7_75t_L g1003 ( .A(n_431), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_431), .B(n_1125), .Y(n_1128) );
INVx1_ASAP7_75t_L g938 ( .A(n_432), .Y(n_938) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_434), .A2(n_479), .B1(n_483), .B2(n_484), .Y(n_478) );
INVx1_ASAP7_75t_L g1008 ( .A(n_435), .Y(n_1008) );
INVx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g575 ( .A(n_440), .Y(n_575) );
INVx2_ASAP7_75t_L g624 ( .A(n_440), .Y(n_624) );
OAI221xp5_ASAP7_75t_L g1208 ( .A1(n_440), .A2(n_995), .B1(n_1209), .B2(n_1210), .C(n_1213), .Y(n_1208) );
INVx1_ASAP7_75t_L g1416 ( .A(n_440), .Y(n_1416) );
INVxp67_ASAP7_75t_L g1117 ( .A(n_441), .Y(n_1117) );
INVx1_ASAP7_75t_L g1125 ( .A(n_441), .Y(n_1125) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g1282 ( .A1(n_444), .A2(n_447), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g733 ( .A(n_445), .Y(n_733) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_445), .B(n_961), .Y(n_1031) );
INVx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_SL g842 ( .A(n_447), .Y(n_842) );
NAND2xp5_ASAP7_75t_R g1206 ( .A(n_447), .B(n_1186), .Y(n_1206) );
BUFx2_ASAP7_75t_L g677 ( .A(n_448), .Y(n_677) );
INVx1_ASAP7_75t_L g1358 ( .A(n_448), .Y(n_1358) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g549 ( .A(n_449), .Y(n_549) );
BUFx3_ASAP7_75t_L g557 ( .A(n_449), .Y(n_557) );
BUFx3_ASAP7_75t_L g617 ( .A(n_449), .Y(n_617) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_450), .A2(n_761), .B(n_772), .Y(n_760) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g577 ( .A(n_451), .Y(n_577) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
OR2x2_ASAP7_75t_L g594 ( .A(n_452), .B(n_595), .Y(n_594) );
OR2x6_ASAP7_75t_L g953 ( .A(n_452), .B(n_595), .Y(n_953) );
AND2x4_ASAP7_75t_L g1012 ( .A(n_452), .B(n_1013), .Y(n_1012) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g603 ( .A(n_453), .Y(n_603) );
AOI21xp5_ASAP7_75t_SL g454 ( .A1(n_455), .A2(n_465), .B(n_466), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g836 ( .A1(n_455), .A2(n_837), .B(n_838), .Y(n_836) );
AOI21xp5_ASAP7_75t_L g1339 ( .A1(n_455), .A2(n_1340), .B(n_1341), .Y(n_1339) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g913 ( .A(n_456), .Y(n_913) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
AND2x4_ASAP7_75t_L g514 ( .A(n_457), .B(n_461), .Y(n_514) );
INVx2_ASAP7_75t_SL g1269 ( .A(n_457), .Y(n_1269) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g965 ( .A(n_461), .Y(n_965) );
INVx3_ASAP7_75t_L g485 ( .A(n_462), .Y(n_485) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx2_ASAP7_75t_L g1058 ( .A(n_463), .Y(n_1058) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_464), .Y(n_1102) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_470), .Y(n_598) );
INVx2_ASAP7_75t_L g795 ( .A(n_470), .Y(n_795) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_470), .Y(n_949) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_470), .B(n_1089), .Y(n_1105) );
INVx2_ASAP7_75t_L g1379 ( .A(n_470), .Y(n_1379) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_471), .Y(n_495) );
BUFx8_ASAP7_75t_L g505 ( .A(n_471), .Y(n_505) );
INVx2_ASAP7_75t_L g534 ( .A(n_471), .Y(n_534) );
INVx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx3_ASAP7_75t_L g878 ( .A(n_474), .Y(n_878) );
CKINVDCx8_ASAP7_75t_R g1381 ( .A(n_474), .Y(n_1381) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_476), .Y(n_518) );
BUFx8_ASAP7_75t_L g876 ( .A(n_476), .Y(n_876) );
BUFx4f_ASAP7_75t_L g1369 ( .A(n_476), .Y(n_1369) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_477), .Y(n_1040) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
BUFx4f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g715 ( .A(n_482), .Y(n_715) );
OR2x4_ASAP7_75t_L g1088 ( .A(n_482), .B(n_1089), .Y(n_1088) );
OAI22xp33_ASAP7_75t_L g877 ( .A1(n_484), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_877) );
OAI22xp33_ASAP7_75t_L g890 ( .A1(n_484), .A2(n_882), .B1(n_891), .B2(n_892), .Y(n_890) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx3_ASAP7_75t_L g1249 ( .A(n_485), .Y(n_1249) );
OAI33xp33_ASAP7_75t_L g875 ( .A1(n_486), .A2(n_876), .A3(n_877), .B1(n_881), .B2(n_886), .B3(n_890), .Y(n_875) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g650 ( .A(n_487), .B(n_651), .C(n_654), .Y(n_650) );
AOI33xp33_ASAP7_75t_L g790 ( .A1(n_487), .A2(n_601), .A3(n_791), .B1(n_793), .B2(n_797), .B3(n_798), .Y(n_790) );
BUFx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g710 ( .A(n_488), .Y(n_710) );
BUFx2_ASAP7_75t_L g830 ( .A(n_488), .Y(n_830) );
BUFx2_ASAP7_75t_L g1191 ( .A(n_488), .Y(n_1191) );
INVx3_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g881 ( .A1(n_493), .A2(n_882), .B1(n_884), .B2(n_885), .Y(n_881) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx8_ASAP7_75t_L g709 ( .A(n_494), .Y(n_709) );
INVx5_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g521 ( .A(n_495), .Y(n_521) );
INVx2_ASAP7_75t_SL g825 ( .A(n_495), .Y(n_825) );
INVx3_ASAP7_75t_L g1039 ( .A(n_495), .Y(n_1039) );
HB1xp67_ASAP7_75t_L g1311 ( .A(n_495), .Y(n_1311) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_497), .A2(n_532), .B1(n_535), .B2(n_536), .C(n_537), .Y(n_531) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g1374 ( .A(n_498), .Y(n_1374) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g538 ( .A(n_502), .Y(n_538) );
INVx1_ASAP7_75t_L g801 ( .A(n_502), .Y(n_801) );
INVx2_ASAP7_75t_L g951 ( .A(n_502), .Y(n_951) );
INVxp67_ASAP7_75t_L g579 ( .A(n_503), .Y(n_579) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g789 ( .A(n_504), .Y(n_789) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_505), .Y(n_641) );
INVx2_ASAP7_75t_SL g887 ( .A(n_505), .Y(n_887) );
INVx3_ASAP7_75t_L g1336 ( .A(n_505), .Y(n_1336) );
INVx2_ASAP7_75t_SL g1422 ( .A(n_505), .Y(n_1422) );
INVx1_ASAP7_75t_L g632 ( .A(n_507), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g507 ( .A(n_508), .B(n_580), .Y(n_507) );
NAND4xp75_ASAP7_75t_L g509 ( .A(n_510), .B(n_516), .C(n_544), .D(n_578), .Y(n_509) );
INVx1_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_529), .B2(n_531), .Y(n_517) );
OAI211xp5_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_522), .C(n_525), .Y(n_519) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_R g1312 ( .A(n_527), .Y(n_1312) );
INVx1_ASAP7_75t_L g1333 ( .A(n_527), .Y(n_1333) );
INVx5_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
BUFx12f_ASAP7_75t_L g597 ( .A(n_528), .Y(n_597) );
BUFx3_ASAP7_75t_L g642 ( .A(n_528), .Y(n_642) );
BUFx3_ASAP7_75t_L g796 ( .A(n_528), .Y(n_796) );
BUFx2_ASAP7_75t_L g826 ( .A(n_528), .Y(n_826) );
AND2x4_ASAP7_75t_L g1065 ( .A(n_528), .B(n_1063), .Y(n_1065) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AOI33xp33_ASAP7_75t_L g1327 ( .A1(n_530), .A2(n_644), .A3(n_1328), .B1(n_1330), .B2(n_1334), .B3(n_1337), .Y(n_1327) );
INVx2_ASAP7_75t_L g1377 ( .A(n_530), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g1426 ( .A(n_530), .Y(n_1426) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g630 ( .A(n_533), .B(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g707 ( .A(n_534), .Y(n_707) );
INVx1_ASAP7_75t_L g1035 ( .A(n_534), .Y(n_1035) );
OR2x6_ASAP7_75t_SL g1061 ( .A(n_534), .B(n_1062), .Y(n_1061) );
BUFx2_ASAP7_75t_L g1332 ( .A(n_534), .Y(n_1332) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_534), .A2(n_1371), .B1(n_1372), .B2(n_1375), .C(n_1376), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_538), .B(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_543), .A2(n_588), .B1(n_589), .B2(n_590), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_561), .B(n_576), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
INVx2_ASAP7_75t_L g923 ( .A(n_547), .Y(n_923) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_548), .B(n_1020), .Y(n_1019) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g684 ( .A(n_549), .Y(n_684) );
BUFx3_ASAP7_75t_L g1203 ( .A(n_551), .Y(n_1203) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_SL g683 ( .A(n_555), .Y(n_683) );
INVx1_ASAP7_75t_L g1148 ( .A(n_555), .Y(n_1148) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_556), .Y(n_847) );
OAI221xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B1(n_565), .B2(n_567), .C(n_568), .Y(n_562) );
BUFx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g1130 ( .A(n_569), .B(n_1100), .Y(n_1130) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_571), .B(n_1125), .Y(n_1132) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx2_ASAP7_75t_L g674 ( .A(n_572), .Y(n_674) );
INVx1_ASAP7_75t_L g727 ( .A(n_573), .Y(n_727) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g681 ( .A(n_574), .Y(n_681) );
OAI21xp33_ASAP7_75t_L g1342 ( .A1(n_576), .A2(n_1343), .B(n_1350), .Y(n_1342) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g606 ( .A(n_577), .Y(n_606) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_605), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_584), .B(n_695), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_584), .A2(n_719), .B(n_720), .Y(n_718) );
AOI21xp33_ASAP7_75t_L g756 ( .A1(n_584), .A2(n_757), .B(n_758), .Y(n_756) );
NAND2xp33_ASAP7_75t_L g831 ( .A(n_584), .B(n_832), .Y(n_831) );
AOI21xp33_ASAP7_75t_L g910 ( .A1(n_584), .A2(n_911), .B(n_912), .Y(n_910) );
AOI211x1_ASAP7_75t_L g1177 ( .A1(n_584), .A2(n_1178), .B(n_1179), .C(n_1193), .Y(n_1177) );
AOI21xp33_ASAP7_75t_SL g1300 ( .A1(n_584), .A2(n_1301), .B(n_1302), .Y(n_1300) );
AOI211x1_ASAP7_75t_L g1319 ( .A1(n_584), .A2(n_1320), .B(n_1321), .C(n_1338), .Y(n_1319) );
AOI21xp5_ASAP7_75t_L g1364 ( .A1(n_584), .A2(n_1365), .B(n_1366), .Y(n_1364) );
AOI21xp5_ASAP7_75t_L g1431 ( .A1(n_584), .A2(n_1432), .B(n_1433), .Y(n_1431) );
AOI222xp33_ASAP7_75t_L g618 ( .A1(n_588), .A2(n_590), .B1(n_619), .B2(n_620), .C1(n_622), .C2(n_625), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B1(n_599), .B2(n_604), .Y(n_591) );
INVx1_ASAP7_75t_L g653 ( .A(n_593), .Y(n_653) );
INVx3_ASAP7_75t_L g1244 ( .A(n_595), .Y(n_1244) );
BUFx2_ASAP7_75t_L g655 ( .A(n_597), .Y(n_655) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx3_ASAP7_75t_L g644 ( .A(n_601), .Y(n_644) );
AOI33xp33_ASAP7_75t_L g820 ( .A1(n_601), .A2(n_821), .A3(n_823), .B1(n_827), .B2(n_828), .B3(n_830), .Y(n_820) );
AOI33xp33_ASAP7_75t_L g944 ( .A1(n_601), .A2(n_945), .A3(n_947), .B1(n_948), .B2(n_950), .B3(n_952), .Y(n_944) );
AOI33xp33_ASAP7_75t_L g1308 ( .A1(n_601), .A2(n_710), .A3(n_1309), .B1(n_1310), .B2(n_1313), .B3(n_1314), .Y(n_1308) );
INVx3_ASAP7_75t_L g1098 ( .A(n_602), .Y(n_1098) );
INVx2_ASAP7_75t_SL g691 ( .A(n_603), .Y(n_691) );
INVx1_ASAP7_75t_L g749 ( .A(n_603), .Y(n_749) );
OAI31xp33_ASAP7_75t_SL g1230 ( .A1(n_603), .A2(n_1231), .A3(n_1232), .B(n_1236), .Y(n_1230) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_607), .B(n_627), .Y(n_605) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_606), .A2(n_841), .B(n_851), .Y(n_840) );
OAI21xp5_ASAP7_75t_L g1197 ( .A1(n_606), .A2(n_1198), .B(n_1207), .Y(n_1197) );
OAI21xp5_ASAP7_75t_L g1385 ( .A1(n_606), .A2(n_1386), .B(n_1393), .Y(n_1385) );
NAND3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .C(n_618), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_609), .A2(n_610), .B1(n_629), .B2(n_630), .Y(n_628) );
BUFx2_ASAP7_75t_L g725 ( .A(n_613), .Y(n_725) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g621 ( .A(n_616), .Y(n_621) );
INVx2_ASAP7_75t_SL g676 ( .A(n_616), .Y(n_676) );
INVx2_ASAP7_75t_L g771 ( .A(n_616), .Y(n_771) );
INVx1_ASAP7_75t_L g903 ( .A(n_616), .Y(n_903) );
INVx2_ASAP7_75t_L g1205 ( .A(n_616), .Y(n_1205) );
BUFx3_ASAP7_75t_L g729 ( .A(n_617), .Y(n_729) );
INVx1_ASAP7_75t_SL g905 ( .A(n_617), .Y(n_905) );
INVx1_ASAP7_75t_L g689 ( .A(n_619), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_625), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_626), .A2(n_934), .B1(n_935), .B2(n_937), .Y(n_933) );
AOI222xp33_ASAP7_75t_L g964 ( .A1(n_629), .A2(n_937), .B1(n_965), .B2(n_966), .C1(n_967), .C2(n_968), .Y(n_964) );
INVx2_ASAP7_75t_SL g958 ( .A(n_630), .Y(n_958) );
INVxp67_ASAP7_75t_L g716 ( .A(n_631), .Y(n_716) );
OAI22x1_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_696), .B2(n_750), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
AND3x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_663), .C(n_694), .Y(n_637) );
NOR2xp33_ASAP7_75t_SL g638 ( .A(n_639), .B(n_656), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_640), .A2(n_643), .B(n_650), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
AOI33xp33_ASAP7_75t_L g703 ( .A1(n_644), .A2(n_704), .A3(n_705), .B1(n_708), .B2(n_710), .B3(n_711), .Y(n_703) );
AOI33xp33_ASAP7_75t_L g1187 ( .A1(n_644), .A2(n_1188), .A3(n_1189), .B1(n_1190), .B2(n_1191), .B3(n_1192), .Y(n_1187) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g1081 ( .A1(n_647), .A2(n_952), .B1(n_1082), .B2(n_1083), .C(n_1084), .Y(n_1081) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NAND3xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .C(n_660), .Y(n_656) );
NAND4xp25_ASAP7_75t_SL g811 ( .A(n_657), .B(n_812), .C(n_817), .D(n_820), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g1184 ( .A(n_657), .B(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1316 ( .A(n_657), .Y(n_1316) );
NAND4xp25_ASAP7_75t_SL g1321 ( .A(n_657), .B(n_1322), .C(n_1325), .D(n_1327), .Y(n_1321) );
AOI21xp5_ASAP7_75t_SL g663 ( .A1(n_664), .A2(n_691), .B(n_692), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .C(n_678), .Y(n_664) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_672), .Y(n_741) );
INVx1_ASAP7_75t_L g768 ( .A(n_672), .Y(n_768) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g1202 ( .A(n_674), .Y(n_1202) );
AOI31xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .A3(n_685), .B(n_688), .Y(n_678) );
BUFx2_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g785 ( .A(n_687), .Y(n_785) );
INVx1_ASAP7_75t_L g750 ( .A(n_696), .Y(n_750) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_698), .B(n_718), .C(n_721), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_712), .C(n_717), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_703), .Y(n_699) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x6_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
OR2x2_ASAP7_75t_L g839 ( .A(n_714), .B(n_716), .Y(n_839) );
INVx2_ASAP7_75t_SL g883 ( .A(n_714), .Y(n_883) );
INVx2_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g1367 ( .A(n_717), .B(n_1368), .C(n_1384), .Y(n_1367) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_737), .B(n_746), .Y(n_721) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_734), .B2(n_735), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_732), .A2(n_907), .B1(n_908), .B2(n_909), .Y(n_906) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx5_ASAP7_75t_L g1219 ( .A(n_738), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
INVxp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g1123 ( .A(n_744), .B(n_1120), .Y(n_1123) );
OR2x6_ASAP7_75t_L g1155 ( .A(n_744), .B(n_1117), .Y(n_1155) );
OAI21xp5_ASAP7_75t_L g894 ( .A1(n_746), .A2(n_895), .B(n_898), .Y(n_894) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g1032 ( .A1(n_748), .A2(n_1033), .B(n_1048), .C(n_1066), .Y(n_1032) );
INVx1_ASAP7_75t_L g1299 ( .A(n_748), .Y(n_1299) );
BUFx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AOI21x1_ASAP7_75t_L g921 ( .A1(n_749), .A2(n_922), .B(n_942), .Y(n_921) );
BUFx2_ASAP7_75t_L g1418 ( .A(n_749), .Y(n_1418) );
XNOR2x1_ASAP7_75t_L g751 ( .A(n_752), .B(n_867), .Y(n_751) );
OAI22x1_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_806), .B1(n_807), .B2(n_866), .Y(n_752) );
INVx2_ASAP7_75t_L g866 ( .A(n_753), .Y(n_866) );
AO21x2_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_755), .B(n_805), .Y(n_753) );
NAND3xp33_ASAP7_75t_SL g755 ( .A(n_756), .B(n_760), .C(n_786), .Y(n_755) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
BUFx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_779), .B1(n_780), .B2(n_783), .C(n_784), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g988 ( .A(n_781), .Y(n_988) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
NAND2x1p5_ASAP7_75t_L g807 ( .A(n_808), .B(n_833), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_831), .Y(n_809) );
INVxp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NOR2xp33_ASAP7_75t_SL g863 ( .A(n_811), .B(n_864), .Y(n_863) );
INVx2_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g1185 ( .A(n_819), .B(n_1186), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_819), .B(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1082 ( .A(n_822), .Y(n_1082) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_831), .B(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_840), .Y(n_835) );
INVx1_ASAP7_75t_L g861 ( .A(n_845), .Y(n_861) );
OAI211xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B(n_859), .C(n_862), .Y(n_853) );
INVx2_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g1395 ( .A(n_856), .Y(n_1395) );
INVx4_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
BUFx4f_ASAP7_75t_L g941 ( .A(n_857), .Y(n_941) );
BUFx4f_ASAP7_75t_L g995 ( .A(n_857), .Y(n_995) );
OR2x6_ASAP7_75t_L g1005 ( .A(n_857), .B(n_1006), .Y(n_1005) );
BUFx4f_ASAP7_75t_L g1288 ( .A(n_857), .Y(n_1288) );
BUFx6f_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx3_ASAP7_75t_L g1025 ( .A(n_858), .Y(n_1025) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
AND3x2_ASAP7_75t_L g869 ( .A(n_870), .B(n_894), .C(n_910), .Y(n_869) );
NOR4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_874), .C(n_875), .D(n_893), .Y(n_870) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_SL g1420 ( .A1(n_876), .A2(n_1421), .B1(n_1426), .B2(n_1427), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_878), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
CKINVDCx14_ASAP7_75t_R g977 ( .A(n_915), .Y(n_977) );
CKINVDCx6p67_ASAP7_75t_R g915 ( .A(n_916), .Y(n_915) );
HB1xp67_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
HB1xp67_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
NAND3xp33_ASAP7_75t_L g919 ( .A(n_920), .B(n_969), .C(n_973), .Y(n_919) );
INVx1_ASAP7_75t_L g970 ( .A(n_921), .Y(n_970) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_925), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_924) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_938), .B1(n_939), .B2(n_940), .Y(n_929) );
INVx3_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
BUFx6f_ASAP7_75t_L g1217 ( .A(n_932), .Y(n_1217) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
INVx1_ASAP7_75t_L g971 ( .A(n_943), .Y(n_971) );
AND2x2_ASAP7_75t_L g943 ( .A(n_944), .B(n_954), .Y(n_943) );
BUFx2_ASAP7_75t_L g1329 ( .A(n_946), .Y(n_1329) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g975 ( .A(n_956), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_957), .B(n_963), .Y(n_956) );
NAND2x1_ASAP7_75t_L g957 ( .A(n_958), .B(n_959), .Y(n_957) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_960), .B(n_1067), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_960), .B(n_1229), .Y(n_1228) );
AND2x4_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
INVx1_ASAP7_75t_L g974 ( .A(n_964), .Y(n_974) );
OAI21xp5_ASAP7_75t_L g969 ( .A1(n_970), .A2(n_971), .B(n_972), .Y(n_969) );
OAI21xp33_ASAP7_75t_L g973 ( .A1(n_972), .A2(n_974), .B(n_975), .Y(n_973) );
NOR3xp33_ASAP7_75t_SL g978 ( .A(n_979), .B(n_1171), .C(n_1436), .Y(n_978) );
NOR3xp33_ASAP7_75t_L g1647 ( .A(n_979), .B(n_1436), .C(n_1648), .Y(n_1647) );
NOR3xp33_ASAP7_75t_L g1649 ( .A(n_979), .B(n_1436), .C(n_1650), .Y(n_1649) );
OAI222xp33_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_1068), .B1(n_1075), .B2(n_1150), .C1(n_1152), .C2(n_1160), .Y(n_979) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
HB1xp67_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
OR2x2_ASAP7_75t_L g984 ( .A(n_985), .B(n_1032), .Y(n_984) );
NAND3xp33_ASAP7_75t_SL g985 ( .A(n_986), .B(n_1014), .C(n_1027), .Y(n_985) );
AOI211xp5_ASAP7_75t_SL g986 ( .A1(n_987), .A2(n_990), .B(n_998), .C(n_1007), .Y(n_986) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_992), .A2(n_995), .B1(n_1010), .B2(n_1011), .C(n_1012), .Y(n_1009) );
BUFx3_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
BUFx2_ASAP7_75t_L g1212 ( .A(n_993), .Y(n_1212) );
INVxp67_ASAP7_75t_SL g994 ( .A(n_995), .Y(n_994) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
AOI33xp33_ASAP7_75t_L g1141 ( .A1(n_997), .A2(n_1142), .A3(n_1144), .B1(n_1145), .B2(n_1146), .B3(n_1147), .Y(n_1141) );
INVx1_ASAP7_75t_L g1268 ( .A(n_999), .Y(n_1268) );
NAND2x2_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1002), .Y(n_999) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1000), .Y(n_1006) );
INVx2_ASAP7_75t_L g1000 ( .A(n_1001), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1002 ( .A(n_1003), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_1005), .Y(n_1272) );
INVx4_ASAP7_75t_L g1143 ( .A(n_1012), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1259 ( .A(n_1012), .Y(n_1259) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_1015), .A2(n_1018), .B1(n_1019), .B2(n_1022), .C1(n_1023), .C2(n_1026), .Y(n_1014) );
AOI21xp33_ASAP7_75t_SL g1270 ( .A1(n_1015), .A2(n_1271), .B(n_1272), .Y(n_1270) );
AND2x4_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
AOI222xp33_ASAP7_75t_L g1266 ( .A1(n_1019), .A2(n_1234), .B1(n_1246), .B2(n_1267), .C1(n_1268), .C2(n_1269), .Y(n_1266) );
INVx1_ASAP7_75t_L g1020 ( .A(n_1021), .Y(n_1020) );
OR2x2_ASAP7_75t_L g1024 ( .A(n_1021), .B(n_1025), .Y(n_1024) );
AOI211xp5_ASAP7_75t_L g1048 ( .A1(n_1022), .A2(n_1049), .B(n_1052), .C(n_1060), .Y(n_1048) );
AOI222xp33_ASAP7_75t_L g1253 ( .A1(n_1023), .A2(n_1235), .B1(n_1254), .B2(n_1259), .C1(n_1260), .C2(n_1263), .Y(n_1253) );
INVx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_SL g1354 ( .A(n_1025), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1029), .Y(n_1027) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx3_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1031), .Y(n_1225) );
AOI221xp5_ASAP7_75t_L g1033 ( .A1(n_1034), .A2(n_1036), .B1(n_1037), .B2(n_1041), .C(n_1042), .Y(n_1033) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
OAI221xp5_ASAP7_75t_L g1237 ( .A1(n_1039), .A2(n_1238), .B1(n_1239), .B2(n_1240), .C(n_1241), .Y(n_1237) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AOI22xp5_ASAP7_75t_L g1245 ( .A1(n_1044), .A2(n_1047), .B1(n_1226), .B2(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
INVx4_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_1054), .A2(n_1056), .B1(n_1234), .B2(n_1235), .Y(n_1233) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
OR2x6_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1059), .Y(n_1057) );
INVx2_ASAP7_75t_L g1062 ( .A(n_1063), .Y(n_1062) );
INVx3_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
INVx1_ASAP7_75t_L g1068 ( .A(n_1069), .Y(n_1068) );
HB1xp67_ASAP7_75t_L g1069 ( .A(n_1070), .Y(n_1069) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NOR2xp33_ASAP7_75t_L g1071 ( .A(n_1072), .B(n_1073), .Y(n_1071) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1072), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1072), .B(n_1164), .Y(n_1170) );
NOR2xp33_ASAP7_75t_L g1158 ( .A(n_1073), .B(n_1159), .Y(n_1158) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1073), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
OR2x2_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1137), .Y(n_1075) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1077), .Y(n_1139) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1079), .B(n_1080), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_1085), .B(n_1112), .Y(n_1138) );
OAI31xp33_ASAP7_75t_SL g1085 ( .A1(n_1086), .A2(n_1090), .A3(n_1103), .B(n_1107), .Y(n_1085) );
NAND3xp33_ASAP7_75t_SL g1090 ( .A(n_1091), .B(n_1093), .C(n_1095), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_1092), .A2(n_1096), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
CKINVDCx8_ASAP7_75t_R g1093 ( .A(n_1094), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_1096), .A2(n_1097), .B1(n_1100), .B2(n_1101), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1099), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1098), .B(n_1102), .Y(n_1101) );
INVx2_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1110), .Y(n_1107) );
INVx1_ASAP7_75t_SL g1108 ( .A(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
AO21x1_ASAP7_75t_L g1112 ( .A1(n_1113), .A2(n_1121), .B(n_1133), .Y(n_1112) );
AOI22xp5_ASAP7_75t_L g1113 ( .A1(n_1114), .A2(n_1115), .B1(n_1118), .B2(n_1119), .Y(n_1113) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
NOR2xp33_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1126), .Y(n_1121) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1130), .C(n_1131), .Y(n_1126) );
INVx2_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
AND2x4_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1136), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g1156 ( .A(n_1135), .B(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1135), .Y(n_1654) );
OAI31xp33_ASAP7_75t_L g1137 ( .A1(n_1138), .A2(n_1139), .A3(n_1140), .B(n_1149), .Y(n_1137) );
INVx1_ASAP7_75t_L g1151 ( .A(n_1141), .Y(n_1151) );
INVx2_ASAP7_75t_SL g1142 ( .A(n_1143), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1151), .Y(n_1149) );
INVx2_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
AND2x4_ASAP7_75t_SL g1153 ( .A(n_1154), .B(n_1156), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1653 ( .A(n_1154), .B(n_1654), .Y(n_1653) );
INVx3_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
OR2x2_ASAP7_75t_L g1651 ( .A(n_1157), .B(n_1652), .Y(n_1651) );
INVx1_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
HB1xp67_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
OAI21xp5_ASAP7_75t_L g1163 ( .A1(n_1164), .A2(n_1165), .B(n_1169), .Y(n_1163) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1438 ( .A(n_1166), .B(n_1439), .Y(n_1438) );
AND2x4_ASAP7_75t_L g1450 ( .A(n_1166), .B(n_1439), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1168), .Y(n_1166) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1171), .Y(n_1648) );
XNOR2xp5_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1360), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1174), .B1(n_1274), .B2(n_1359), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
AOI22xp5_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1221), .B1(n_1222), .B2(n_1273), .Y(n_1174) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1175), .Y(n_1273) );
XOR2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1220), .Y(n_1175) );
NAND2xp5_ASAP7_75t_SL g1176 ( .A(n_1177), .B(n_1197), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1187), .Y(n_1179) );
NOR2xp33_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1184), .Y(n_1180) );
NAND3xp33_ASAP7_75t_SL g1198 ( .A(n_1199), .B(n_1200), .C(n_1206), .Y(n_1198) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx4_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
OAI22xp5_ASAP7_75t_L g1214 ( .A1(n_1215), .A2(n_1216), .B1(n_1218), .B2(n_1219), .Y(n_1214) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
AOI211x1_ASAP7_75t_L g1224 ( .A1(n_1225), .A2(n_1226), .B(n_1227), .C(n_1252), .Y(n_1224) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1230), .Y(n_1227) );
NAND3xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1245), .C(n_1247), .Y(n_1236) );
INVx3_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
OAI211xp5_ASAP7_75t_L g1247 ( .A1(n_1248), .A2(n_1249), .B(n_1250), .C(n_1251), .Y(n_1247) );
NAND3xp33_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1266), .C(n_1270), .Y(n_1252) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx2_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
HB1xp67_ASAP7_75t_L g1359 ( .A(n_1275), .Y(n_1359) );
XNOR2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1317), .Y(n_1275) );
NAND3xp33_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1300), .C(n_1303), .Y(n_1277) );
OAI31xp33_ASAP7_75t_L g1278 ( .A1(n_1279), .A2(n_1285), .A3(n_1297), .B(n_1298), .Y(n_1278) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1282), .Y(n_1279) );
OAI211xp5_ASAP7_75t_L g1286 ( .A1(n_1287), .A2(n_1288), .B(n_1289), .C(n_1290), .Y(n_1286) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
NOR3xp33_ASAP7_75t_L g1303 ( .A(n_1304), .B(n_1315), .C(n_1316), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1308), .Y(n_1304) );
XNOR2x2_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1338 ( .A(n_1339), .B(n_1342), .Y(n_1338) );
OAI211xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1353), .B(n_1355), .C(n_1356), .Y(n_1351) );
OAI211xp5_ASAP7_75t_L g1413 ( .A1(n_1353), .A2(n_1414), .B(n_1415), .C(n_1417), .Y(n_1413) );
INVx5_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
HB1xp67_ASAP7_75t_L g1360 ( .A(n_1361), .Y(n_1360) );
AO22x2_ASAP7_75t_L g1361 ( .A1(n_1362), .A2(n_1399), .B1(n_1400), .B2(n_1435), .Y(n_1361) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1362), .Y(n_1435) );
AND4x1_ASAP7_75t_L g1363 ( .A(n_1364), .B(n_1367), .C(n_1385), .D(n_1398), .Y(n_1363) );
OAI22xp5_ASAP7_75t_SL g1368 ( .A1(n_1369), .A2(n_1370), .B1(n_1377), .B2(n_1378), .Y(n_1368) );
OAI221xp5_ASAP7_75t_L g1421 ( .A1(n_1372), .A2(n_1422), .B1(n_1423), .B2(n_1424), .C(n_1425), .Y(n_1421) );
INVx3_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
BUFx2_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
OAI221xp5_ASAP7_75t_L g1378 ( .A1(n_1379), .A2(n_1380), .B1(n_1381), .B2(n_1382), .C(n_1383), .Y(n_1378) );
OAI211xp5_ASAP7_75t_L g1394 ( .A1(n_1380), .A2(n_1395), .B(n_1396), .C(n_1397), .Y(n_1394) );
OAI221xp5_ASAP7_75t_L g1427 ( .A1(n_1381), .A2(n_1414), .B1(n_1422), .B2(n_1428), .C(n_1429), .Y(n_1427) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
AND4x1_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1419), .C(n_1431), .D(n_1434), .Y(n_1401) );
OAI21xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1412), .B(n_1418), .Y(n_1402) );
INVx2_ASAP7_75t_SL g1406 ( .A(n_1407), .Y(n_1406) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1437), .B(n_1440), .Y(n_1436) );
BUFx2_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AND2x6_ASAP7_75t_L g1445 ( .A(n_1439), .B(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1439), .B(n_1448), .Y(n_1447) );
AND2x6_ASAP7_75t_L g1451 ( .A(n_1439), .B(n_1452), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1458 ( .A(n_1439), .B(n_1448), .Y(n_1458) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1439), .B(n_1448), .Y(n_1468) );
AOI21xp5_ASAP7_75t_L g1440 ( .A1(n_1441), .A2(n_1559), .B(n_1603), .Y(n_1440) );
OAI211xp5_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1453), .B(n_1499), .C(n_1545), .Y(n_1441) );
AOI22xp5_ASAP7_75t_L g1628 ( .A1(n_1442), .A2(n_1551), .B1(n_1629), .B2(n_1635), .Y(n_1628) );
CKINVDCx5p33_ASAP7_75t_R g1442 ( .A(n_1443), .Y(n_1442) );
CKINVDCx6p67_ASAP7_75t_R g1511 ( .A(n_1443), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1612 ( .A(n_1443), .B(n_1471), .Y(n_1612) );
OR2x2_ASAP7_75t_L g1630 ( .A(n_1443), .B(n_1471), .Y(n_1630) );
OR2x2_ASAP7_75t_L g1645 ( .A(n_1443), .B(n_1535), .Y(n_1645) );
OR2x6_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1449), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1532 ( .A(n_1444), .B(n_1449), .Y(n_1532) );
INVx2_ASAP7_75t_L g1542 ( .A(n_1445), .Y(n_1542) );
O2A1O1Ixp33_ASAP7_75t_L g1453 ( .A1(n_1454), .A2(n_1469), .B(n_1474), .C(n_1488), .Y(n_1453) );
NOR2xp33_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1459), .Y(n_1454) );
INVx2_ASAP7_75t_L g1482 ( .A(n_1455), .Y(n_1482) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1455), .B(n_1490), .Y(n_1489) );
AND2x2_ASAP7_75t_L g1496 ( .A(n_1455), .B(n_1464), .Y(n_1496) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1455), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1455), .B(n_1527), .Y(n_1526) );
OR2x2_ASAP7_75t_L g1569 ( .A(n_1455), .B(n_1531), .Y(n_1569) );
AND2x2_ASAP7_75t_L g1601 ( .A(n_1455), .B(n_1484), .Y(n_1601) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1455), .B(n_1484), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
INVxp67_ASAP7_75t_L g1544 ( .A(n_1458), .Y(n_1544) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1464), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1460), .B(n_1493), .Y(n_1498) );
AND3x1_ASAP7_75t_L g1515 ( .A(n_1460), .B(n_1476), .C(n_1481), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1522 ( .A(n_1460), .B(n_1476), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1460), .B(n_1464), .Y(n_1634) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1461), .B(n_1476), .Y(n_1475) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_1461), .B(n_1493), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1531 ( .A(n_1461), .B(n_1464), .Y(n_1531) );
OR2x2_ASAP7_75t_L g1461 ( .A(n_1462), .B(n_1463), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1492 ( .A(n_1464), .B(n_1493), .Y(n_1492) );
OR2x2_ASAP7_75t_L g1517 ( .A(n_1464), .B(n_1476), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1584 ( .A(n_1464), .B(n_1522), .Y(n_1584) );
AND2x2_ASAP7_75t_L g1599 ( .A(n_1464), .B(n_1476), .Y(n_1599) );
BUFx2_ASAP7_75t_L g1464 ( .A(n_1465), .Y(n_1464) );
INVx2_ASAP7_75t_L g1481 ( .A(n_1465), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1513 ( .A(n_1465), .B(n_1475), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1534 ( .A(n_1465), .B(n_1498), .Y(n_1534) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1465), .B(n_1506), .Y(n_1566) );
OR2x2_ASAP7_75t_L g1587 ( .A(n_1465), .B(n_1588), .Y(n_1587) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1466), .B(n_1467), .Y(n_1465) );
O2A1O1Ixp33_ASAP7_75t_L g1474 ( .A1(n_1469), .A2(n_1475), .B(n_1479), .C(n_1483), .Y(n_1474) );
CKINVDCx14_ASAP7_75t_R g1469 ( .A(n_1470), .Y(n_1469) );
OAI22xp5_ASAP7_75t_L g1552 ( .A1(n_1470), .A2(n_1550), .B1(n_1553), .B2(n_1556), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1470), .B(n_1538), .Y(n_1570) );
AOI211xp5_ASAP7_75t_L g1594 ( .A1(n_1470), .A2(n_1595), .B(n_1596), .C(n_1597), .Y(n_1594) );
AOI221xp5_ASAP7_75t_L g1604 ( .A1(n_1470), .A2(n_1515), .B1(n_1605), .B2(n_1607), .C(n_1608), .Y(n_1604) );
INVx3_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1471), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1501 ( .A(n_1471), .B(n_1484), .Y(n_1501) );
AOI22xp5_ASAP7_75t_L g1525 ( .A1(n_1471), .A2(n_1526), .B1(n_1529), .B2(n_1530), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1529 ( .A(n_1471), .B(n_1484), .Y(n_1529) );
AND2x2_ASAP7_75t_L g1536 ( .A(n_1471), .B(n_1490), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1582 ( .A(n_1471), .B(n_1511), .Y(n_1582) );
AND2x2_ASAP7_75t_L g1600 ( .A(n_1471), .B(n_1601), .Y(n_1600) );
AND2x2_ASAP7_75t_L g1627 ( .A(n_1471), .B(n_1511), .Y(n_1627) );
AND2x4_ASAP7_75t_L g1471 ( .A(n_1472), .B(n_1473), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1549 ( .A(n_1475), .B(n_1482), .Y(n_1549) );
INVx1_ASAP7_75t_L g1588 ( .A(n_1475), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1632 ( .A(n_1475), .B(n_1496), .Y(n_1632) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1476), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1528 ( .A(n_1476), .B(n_1481), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1478), .Y(n_1476) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1637 ( .A(n_1480), .B(n_1498), .Y(n_1637) );
AND2x2_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1482), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1481), .B(n_1506), .Y(n_1505) );
OR2x2_ASAP7_75t_L g1548 ( .A(n_1481), .B(n_1549), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1591 ( .A(n_1481), .B(n_1498), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1640 ( .A(n_1481), .B(n_1558), .Y(n_1640) );
NAND2xp5_ASAP7_75t_SL g1642 ( .A(n_1481), .B(n_1643), .Y(n_1642) );
NOR2xp33_ASAP7_75t_L g1520 ( .A(n_1482), .B(n_1521), .Y(n_1520) );
NOR2xp33_ASAP7_75t_L g1555 ( .A(n_1482), .B(n_1517), .Y(n_1555) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1482), .B(n_1510), .Y(n_1565) );
INVx1_ASAP7_75t_L g1593 ( .A(n_1482), .Y(n_1593) );
NAND2xp5_ASAP7_75t_L g1625 ( .A(n_1482), .B(n_1599), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1518 ( .A(n_1483), .B(n_1511), .Y(n_1518) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1483), .Y(n_1576) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1487), .Y(n_1483) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1484), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
OAI21xp33_ASAP7_75t_L g1488 ( .A1(n_1489), .A2(n_1491), .B(n_1494), .Y(n_1488) );
INVx2_ASAP7_75t_L g1510 ( .A(n_1490), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1523 ( .A(n_1490), .B(n_1511), .Y(n_1523) );
OAI211xp5_ASAP7_75t_SL g1561 ( .A1(n_1491), .A2(n_1562), .B(n_1563), .C(n_1567), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1586 ( .A(n_1491), .B(n_1587), .Y(n_1586) );
INVx1_ASAP7_75t_L g1491 ( .A(n_1492), .Y(n_1491) );
A2O1A1Ixp33_ASAP7_75t_L g1519 ( .A1(n_1492), .A2(n_1504), .B(n_1520), .C(n_1523), .Y(n_1519) );
AOI221xp5_ASAP7_75t_L g1545 ( .A1(n_1492), .A2(n_1546), .B1(n_1547), .B2(n_1550), .C(n_1552), .Y(n_1545) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1494), .Y(n_1595) );
OR2x2_ASAP7_75t_L g1622 ( .A(n_1494), .B(n_1510), .Y(n_1622) );
OR2x2_ASAP7_75t_L g1494 ( .A(n_1495), .B(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
NAND2xp5_ASAP7_75t_L g1558 ( .A(n_1498), .B(n_1504), .Y(n_1558) );
AOI211xp5_ASAP7_75t_L g1499 ( .A1(n_1500), .A2(n_1502), .B(n_1507), .C(n_1524), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1546 ( .A(n_1500), .B(n_1504), .Y(n_1546) );
OAI322xp33_ASAP7_75t_L g1573 ( .A1(n_1500), .A2(n_1517), .A3(n_1532), .B1(n_1549), .B2(n_1574), .C1(n_1577), .C2(n_1579), .Y(n_1573) );
AND2x2_ASAP7_75t_SL g1596 ( .A(n_1500), .B(n_1515), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1606 ( .A(n_1500), .B(n_1503), .Y(n_1606) );
INVx2_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1505), .Y(n_1502) );
NOR2xp33_ASAP7_75t_L g1516 ( .A(n_1503), .B(n_1517), .Y(n_1516) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1503), .Y(n_1578) );
AOI31xp33_ASAP7_75t_L g1585 ( .A1(n_1503), .A2(n_1581), .A3(n_1586), .B(n_1589), .Y(n_1585) );
AND2x2_ASAP7_75t_L g1626 ( .A(n_1503), .B(n_1515), .Y(n_1626) );
INVx2_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
NAND2xp5_ASAP7_75t_SL g1562 ( .A(n_1504), .B(n_1529), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_1504), .B(n_1584), .Y(n_1583) );
NAND2xp5_ASAP7_75t_L g1577 ( .A(n_1505), .B(n_1578), .Y(n_1577) );
OR2x2_ASAP7_75t_L g1643 ( .A(n_1506), .B(n_1522), .Y(n_1643) );
OAI211xp5_ASAP7_75t_L g1507 ( .A1(n_1508), .A2(n_1512), .B(n_1514), .C(n_1519), .Y(n_1507) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1510), .B(n_1511), .Y(n_1509) );
INVx2_ASAP7_75t_L g1551 ( .A(n_1510), .Y(n_1551) );
A2O1A1Ixp33_ASAP7_75t_L g1623 ( .A1(n_1510), .A2(n_1624), .B(n_1626), .C(n_1627), .Y(n_1623) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1511), .B(n_1572), .Y(n_1571) );
NOR2xp33_ASAP7_75t_SL g1575 ( .A(n_1511), .B(n_1576), .Y(n_1575) );
NOR2xp33_ASAP7_75t_L g1617 ( .A(n_1511), .B(n_1618), .Y(n_1617) );
O2A1O1Ixp33_ASAP7_75t_L g1608 ( .A1(n_1512), .A2(n_1609), .B(n_1610), .C(n_1611), .Y(n_1608) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
OAI21xp33_ASAP7_75t_L g1514 ( .A1(n_1515), .A2(n_1516), .B(n_1518), .Y(n_1514) );
NAND2xp5_ASAP7_75t_L g1602 ( .A(n_1518), .B(n_1534), .Y(n_1602) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1523), .Y(n_1579) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_1525), .A2(n_1532), .B1(n_1533), .B2(n_1535), .C(n_1537), .Y(n_1524) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
AOI22xp5_ASAP7_75t_L g1613 ( .A1(n_1532), .A2(n_1614), .B1(n_1619), .B2(n_1621), .Y(n_1613) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
CKINVDCx6p67_ASAP7_75t_R g1535 ( .A(n_1536), .Y(n_1535) );
NAND2xp5_ASAP7_75t_L g1592 ( .A(n_1536), .B(n_1593), .Y(n_1592) );
INVx3_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx2_ASAP7_75t_SL g1538 ( .A(n_1539), .Y(n_1538) );
OAI21xp33_ASAP7_75t_L g1567 ( .A1(n_1539), .A2(n_1568), .B(n_1570), .Y(n_1567) );
INVx2_ASAP7_75t_SL g1572 ( .A(n_1539), .Y(n_1572) );
OAI22xp5_ASAP7_75t_SL g1540 ( .A1(n_1541), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1540) );
INVx1_ASAP7_75t_L g1615 ( .A(n_1546), .Y(n_1615) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
AND2x2_ASAP7_75t_L g1554 ( .A(n_1550), .B(n_1555), .Y(n_1554) );
AND2x2_ASAP7_75t_L g1607 ( .A(n_1550), .B(n_1595), .Y(n_1607) );
NAND2xp5_ASAP7_75t_L g1636 ( .A(n_1550), .B(n_1637), .Y(n_1636) );
INVx2_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1556 ( .A(n_1557), .Y(n_1556) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
NAND5xp2_ASAP7_75t_L g1559 ( .A(n_1560), .B(n_1580), .C(n_1585), .D(n_1594), .E(n_1602), .Y(n_1559) );
AOI21xp5_ASAP7_75t_L g1560 ( .A1(n_1561), .A2(n_1571), .B(n_1573), .Y(n_1560) );
NAND2xp5_ASAP7_75t_L g1563 ( .A(n_1564), .B(n_1566), .Y(n_1563) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
NAND3xp33_ASAP7_75t_L g1624 ( .A(n_1569), .B(n_1590), .C(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
NAND2xp5_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1583), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
OAI22xp5_ASAP7_75t_L g1629 ( .A1(n_1582), .A2(n_1630), .B1(n_1631), .B2(n_1633), .Y(n_1629) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1584), .Y(n_1620) );
AOI21xp33_ASAP7_75t_L g1589 ( .A1(n_1588), .A2(n_1590), .B(n_1592), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1619 ( .A(n_1590), .B(n_1620), .Y(n_1619) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVxp67_ASAP7_75t_SL g1597 ( .A(n_1598), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1598 ( .A(n_1599), .B(n_1600), .Y(n_1598) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1599), .Y(n_1609) );
CKINVDCx14_ASAP7_75t_R g1610 ( .A(n_1601), .Y(n_1610) );
NAND5xp2_ASAP7_75t_L g1603 ( .A(n_1604), .B(n_1613), .C(n_1623), .D(n_1628), .E(n_1638), .Y(n_1603) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
NAND2xp5_ASAP7_75t_SL g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
INVxp67_ASAP7_75t_L g1616 ( .A(n_1617), .Y(n_1616) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
INVx1_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
CKINVDCx14_ASAP7_75t_R g1633 ( .A(n_1634), .Y(n_1633) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
OAI21xp5_ASAP7_75t_L g1638 ( .A1(n_1639), .A2(n_1641), .B(n_1644), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
INVxp67_ASAP7_75t_SL g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVx1_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1652 ( .A(n_1653), .Y(n_1652) );
endmodule