module fake_netlist_1_7838_n_697 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_697);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_697;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_56), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_51), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_20), .Y(n_79) );
INVxp33_ASAP7_75t_SL g80 ( .A(n_42), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_36), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_1), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_5), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_50), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_26), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_69), .Y(n_87) );
INVxp33_ASAP7_75t_L g88 ( .A(n_7), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_8), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_15), .Y(n_90) );
INVxp67_ASAP7_75t_L g91 ( .A(n_64), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_33), .Y(n_92) );
CKINVDCx14_ASAP7_75t_R g93 ( .A(n_54), .Y(n_93) );
HB1xp67_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_63), .Y(n_95) );
INVxp33_ASAP7_75t_L g96 ( .A(n_62), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_74), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_71), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_59), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_30), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_28), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_70), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_43), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_6), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_35), .Y(n_105) );
INVxp33_ASAP7_75t_L g106 ( .A(n_15), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_6), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_27), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_52), .Y(n_111) );
BUFx2_ASAP7_75t_L g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_48), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_38), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_72), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_37), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_1), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_53), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_29), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_68), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_112), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_124), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_112), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_94), .B(n_0), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_110), .Y(n_130) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_91), .B(n_0), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_110), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_124), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_93), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_100), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_77), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_80), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_88), .B(n_2), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_120), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_78), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_79), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_120), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_78), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_79), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_95), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_81), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_81), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_82), .Y(n_153) );
INVx3_ASAP7_75t_L g154 ( .A(n_123), .Y(n_154) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_85), .B(n_76), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_85), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_86), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_86), .B(n_32), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_87), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_82), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_83), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_87), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g164 ( .A(n_117), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_92), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_97), .Y(n_166) );
BUFx2_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_152), .Y(n_168) );
AND2x6_ASAP7_75t_L g169 ( .A(n_154), .B(n_123), .Y(n_169) );
AND2x2_ASAP7_75t_L g170 ( .A(n_146), .B(n_106), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_125), .B(n_96), .Y(n_171) );
INVx4_ASAP7_75t_SL g172 ( .A(n_158), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_141), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_146), .B(n_122), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_153), .Y(n_175) );
INVx1_ASAP7_75t_SL g176 ( .A(n_128), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_141), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_153), .B(n_122), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_160), .B(n_83), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
BUFx2_ASAP7_75t_L g181 ( .A(n_150), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_154), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
INVx1_ASAP7_75t_SL g185 ( .A(n_149), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_152), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_152), .Y(n_187) );
INVx8_ASAP7_75t_L g188 ( .A(n_158), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_126), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_126), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_126), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_142), .B(n_103), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_160), .B(n_119), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_143), .B(n_119), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g195 ( .A(n_134), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_138), .B(n_90), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_155), .A2(n_161), .B1(n_143), .B2(n_159), .Y(n_197) );
OAI22x1_ASAP7_75t_L g198 ( .A1(n_143), .A2(n_89), .B1(n_90), .B2(n_104), .Y(n_198) );
BUFx6f_ASAP7_75t_L g199 ( .A(n_152), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_126), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
CKINVDCx5p33_ASAP7_75t_R g204 ( .A(n_164), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_126), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_126), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_138), .B(n_104), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_126), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_139), .B(n_113), .Y(n_211) );
OAI22xp33_ASAP7_75t_SL g212 ( .A1(n_129), .A2(n_113), .B1(n_107), .B2(n_116), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_158), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_139), .B(n_121), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_133), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_148), .Y(n_216) );
NAND2x1p5_ASAP7_75t_L g217 ( .A(n_155), .B(n_121), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_148), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_158), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_133), .Y(n_220) );
INVx2_ASAP7_75t_SL g221 ( .A(n_165), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_145), .B(n_118), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_157), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_133), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_133), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_145), .B(n_118), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_151), .A2(n_116), .B1(n_115), .B2(n_114), .Y(n_228) );
BUFx4f_ASAP7_75t_L g229 ( .A(n_158), .Y(n_229) );
INVx3_ASAP7_75t_SL g230 ( .A(n_204), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_175), .B(n_131), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_175), .Y(n_232) );
NOR2xp33_ASAP7_75t_R g233 ( .A(n_204), .B(n_158), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_213), .Y(n_234) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_213), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_221), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_178), .B(n_131), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_206), .A2(n_151), .B1(n_163), .B2(n_162), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_181), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_178), .B(n_159), .Y(n_240) );
BUFx4f_ASAP7_75t_L g241 ( .A(n_217), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_221), .Y(n_242) );
INVxp67_ASAP7_75t_SL g243 ( .A(n_222), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_178), .B(n_163), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_213), .Y(n_245) );
OR2x2_ASAP7_75t_SL g246 ( .A(n_176), .B(n_162), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_193), .B(n_156), .Y(n_247) );
INVx5_ASAP7_75t_L g248 ( .A(n_169), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx5_ASAP7_75t_L g250 ( .A(n_169), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_196), .Y(n_251) );
AO22x1_ASAP7_75t_L g252 ( .A1(n_197), .A2(n_158), .B1(n_156), .B2(n_98), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_210), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_216), .Y(n_254) );
INVxp67_ASAP7_75t_SL g255 ( .A(n_222), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_216), .Y(n_256) );
NAND3xp33_ASAP7_75t_L g257 ( .A(n_171), .B(n_133), .C(n_165), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_214), .A2(n_165), .B(n_166), .C(n_157), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_193), .B(n_166), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_213), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_218), .Y(n_262) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_195), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_193), .B(n_135), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_224), .Y(n_267) );
INVxp67_ASAP7_75t_L g268 ( .A(n_170), .Y(n_268) );
NAND3xp33_ASAP7_75t_SL g269 ( .A(n_217), .B(n_114), .C(n_98), .Y(n_269) );
NOR3xp33_ASAP7_75t_SL g270 ( .A(n_195), .B(n_192), .C(n_177), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g271 ( .A1(n_206), .A2(n_158), .B1(n_166), .B2(n_137), .Y(n_271) );
BUFx12f_ASAP7_75t_L g272 ( .A(n_167), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_224), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_185), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_196), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_222), .B(n_137), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_170), .B(n_137), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_219), .B(n_115), .Y(n_280) );
CKINVDCx5p33_ASAP7_75t_R g281 ( .A(n_181), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_174), .B(n_135), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_219), .B(n_97), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_183), .Y(n_284) );
AOI22xp5_ASAP7_75t_L g285 ( .A1(n_217), .A2(n_158), .B1(n_147), .B2(n_144), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_167), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_211), .A2(n_147), .B1(n_144), .B2(n_140), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
O2A1O1Ixp33_ASAP7_75t_L g289 ( .A1(n_173), .A2(n_147), .B(n_144), .C(n_140), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_174), .Y(n_290) );
BUFx2_ASAP7_75t_L g291 ( .A(n_180), .Y(n_291) );
AND3x1_ASAP7_75t_SL g292 ( .A(n_198), .B(n_99), .C(n_101), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_208), .Y(n_293) );
NOR2xp33_ASAP7_75t_R g294 ( .A(n_188), .B(n_135), .Y(n_294) );
AO22x1_ASAP7_75t_L g295 ( .A1(n_180), .A2(n_111), .B1(n_101), .B2(n_102), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_243), .B(n_194), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_234), .Y(n_297) );
NOR2x1_ASAP7_75t_L g298 ( .A(n_269), .B(n_219), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_243), .B(n_194), .Y(n_299) );
AND2x2_ASAP7_75t_SL g300 ( .A(n_241), .B(n_229), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_255), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_255), .B(n_179), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_290), .B(n_179), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_232), .B(n_208), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_249), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_293), .B(n_172), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_248), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_253), .Y(n_308) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_248), .B(n_229), .Y(n_309) );
NOR2xp33_ASAP7_75t_L g310 ( .A(n_268), .B(n_212), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_254), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_239), .B(n_172), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_256), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_248), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_251), .Y(n_316) );
INVx4_ASAP7_75t_L g317 ( .A(n_248), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_259), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_290), .A2(n_169), .B1(n_198), .B2(n_188), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_250), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_240), .B(n_169), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_262), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_268), .B(n_229), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_247), .B(n_169), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_274), .B(n_227), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_238), .A2(n_188), .B1(n_213), .B2(n_228), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_264), .Y(n_327) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_230), .Y(n_328) );
BUFx4f_ASAP7_75t_SL g329 ( .A(n_272), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_266), .Y(n_330) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_258), .A2(n_203), .B(n_201), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_265), .B(n_169), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_265), .B(n_172), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_251), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_244), .A2(n_188), .B(n_202), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g336 ( .A1(n_280), .A2(n_283), .B(n_260), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_250), .B(n_172), .Y(n_337) );
AND2x4_ASAP7_75t_L g338 ( .A(n_276), .B(n_135), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_267), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_276), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_273), .Y(n_341) );
AND2x4_ASAP7_75t_L g342 ( .A(n_282), .B(n_140), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_282), .B(n_136), .Y(n_343) );
AOI222xp33_ASAP7_75t_L g344 ( .A1(n_286), .A2(n_136), .B1(n_127), .B2(n_105), .C1(n_108), .C2(n_99), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_275), .B(n_127), .Y(n_345) );
CKINVDCx14_ASAP7_75t_R g346 ( .A(n_281), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_301), .B(n_238), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_301), .B(n_277), .Y(n_348) );
AND2x2_ASAP7_75t_SL g349 ( .A(n_300), .B(n_241), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_303), .A2(n_230), .B1(n_291), .B2(n_269), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_303), .A2(n_288), .B1(n_263), .B2(n_237), .Y(n_351) );
CKINVDCx6p67_ASAP7_75t_R g352 ( .A(n_325), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_329), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_305), .Y(n_354) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_297), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_305), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g358 ( .A(n_315), .B(n_250), .Y(n_358) );
AO31x2_ASAP7_75t_L g359 ( .A1(n_308), .A2(n_136), .A3(n_127), .B(n_215), .Y(n_359) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_310), .A2(n_279), .B1(n_295), .B2(n_270), .C(n_231), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_325), .A2(n_271), .B1(n_285), .B2(n_278), .Y(n_361) );
OAI221xp5_ASAP7_75t_L g362 ( .A1(n_302), .A2(n_270), .B1(n_287), .B2(n_289), .C(n_257), .Y(n_362) );
BUFx2_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_297), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_296), .B(n_299), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_307), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_318), .B(n_252), .Y(n_367) );
AOI21xp5_ASAP7_75t_L g368 ( .A1(n_331), .A2(n_284), .B(n_242), .Y(n_368) );
CKINVDCx11_ASAP7_75t_R g369 ( .A(n_346), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_304), .A2(n_287), .B1(n_236), .B2(n_233), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_304), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_328), .A2(n_246), .B1(n_233), .B2(n_294), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_318), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_304), .A2(n_294), .B1(n_250), .B2(n_102), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g375 ( .A1(n_323), .A2(n_105), .B(n_108), .C(n_111), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_297), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_327), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_297), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_365), .B(n_327), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_354), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_352), .A2(n_319), .B1(n_344), .B2(n_342), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_351), .A2(n_326), .B1(n_321), .B2(n_324), .C(n_341), .Y(n_382) );
OAI22xp5_ASAP7_75t_L g383 ( .A1(n_365), .A2(n_313), .B1(n_311), .B2(n_322), .Y(n_383) );
OAI211xp5_ASAP7_75t_L g384 ( .A1(n_360), .A2(n_343), .B(n_330), .C(n_341), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_369), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_352), .A2(n_330), .B1(n_334), .B2(n_342), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_354), .Y(n_387) );
OAI22xp33_ASAP7_75t_L g388 ( .A1(n_371), .A2(n_311), .B1(n_322), .B2(n_313), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_360), .A2(n_342), .B1(n_338), .B2(n_345), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_368), .A2(n_314), .B(n_297), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_347), .A2(n_338), .B1(n_345), .B2(n_343), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_356), .B(n_339), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_347), .A2(n_338), .B1(n_345), .B2(n_339), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_362), .A2(n_340), .B1(n_316), .B2(n_336), .C(n_334), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_356), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_371), .B(n_316), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_368), .A2(n_225), .B(n_220), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_375), .A2(n_298), .B(n_335), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_357), .Y(n_399) );
AO21x2_ASAP7_75t_L g400 ( .A1(n_367), .A2(n_225), .B(n_220), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_350), .A2(n_298), .B(n_332), .Y(n_401) );
OAI22xp33_ASAP7_75t_L g402 ( .A1(n_363), .A2(n_340), .B1(n_316), .B2(n_292), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_349), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_361), .A2(n_292), .B1(n_300), .B2(n_340), .Y(n_404) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_362), .A2(n_300), .B1(n_312), .B2(n_333), .Y(n_405) );
AOI211xp5_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_312), .B(n_333), .C(n_133), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_397), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_380), .Y(n_408) );
OAI211xp5_ASAP7_75t_L g409 ( .A1(n_381), .A2(n_372), .B(n_377), .C(n_373), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_383), .A2(n_373), .B1(n_377), .B2(n_357), .Y(n_410) );
INVxp67_ASAP7_75t_L g411 ( .A(n_379), .Y(n_411) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_403), .A2(n_348), .B1(n_367), .B2(n_353), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_380), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_379), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_392), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_399), .B(n_348), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_389), .A2(n_349), .B1(n_370), .B2(n_374), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_403), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_392), .B(n_359), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_387), .B(n_359), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_387), .Y(n_421) );
NAND3xp33_ASAP7_75t_L g422 ( .A(n_394), .B(n_207), .C(n_366), .Y(n_422) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_403), .B(n_355), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_395), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_395), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_399), .B(n_359), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_386), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_393), .A2(n_349), .B1(n_366), .B2(n_355), .Y(n_428) );
OAI211xp5_ASAP7_75t_L g429 ( .A1(n_404), .A2(n_366), .B(n_215), .C(n_226), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_402), .A2(n_312), .B1(n_306), .B2(n_364), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_391), .B(n_359), .Y(n_431) );
AOI222xp33_ASAP7_75t_L g432 ( .A1(n_384), .A2(n_312), .B1(n_306), .B2(n_309), .C1(n_5), .C2(n_8), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_397), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_404), .B(n_359), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_405), .B(n_364), .Y(n_435) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_401), .A2(n_306), .B1(n_376), .B2(n_364), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_396), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g438 ( .A1(n_382), .A2(n_168), .B1(n_182), .B2(n_184), .C(n_186), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_400), .Y(n_439) );
OAI221xp5_ASAP7_75t_L g440 ( .A1(n_405), .A2(n_358), .B1(n_226), .B2(n_184), .C(n_182), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_406), .A2(n_378), .B(n_376), .C(n_307), .Y(n_442) );
INVx4_ASAP7_75t_L g443 ( .A(n_418), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_419), .B(n_359), .Y(n_444) );
AOI31xp33_ASAP7_75t_L g445 ( .A1(n_432), .A2(n_385), .A3(n_388), .B(n_358), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_424), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_400), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_426), .B(n_400), .Y(n_448) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_422), .A2(n_390), .B(n_398), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_425), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_425), .Y(n_451) );
INVx4_ASAP7_75t_L g452 ( .A(n_418), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_SL g453 ( .A1(n_429), .A2(n_168), .B(n_186), .C(n_187), .Y(n_453) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_411), .B(n_385), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_418), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_414), .B(n_2), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_418), .Y(n_457) );
NAND2x1_ASAP7_75t_L g458 ( .A(n_421), .B(n_397), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_426), .B(n_397), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_408), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_432), .B(n_187), .C(n_189), .D(n_190), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_420), .B(n_378), .Y(n_462) );
BUFx2_ASAP7_75t_L g463 ( .A(n_425), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_409), .A2(n_358), .B(n_190), .Y(n_465) );
OAI33xp33_ASAP7_75t_L g466 ( .A1(n_412), .A2(n_3), .A3(n_4), .B1(n_9), .B2(n_10), .B3(n_11), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
NOR2x1_ASAP7_75t_L g468 ( .A(n_422), .B(n_420), .Y(n_468) );
OAI31xp33_ASAP7_75t_L g469 ( .A1(n_427), .A2(n_378), .A3(n_376), .B(n_337), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_415), .B(n_3), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_413), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_424), .B(n_4), .Y(n_472) );
NAND4xp25_ASAP7_75t_L g473 ( .A(n_427), .B(n_189), .C(n_191), .D(n_200), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_434), .B(n_9), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_407), .Y(n_475) );
AOI21xp33_ASAP7_75t_SL g476 ( .A1(n_428), .A2(n_11), .B(n_12), .Y(n_476) );
AOI31xp33_ASAP7_75t_L g477 ( .A1(n_428), .A2(n_12), .A3(n_13), .B(n_14), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_421), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_437), .B(n_13), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_407), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_434), .B(n_14), .Y(n_483) );
AND2x4_ASAP7_75t_L g484 ( .A(n_435), .B(n_355), .Y(n_484) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
AOI33xp33_ASAP7_75t_L g486 ( .A1(n_431), .A2(n_209), .A3(n_200), .B1(n_205), .B2(n_191), .B3(n_19), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_415), .B(n_16), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_423), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_427), .A2(n_355), .B1(n_320), .B2(n_317), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_416), .B(n_16), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_431), .B(n_17), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_417), .A2(n_355), .B1(n_320), .B2(n_317), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_474), .B(n_437), .Y(n_494) );
NOR3xp33_ASAP7_75t_L g495 ( .A(n_466), .B(n_440), .C(n_410), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_460), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_474), .B(n_441), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_444), .B(n_435), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_483), .B(n_441), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_464), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_444), .B(n_435), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_464), .Y(n_504) );
OR2x4_ASAP7_75t_L g505 ( .A(n_445), .B(n_416), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_447), .B(n_435), .Y(n_506) );
AND2x4_ASAP7_75t_L g507 ( .A(n_443), .B(n_423), .Y(n_507) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_446), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_475), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_483), .A2(n_417), .B1(n_440), .B2(n_410), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_467), .Y(n_511) );
INVxp67_ASAP7_75t_L g512 ( .A(n_454), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_467), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g515 ( .A1(n_477), .A2(n_441), .B1(n_430), .B2(n_438), .C(n_436), .Y(n_515) );
INVx1_ASAP7_75t_SL g516 ( .A(n_489), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_456), .A2(n_442), .B1(n_433), .B2(n_199), .C(n_207), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_492), .B(n_423), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_492), .B(n_447), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_471), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_462), .B(n_433), .Y(n_521) );
AOI31xp33_ASAP7_75t_L g522 ( .A1(n_476), .A2(n_18), .A3(n_19), .B(n_209), .Y(n_522) );
INVx4_ASAP7_75t_L g523 ( .A(n_443), .Y(n_523) );
INVxp67_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_451), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_462), .B(n_18), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_448), .B(n_205), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_480), .B(n_355), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_472), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_448), .B(n_207), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_491), .B(n_207), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_472), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_478), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_478), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_459), .B(n_207), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_481), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_481), .Y(n_538) );
NAND2xp33_ASAP7_75t_SL g539 ( .A(n_443), .B(n_320), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_452), .B(n_21), .Y(n_540) );
CKINVDCx16_ASAP7_75t_R g541 ( .A(n_452), .Y(n_541) );
NAND3xp33_ASAP7_75t_L g542 ( .A(n_476), .B(n_199), .C(n_314), .Y(n_542) );
AND2x2_ASAP7_75t_SL g543 ( .A(n_463), .B(n_317), .Y(n_543) );
AOI21xp5_ASAP7_75t_SL g544 ( .A1(n_452), .A2(n_315), .B(n_314), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_488), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_463), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_459), .B(n_199), .Y(n_547) );
AOI211xp5_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_199), .B(n_314), .C(n_34), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_488), .B(n_22), .Y(n_549) );
OAI222xp33_ASAP7_75t_L g550 ( .A1(n_468), .A2(n_315), .B1(n_39), .B2(n_41), .C1(n_44), .C2(n_45), .Y(n_550) );
NAND2x1_ASAP7_75t_SL g551 ( .A(n_455), .B(n_24), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_479), .B(n_46), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g553 ( .A1(n_524), .A2(n_487), .B1(n_461), .B2(n_493), .C(n_473), .Y(n_553) );
INVxp67_ASAP7_75t_SL g554 ( .A(n_525), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_497), .Y(n_555) );
NAND2xp33_ASAP7_75t_SL g556 ( .A(n_523), .B(n_450), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_509), .Y(n_557) );
OAI221xp5_ASAP7_75t_L g558 ( .A1(n_512), .A2(n_469), .B1(n_468), .B2(n_490), .C(n_450), .Y(n_558) );
OAI21xp5_ASAP7_75t_SL g559 ( .A1(n_522), .A2(n_510), .B(n_505), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_530), .B(n_486), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_505), .B(n_455), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_544), .A2(n_458), .B(n_453), .Y(n_564) );
AND2x4_ASAP7_75t_L g565 ( .A(n_523), .B(n_455), .Y(n_565) );
NAND3xp33_ASAP7_75t_L g566 ( .A(n_495), .B(n_465), .C(n_457), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_533), .B(n_457), .C(n_485), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_519), .B(n_534), .Y(n_568) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_539), .A2(n_457), .B(n_458), .C(n_482), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_535), .B(n_482), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_518), .B(n_499), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_510), .A2(n_479), .B(n_484), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_496), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_499), .B(n_484), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_508), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_504), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_511), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_516), .B(n_484), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_503), .B(n_485), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
OAI21xp33_ASAP7_75t_L g583 ( .A1(n_546), .A2(n_485), .B(n_199), .Y(n_583) );
AOI22x1_ASAP7_75t_L g584 ( .A1(n_541), .A2(n_485), .B1(n_314), .B2(n_57), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_494), .B(n_485), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_520), .B(n_449), .Y(n_586) );
OAI32xp33_ASAP7_75t_L g587 ( .A1(n_523), .A2(n_449), .A3(n_55), .B1(n_58), .B2(n_60), .Y(n_587) );
OA21x2_ASAP7_75t_L g588 ( .A1(n_536), .A2(n_449), .B(n_61), .Y(n_588) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_542), .B(n_261), .C(n_245), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_526), .B(n_47), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_537), .B(n_65), .Y(n_591) );
NAND4xp25_ASAP7_75t_SL g592 ( .A(n_515), .B(n_66), .C(n_67), .D(n_73), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_538), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_545), .Y(n_594) );
AND2x2_ASAP7_75t_SL g595 ( .A(n_507), .B(n_543), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_527), .A2(n_75), .B1(n_234), .B2(n_235), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_528), .B(n_234), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_528), .Y(n_599) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_548), .B(n_235), .C(n_245), .Y(n_600) );
O2A1O1Ixp5_ASAP7_75t_L g601 ( .A1(n_539), .A2(n_235), .B(n_245), .C(n_261), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_550), .A2(n_235), .B(n_245), .C(n_261), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_503), .A2(n_261), .B(n_506), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_506), .B(n_498), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_568), .B(n_531), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_604), .B(n_581), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_571), .B(n_521), .Y(n_607) );
NAND2xp5_ASAP7_75t_SL g608 ( .A(n_595), .B(n_543), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_595), .B(n_507), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_562), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_555), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_574), .B(n_531), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_562), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_575), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_599), .B(n_513), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_557), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_576), .Y(n_617) );
AND4x1_ASAP7_75t_L g618 ( .A(n_561), .B(n_544), .C(n_517), .D(n_500), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_565), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_554), .B(n_513), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_554), .B(n_547), .Y(n_621) );
NAND2x1_ASAP7_75t_L g622 ( .A(n_565), .B(n_507), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_575), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_577), .B(n_529), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_578), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_598), .Y(n_626) );
XNOR2xp5_ASAP7_75t_L g627 ( .A(n_556), .B(n_540), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_585), .B(n_549), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_563), .B(n_549), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_579), .Y(n_630) );
NOR2xp33_ASAP7_75t_SL g631 ( .A(n_559), .B(n_540), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_580), .Y(n_632) );
XNOR2x1_ASAP7_75t_L g633 ( .A(n_560), .B(n_540), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_582), .B(n_532), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_593), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_573), .B(n_552), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_570), .Y(n_638) );
OR2x2_ASAP7_75t_L g639 ( .A(n_573), .B(n_552), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_572), .B(n_551), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_638), .B(n_586), .Y(n_641) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_633), .B(n_627), .Y(n_642) );
OAI21xp33_ASAP7_75t_SL g643 ( .A1(n_609), .A2(n_564), .B(n_592), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_631), .A2(n_558), .B1(n_603), .B2(n_566), .C(n_553), .Y(n_644) );
A2O1A1Ixp33_ASAP7_75t_L g645 ( .A1(n_608), .A2(n_602), .B(n_564), .C(n_583), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_635), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_635), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_638), .B(n_567), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_626), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_626), .B(n_569), .Y(n_650) );
AOI22xp33_ASAP7_75t_SL g651 ( .A1(n_633), .A2(n_584), .B1(n_588), .B2(n_600), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_610), .B(n_588), .Y(n_652) );
NAND4xp75_ASAP7_75t_L g653 ( .A(n_640), .B(n_601), .C(n_596), .D(n_590), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_630), .Y(n_654) );
INVx2_ASAP7_75t_SL g655 ( .A(n_622), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_614), .Y(n_656) );
INVxp67_ASAP7_75t_L g657 ( .A(n_614), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_606), .B(n_607), .Y(n_658) );
AOI211xp5_ASAP7_75t_SL g659 ( .A1(n_619), .A2(n_591), .B(n_597), .C(n_602), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_630), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_637), .Y(n_661) );
INVx1_ASAP7_75t_SL g662 ( .A(n_632), .Y(n_662) );
AO21x1_ASAP7_75t_L g663 ( .A1(n_622), .A2(n_589), .B(n_601), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g664 ( .A(n_655), .B(n_627), .Y(n_664) );
BUFx12f_ASAP7_75t_L g665 ( .A(n_655), .Y(n_665) );
INVx1_ASAP7_75t_SL g666 ( .A(n_662), .Y(n_666) );
AOI221xp5_ASAP7_75t_L g667 ( .A1(n_644), .A2(n_617), .B1(n_625), .B2(n_611), .C(n_623), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g668 ( .A1(n_645), .A2(n_623), .B(n_610), .C(n_613), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_649), .B(n_613), .Y(n_669) );
NAND3x1_ASAP7_75t_L g670 ( .A(n_642), .B(n_619), .C(n_618), .Y(n_670) );
NOR4xp25_ASAP7_75t_L g671 ( .A(n_643), .B(n_637), .C(n_620), .D(n_621), .Y(n_671) );
OAI31xp33_ASAP7_75t_L g672 ( .A1(n_642), .A2(n_619), .A3(n_607), .B(n_612), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_658), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_657), .A2(n_650), .B1(n_641), .B2(n_658), .C1(n_648), .C2(n_652), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_651), .B(n_587), .C(n_634), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_654), .B(n_615), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_660), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_663), .A2(n_639), .B(n_636), .C(n_605), .Y(n_678) );
INVx2_ASAP7_75t_L g679 ( .A(n_656), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_661), .Y(n_680) );
OAI21xp33_ASAP7_75t_SL g681 ( .A1(n_656), .A2(n_606), .B(n_612), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g682 ( .A1(n_646), .A2(n_624), .B1(n_615), .B2(n_628), .C(n_616), .Y(n_682) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_645), .A2(n_639), .B1(n_636), .B2(n_628), .Y(n_683) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_659), .B(n_647), .C(n_616), .Y(n_684) );
OAI211xp5_ASAP7_75t_SL g685 ( .A1(n_653), .A2(n_629), .B(n_644), .C(n_559), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_666), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_667), .B(n_674), .Y(n_687) );
OR4x2_ASAP7_75t_L g688 ( .A(n_670), .B(n_672), .C(n_671), .D(n_685), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g689 ( .A1(n_668), .A2(n_683), .B1(n_678), .B2(n_664), .C(n_675), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_686), .Y(n_690) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_689), .B(n_684), .C(n_681), .Y(n_691) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_687), .B(n_682), .C(n_680), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_690), .Y(n_693) );
AND2x2_ASAP7_75t_L g694 ( .A(n_691), .B(n_665), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_693), .A2(n_692), .B1(n_688), .B2(n_663), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g696 ( .A1(n_695), .A2(n_694), .B1(n_679), .B2(n_673), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_677), .B1(n_669), .B2(n_676), .C(n_629), .Y(n_697) );
endmodule