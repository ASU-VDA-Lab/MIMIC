module fake_ibex_83_n_964 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_964);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_964;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_845;
wire n_947;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_375;
wire n_317;
wire n_340;
wire n_280;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_278;
wire n_242;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_185;
wire n_388;
wire n_953;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_797;
wire n_796;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_801;
wire n_918;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_581;
wire n_416;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_955;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_392;
wire n_206;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_188;
wire n_200;
wire n_506;
wire n_444;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_927;
wire n_934;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_285;
wire n_320;
wire n_247;
wire n_379;
wire n_288;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_385;
wire n_233;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_631;
wire n_683;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_874;
wire n_890;
wire n_912;
wire n_921;
wire n_816;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_231;
wire n_298;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_69),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_92),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_60),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_30),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_71),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_4),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_67),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_52),
.Y(n_186)
);

INVxp33_ASAP7_75t_SL g187 ( 
.A(n_25),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_114),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_126),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_90),
.B(n_150),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_78),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_125),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_48),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_80),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_66),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_102),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_135),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_155),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_54),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_3),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_99),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_106),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_26),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_65),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_134),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_154),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_137),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_62),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_74),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_59),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_8),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_122),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_55),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_107),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_25),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_27),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_81),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_105),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_47),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_17),
.B(n_84),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_91),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_131),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_22),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_95),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_161),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_6),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_108),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_29),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_75),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_35),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_93),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_9),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_39),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_103),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_79),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_144),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_15),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_1),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_133),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_120),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_170),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_82),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_173),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_72),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_53),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_109),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_64),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_151),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_124),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_73),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_13),
.B(n_164),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_153),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_3),
.B(n_77),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_87),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_63),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_119),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g280 ( 
.A(n_76),
.B(n_116),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_7),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g283 ( 
.A(n_88),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_43),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_26),
.Y(n_286)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_49),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_L g288 ( 
.A(n_96),
.B(n_47),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_40),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_110),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_143),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_50),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_152),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_49),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_233),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_0),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_184),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_245),
.B(n_2),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_287),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_184),
.A2(n_6),
.B1(n_8),
.B2(n_10),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_233),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_202),
.Y(n_303)
);

OAI22x1_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_230),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_210),
.B(n_13),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_230),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_178),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_273),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_233),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_175),
.B(n_182),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_261),
.B(n_14),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_179),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_175),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_268),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_180),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_178),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_183),
.B(n_16),
.Y(n_319)
);

CKINVDCx11_ASAP7_75t_R g320 ( 
.A(n_258),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_178),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_193),
.B(n_207),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_188),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_233),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

OA21x2_ASAP7_75t_L g327 ( 
.A1(n_182),
.A2(n_83),
.B(n_169),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_189),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_197),
.Y(n_329)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_178),
.Y(n_331)
);

AND2x2_ASAP7_75t_R g332 ( 
.A(n_258),
.B(n_17),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_226),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_187),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_186),
.B(n_204),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_207),
.B(n_19),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g338 ( 
.A1(n_186),
.A2(n_85),
.B(n_165),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_202),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_207),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_281),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_209),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_209),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_226),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_226),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_198),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_244),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_176),
.B(n_20),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_294),
.B(n_181),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_199),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_204),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_201),
.B(n_23),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_283),
.B(n_23),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_244),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_223),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_223),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_187),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_360)
);

OA21x2_ASAP7_75t_L g361 ( 
.A1(n_263),
.A2(n_89),
.B(n_160),
.Y(n_361)
);

CKINVDCx8_ASAP7_75t_R g362 ( 
.A(n_174),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_216),
.B(n_28),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_283),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_224),
.B(n_29),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_205),
.Y(n_367)
);

CKINVDCx11_ASAP7_75t_R g368 ( 
.A(n_241),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_231),
.B(n_30),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_242),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_263),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_283),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_211),
.Y(n_374)
);

AND2x6_ASAP7_75t_L g375 ( 
.A(n_291),
.B(n_51),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_283),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_283),
.Y(n_377)
);

OA21x2_ASAP7_75t_L g378 ( 
.A1(n_291),
.A2(n_97),
.B(n_159),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_293),
.B(n_31),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_213),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_241),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_381)
);

BUFx8_ASAP7_75t_L g382 ( 
.A(n_283),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_293),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_215),
.Y(n_384)
);

OA21x2_ASAP7_75t_L g385 ( 
.A1(n_217),
.A2(n_98),
.B(n_158),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_218),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_326),
.B(n_174),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_354),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_379),
.A2(n_351),
.B1(n_365),
.B2(n_363),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_379),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_195),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_296),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_351),
.A2(n_246),
.B1(n_251),
.B2(n_252),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_310),
.B(n_266),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_296),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_300),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_300),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_312),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_354),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_286),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_363),
.A2(n_365),
.B1(n_369),
.B2(n_337),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_326),
.B(n_191),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_312),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_354),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g412 ( 
.A(n_343),
.B(n_289),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_326),
.B(n_191),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_303),
.B(n_257),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_358),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_358),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_309),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_375),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

AND3x2_ASAP7_75t_L g421 ( 
.A(n_340),
.B(n_254),
.C(n_232),
.Y(n_421)
);

OR2x6_ASAP7_75t_L g422 ( 
.A(n_340),
.B(n_285),
.Y(n_422)
);

OR2x6_ASAP7_75t_L g423 ( 
.A(n_337),
.B(n_292),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_SL g424 ( 
.A1(n_314),
.A2(n_324),
.B(n_317),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_323),
.B(n_235),
.Y(n_425)
);

BUFx2_ASAP7_75t_L g426 ( 
.A(n_323),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g427 ( 
.A1(n_369),
.A2(n_244),
.B1(n_239),
.B2(n_284),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_339),
.B(n_203),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_315),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_330),
.B(n_314),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_359),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_342),
.A2(n_266),
.B1(n_249),
.B2(n_236),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_324),
.A2(n_247),
.B1(n_279),
.B2(n_277),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_330),
.B(n_194),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_383),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_382),
.B(n_219),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_384),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_328),
.B(n_196),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_384),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_328),
.B(n_214),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_386),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_309),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_306),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_382),
.B(n_220),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_345),
.B(n_346),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_309),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_305),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_362),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_382),
.B(n_221),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_329),
.B(n_262),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_382),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_371),
.Y(n_460)
);

CKINVDCx14_ASAP7_75t_R g461 ( 
.A(n_368),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_362),
.B(n_262),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_329),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_349),
.B(n_265),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_349),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_353),
.B(n_222),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_371),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_367),
.B(n_274),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_372),
.A2(n_260),
.B1(n_238),
.B2(n_234),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_372),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_374),
.A2(n_237),
.B1(n_229),
.B2(n_243),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_295),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_374),
.B(n_267),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_302),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_302),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_320),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_309),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_345),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_307),
.Y(n_480)
);

OAI22xp33_ASAP7_75t_L g481 ( 
.A1(n_301),
.A2(n_276),
.B1(n_288),
.B2(n_275),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_346),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_307),
.Y(n_483)
);

OR2x6_ASAP7_75t_L g484 ( 
.A(n_304),
.B(n_248),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_311),
.Y(n_485)
);

CKINVDCx11_ASAP7_75t_R g486 ( 
.A(n_332),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_322),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_322),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_308),
.B(n_185),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_318),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_325),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_325),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_297),
.A2(n_269),
.B1(n_250),
.B2(n_225),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_341),
.Y(n_494)
);

CKINVDCx6p67_ASAP7_75t_R g495 ( 
.A(n_299),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_308),
.B(n_200),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_313),
.A2(n_270),
.B1(n_255),
.B2(n_227),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_364),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_364),
.B(n_228),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_373),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_319),
.A2(n_272),
.B1(n_264),
.B2(n_253),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_375),
.B(n_192),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_318),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_376),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_377),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_318),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_316),
.A2(n_256),
.B1(n_259),
.B2(n_271),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_355),
.B(n_208),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_390),
.A2(n_301),
.B1(n_298),
.B2(n_335),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_459),
.B(n_212),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_387),
.B(n_356),
.Y(n_513)
);

NOR2x2_ASAP7_75t_L g514 ( 
.A(n_414),
.B(n_381),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_432),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_439),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_441),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_452),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_426),
.A2(n_381),
.B1(n_360),
.B2(n_370),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_405),
.B(n_177),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_413),
.B(n_190),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_425),
.B(n_240),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_448),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_389),
.A2(n_375),
.B1(n_378),
.B2(n_338),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_464),
.A2(n_375),
.B1(n_290),
.B2(n_338),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_408),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_463),
.B(n_280),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_464),
.B(n_327),
.Y(n_530)
);

NAND2x1p5_ASAP7_75t_L g531 ( 
.A(n_420),
.B(n_327),
.Y(n_531)
);

OAI21xp5_ASAP7_75t_L g532 ( 
.A1(n_502),
.A2(n_378),
.B(n_361),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_338),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_401),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_428),
.B(n_338),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_437),
.A2(n_378),
.B(n_361),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_473),
.B(n_318),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_391),
.A2(n_470),
.B1(n_479),
.B2(n_465),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_473),
.A2(n_378),
.B1(n_361),
.B2(n_385),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_435),
.B(n_350),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_404),
.A2(n_366),
.B1(n_357),
.B2(n_361),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_431),
.B(n_357),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_407),
.B(n_321),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_423),
.A2(n_385),
.B1(n_366),
.B2(n_357),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_431),
.B(n_442),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_409),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_458),
.B(n_366),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_394),
.B(n_385),
.Y(n_550)
);

NAND2x1p5_ASAP7_75t_L g551 ( 
.A(n_462),
.B(n_321),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_423),
.A2(n_348),
.B1(n_347),
.B2(n_334),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_438),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_440),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_423),
.A2(n_348),
.B1(n_347),
.B2(n_334),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_419),
.Y(n_556)
);

AND2x6_ASAP7_75t_SL g557 ( 
.A(n_484),
.B(n_34),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_395),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_SL g559 ( 
.A(n_418),
.B(n_348),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_398),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_443),
.Y(n_562)
);

NOR3xp33_ASAP7_75t_L g563 ( 
.A(n_481),
.B(n_35),
.C(n_36),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_453),
.B(n_348),
.Y(n_564)
);

OR2x2_ASAP7_75t_L g565 ( 
.A(n_403),
.B(n_36),
.Y(n_565)
);

NOR2x1p5_ASAP7_75t_L g566 ( 
.A(n_478),
.B(n_37),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_424),
.A2(n_347),
.B1(n_334),
.B2(n_333),
.Y(n_567)
);

BUFx12f_ASAP7_75t_L g568 ( 
.A(n_486),
.Y(n_568)
);

NOR3xp33_ASAP7_75t_L g569 ( 
.A(n_508),
.B(n_38),
.C(n_39),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_400),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_446),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_347),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_461),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_429),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_509),
.B(n_334),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_333),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_500),
.B(n_333),
.Y(n_577)
);

AND2x2_ASAP7_75t_SL g578 ( 
.A(n_418),
.B(n_333),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_468),
.Y(n_579)
);

OAI221xp5_ASAP7_75t_L g580 ( 
.A1(n_396),
.A2(n_331),
.B1(n_321),
.B2(n_41),
.C(n_42),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_489),
.B(n_496),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_472),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_422),
.B(n_38),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_497),
.B(n_331),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_437),
.B(n_331),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_501),
.B(n_331),
.Y(n_586)
);

O2A1O1Ixp5_ASAP7_75t_L g587 ( 
.A1(n_449),
.A2(n_111),
.B(n_148),
.C(n_147),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_484),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_434),
.B(n_45),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_449),
.B(n_112),
.Y(n_590)
);

BUFx12f_ASAP7_75t_L g591 ( 
.A(n_486),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_493),
.B(n_113),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_422),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_469),
.B(n_45),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_422),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_412),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_471),
.B(n_56),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_466),
.B(n_57),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_454),
.B(n_58),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_484),
.B(n_61),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_433),
.B(n_70),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_596),
.B(n_495),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_530),
.A2(n_537),
.B(n_536),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_596),
.B(n_495),
.Y(n_605)
);

O2A1O1Ixp33_ASAP7_75t_L g606 ( 
.A1(n_510),
.A2(n_499),
.B(n_482),
.C(n_427),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_547),
.B(n_468),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_539),
.B(n_421),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_512),
.Y(n_609)
);

OAI22xp5_ASAP7_75t_L g610 ( 
.A1(n_547),
.A2(n_478),
.B1(n_397),
.B2(n_450),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_522),
.B(n_523),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_583),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_544),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_540),
.A2(n_498),
.B(n_487),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_517),
.Y(n_615)
);

AO32x1_ASAP7_75t_L g616 ( 
.A1(n_542),
.A2(n_411),
.A3(n_388),
.B1(n_402),
.B2(n_406),
.Y(n_616)
);

BUFx3_ASAP7_75t_L g617 ( 
.A(n_573),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_522),
.B(n_492),
.Y(n_618)
);

OAI22xp5_ASAP7_75t_L g619 ( 
.A1(n_602),
.A2(n_488),
.B1(n_474),
.B2(n_505),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_L g620 ( 
.A1(n_525),
.A2(n_494),
.B(n_506),
.C(n_504),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_525),
.A2(n_491),
.B(n_506),
.C(n_504),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_523),
.B(n_488),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_546),
.B(n_474),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_593),
.B(n_485),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_583),
.B(n_593),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_556),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_581),
.B(n_485),
.Y(n_627)
);

INVx11_ASAP7_75t_L g628 ( 
.A(n_568),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g629 ( 
.A1(n_595),
.A2(n_475),
.B1(n_491),
.B2(n_480),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_513),
.A2(n_475),
.B(n_480),
.C(n_483),
.Y(n_630)
);

CKINVDCx11_ASAP7_75t_R g631 ( 
.A(n_591),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_565),
.B(n_483),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_601),
.B(n_507),
.Y(n_633)
);

A2O1A1Ixp33_ASAP7_75t_L g634 ( 
.A1(n_513),
.A2(n_444),
.B(n_406),
.C(n_410),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_526),
.A2(n_444),
.B(n_410),
.Y(n_635)
);

OA22x2_ASAP7_75t_L g636 ( 
.A1(n_521),
.A2(n_467),
.B1(n_460),
.B2(n_457),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_515),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_595),
.A2(n_460),
.B1(n_456),
.B2(n_455),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_L g639 ( 
.A1(n_550),
.A2(n_415),
.B(n_455),
.C(n_416),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_519),
.Y(n_640)
);

OA21x2_ASAP7_75t_L g641 ( 
.A1(n_545),
.A2(n_416),
.B(n_451),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_558),
.A2(n_503),
.B(n_490),
.C(n_477),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_524),
.B(n_490),
.Y(n_643)
);

A2O1A1Ixp33_ASAP7_75t_L g644 ( 
.A1(n_560),
.A2(n_477),
.B(n_451),
.C(n_447),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_516),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_602),
.A2(n_451),
.B1(n_447),
.B2(n_417),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_561),
.A2(n_451),
.B(n_447),
.C(n_417),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_602),
.A2(n_417),
.B1(n_393),
.B2(n_447),
.Y(n_648)
);

AOI221xp5_ASAP7_75t_L g649 ( 
.A1(n_518),
.A2(n_579),
.B1(n_599),
.B2(n_563),
.C(n_569),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_570),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_601),
.A2(n_393),
.B1(n_100),
.B2(n_104),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_531),
.A2(n_115),
.B(n_117),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_534),
.B(n_127),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_528),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_130),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_601),
.B(n_136),
.Y(n_656)
);

BUFx6f_ASAP7_75t_L g657 ( 
.A(n_544),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_548),
.B(n_520),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_566),
.B(n_146),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_578),
.B(n_138),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g661 ( 
.A1(n_535),
.A2(n_140),
.B1(n_142),
.B2(n_145),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_554),
.B(n_571),
.Y(n_662)
);

OAI22x1_ASAP7_75t_L g663 ( 
.A1(n_514),
.A2(n_557),
.B1(n_588),
.B2(n_563),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_578),
.B(n_564),
.Y(n_664)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_531),
.A2(n_533),
.B(n_541),
.Y(n_665)
);

AOI22x1_ASAP7_75t_L g666 ( 
.A1(n_533),
.A2(n_551),
.B1(n_582),
.B2(n_562),
.Y(n_666)
);

AOI21xp5_ASAP7_75t_L g667 ( 
.A1(n_549),
.A2(n_585),
.B(n_575),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_553),
.A2(n_527),
.B1(n_594),
.B2(n_589),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_544),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_511),
.B(n_574),
.Y(n_670)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_572),
.A2(n_576),
.B(n_586),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g672 ( 
.A1(n_587),
.A2(n_600),
.B(n_590),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_551),
.B(n_529),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_577),
.A2(n_543),
.B(n_584),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_544),
.Y(n_675)
);

OAI22xp5_ASAP7_75t_L g676 ( 
.A1(n_588),
.A2(n_580),
.B1(n_597),
.B2(n_590),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_600),
.B(n_552),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_555),
.B(n_592),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_598),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_567),
.B(n_559),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_587),
.A2(n_390),
.B1(n_539),
.B2(n_602),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_596),
.B(n_495),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_530),
.A2(n_537),
.B(n_536),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_512),
.Y(n_684)
);

NOR2x1_ASAP7_75t_L g685 ( 
.A(n_601),
.B(n_414),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_650),
.Y(n_686)
);

AO21x1_ASAP7_75t_L g687 ( 
.A1(n_681),
.A2(n_619),
.B(n_656),
.Y(n_687)
);

AO21x1_ASAP7_75t_L g688 ( 
.A1(n_681),
.A2(n_619),
.B(n_656),
.Y(n_688)
);

INVx3_ASAP7_75t_SL g689 ( 
.A(n_640),
.Y(n_689)
);

AO31x2_ASAP7_75t_L g690 ( 
.A1(n_676),
.A2(n_668),
.A3(n_644),
.B(n_647),
.Y(n_690)
);

OA21x2_ASAP7_75t_L g691 ( 
.A1(n_672),
.A2(n_652),
.B(n_635),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_603),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_649),
.B(n_682),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_666),
.A2(n_665),
.B(n_614),
.Y(n_694)
);

AOI221xp5_ASAP7_75t_L g695 ( 
.A1(n_663),
.A2(n_610),
.B1(n_608),
.B2(n_637),
.C(n_645),
.Y(n_695)
);

BUFx8_ASAP7_75t_L g696 ( 
.A(n_617),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_627),
.B(n_625),
.Y(n_697)
);

AOI31xp67_ASAP7_75t_L g698 ( 
.A1(n_636),
.A2(n_638),
.A3(n_646),
.B(n_653),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_613),
.Y(n_699)
);

AO31x2_ASAP7_75t_L g700 ( 
.A1(n_671),
.A2(n_634),
.A3(n_642),
.B(n_674),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_685),
.B(n_607),
.Y(n_701)
);

NOR2x1_ASAP7_75t_L g702 ( 
.A(n_659),
.B(n_632),
.Y(n_702)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_628),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_662),
.Y(n_704)
);

AO32x2_ASAP7_75t_L g705 ( 
.A1(n_651),
.A2(n_629),
.A3(n_616),
.B1(n_661),
.B2(n_641),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_620),
.A2(n_621),
.B(n_667),
.C(n_618),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_607),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_623),
.A2(n_622),
.B1(n_677),
.B2(n_624),
.Y(n_708)
);

BUFx3_ASAP7_75t_L g709 ( 
.A(n_631),
.Y(n_709)
);

BUFx8_ASAP7_75t_L g710 ( 
.A(n_670),
.Y(n_710)
);

OAI22x1_ASAP7_75t_L g711 ( 
.A1(n_633),
.A2(n_670),
.B1(n_673),
.B2(n_660),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_626),
.A2(n_643),
.B1(n_679),
.B2(n_630),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_669),
.B(n_684),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_657),
.B(n_675),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_654),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_609),
.B(n_615),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_680),
.A2(n_678),
.B(n_655),
.Y(n_717)
);

AOI31xp67_ASAP7_75t_L g718 ( 
.A1(n_616),
.A2(n_636),
.A3(n_545),
.B(n_540),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_664),
.A2(n_596),
.B1(n_346),
.B2(n_345),
.Y(n_719)
);

AOI221x1_ASAP7_75t_L g720 ( 
.A1(n_604),
.A2(n_683),
.B1(n_681),
.B2(n_672),
.C(n_619),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_603),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_625),
.A2(n_510),
.B1(n_583),
.B2(n_596),
.Y(n_722)
);

BUFx3_ASAP7_75t_L g723 ( 
.A(n_640),
.Y(n_723)
);

AO31x2_ASAP7_75t_L g724 ( 
.A1(n_604),
.A2(n_683),
.A3(n_639),
.B(n_536),
.Y(n_724)
);

BUFx2_ASAP7_75t_R g725 ( 
.A(n_617),
.Y(n_725)
);

BUFx2_ASAP7_75t_L g726 ( 
.A(n_625),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_619),
.A2(n_625),
.B1(n_627),
.B2(n_612),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_604),
.A2(n_683),
.B(n_530),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_649),
.B(n_596),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_640),
.Y(n_730)
);

AO31x2_ASAP7_75t_L g731 ( 
.A1(n_604),
.A2(n_683),
.A3(n_639),
.B(n_536),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_637),
.Y(n_732)
);

OAI21xp5_ASAP7_75t_L g733 ( 
.A1(n_604),
.A2(n_683),
.B(n_536),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_603),
.B(n_596),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_603),
.A2(n_596),
.B1(n_346),
.B2(n_345),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_604),
.A2(n_683),
.A3(n_639),
.B(n_536),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_SL g737 ( 
.A(n_656),
.B(n_476),
.C(n_478),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_649),
.B(n_596),
.Y(n_738)
);

AOI221x1_ASAP7_75t_L g739 ( 
.A1(n_604),
.A2(n_683),
.B1(n_681),
.B2(n_672),
.C(n_619),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_640),
.Y(n_740)
);

OAI22x1_ASAP7_75t_L g741 ( 
.A1(n_685),
.A2(n_346),
.B1(n_345),
.B2(n_583),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_637),
.Y(n_742)
);

NOR2xp67_ASAP7_75t_L g743 ( 
.A(n_610),
.B(n_568),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_649),
.B(n_596),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_625),
.A2(n_510),
.B1(n_583),
.B2(n_596),
.Y(n_745)
);

AO31x2_ASAP7_75t_L g746 ( 
.A1(n_604),
.A2(n_683),
.A3(n_639),
.B(n_536),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_SL g747 ( 
.A(n_656),
.B(n_476),
.C(n_478),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_649),
.B(n_596),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_604),
.A2(n_683),
.B(n_536),
.Y(n_749)
);

AOI21xp5_ASAP7_75t_L g750 ( 
.A1(n_604),
.A2(n_683),
.B(n_530),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_637),
.Y(n_751)
);

AO32x2_ASAP7_75t_L g752 ( 
.A1(n_681),
.A2(n_619),
.A3(n_648),
.B1(n_676),
.B2(n_542),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_605),
.B(n_596),
.Y(n_753)
);

AOI221x1_ASAP7_75t_L g754 ( 
.A1(n_604),
.A2(n_683),
.B1(n_681),
.B2(n_672),
.C(n_619),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_640),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_649),
.B(n_596),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_605),
.B(n_596),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_604),
.A2(n_683),
.A3(n_639),
.B(n_536),
.Y(n_758)
);

AO32x2_ASAP7_75t_L g759 ( 
.A1(n_681),
.A2(n_619),
.A3(n_648),
.B1(n_676),
.B2(n_542),
.Y(n_759)
);

INVx1_ASAP7_75t_SL g760 ( 
.A(n_640),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_649),
.B(n_596),
.Y(n_761)
);

BUFx12f_ASAP7_75t_L g762 ( 
.A(n_631),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_649),
.B(n_596),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_604),
.A2(n_683),
.B(n_530),
.Y(n_764)
);

AOI21xp33_ASAP7_75t_L g765 ( 
.A1(n_603),
.A2(n_482),
.B(n_478),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_604),
.A2(n_683),
.B(n_530),
.Y(n_766)
);

OAI21xp5_ASAP7_75t_L g767 ( 
.A1(n_604),
.A2(n_683),
.B(n_536),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_603),
.B(n_596),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_610),
.B(n_568),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_649),
.B(n_596),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_619),
.A2(n_625),
.B1(n_627),
.B2(n_612),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_658),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_603),
.A2(n_596),
.B1(n_346),
.B2(n_345),
.Y(n_773)
);

AOI221xp5_ASAP7_75t_SL g774 ( 
.A1(n_606),
.A2(n_649),
.B1(n_611),
.B2(n_681),
.C(n_481),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_604),
.A2(n_683),
.B(n_532),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_649),
.B(n_596),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_685),
.B(n_547),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_603),
.A2(n_596),
.B1(n_346),
.B2(n_345),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_723),
.B(n_730),
.Y(n_779)
);

BUFx3_ASAP7_75t_L g780 ( 
.A(n_689),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_772),
.Y(n_781)
);

OR2x2_ASAP7_75t_L g782 ( 
.A(n_760),
.B(n_734),
.Y(n_782)
);

AO21x2_ASAP7_75t_L g783 ( 
.A1(n_687),
.A2(n_688),
.B(n_733),
.Y(n_783)
);

AO21x2_ASAP7_75t_L g784 ( 
.A1(n_749),
.A2(n_767),
.B(n_694),
.Y(n_784)
);

BUFx2_ASAP7_75t_L g785 ( 
.A(n_740),
.Y(n_785)
);

OA21x2_ASAP7_75t_L g786 ( 
.A1(n_720),
.A2(n_754),
.B(n_739),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_768),
.B(n_753),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_775),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_757),
.A2(n_692),
.B1(n_722),
.B2(n_745),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_SL g790 ( 
.A1(n_727),
.A2(n_771),
.B(n_747),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_696),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_697),
.B(n_735),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_755),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_732),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_774),
.A2(n_706),
.B(n_704),
.C(n_717),
.Y(n_795)
);

CKINVDCx16_ASAP7_75t_R g796 ( 
.A(n_762),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_704),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_693),
.B(n_729),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_738),
.A2(n_761),
.B(n_744),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_728),
.A2(n_766),
.A3(n_750),
.B(n_764),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_742),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_748),
.A2(n_756),
.B(n_770),
.C(n_763),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_695),
.A2(n_708),
.B1(n_776),
.B2(n_769),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_751),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_743),
.A2(n_737),
.B1(n_702),
.B2(n_726),
.Y(n_805)
);

OA21x2_ASAP7_75t_L g806 ( 
.A1(n_712),
.A2(n_718),
.B(n_752),
.Y(n_806)
);

AO31x2_ASAP7_75t_L g807 ( 
.A1(n_711),
.A2(n_752),
.A3(n_759),
.B(n_690),
.Y(n_807)
);

OA21x2_ASAP7_75t_L g808 ( 
.A1(n_752),
.A2(n_759),
.B(n_691),
.Y(n_808)
);

BUFx12f_ASAP7_75t_L g809 ( 
.A(n_703),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_696),
.Y(n_810)
);

CKINVDCx6p67_ASAP7_75t_R g811 ( 
.A(n_709),
.Y(n_811)
);

AO31x2_ASAP7_75t_L g812 ( 
.A1(n_759),
.A2(n_690),
.A3(n_716),
.B(n_736),
.Y(n_812)
);

OA21x2_ASAP7_75t_L g813 ( 
.A1(n_698),
.A2(n_690),
.B(n_705),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_710),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_715),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_721),
.B(n_707),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_710),
.A2(n_741),
.B1(n_765),
.B2(n_701),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_703),
.B(n_777),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_725),
.Y(n_819)
);

AO21x2_ASAP7_75t_L g820 ( 
.A1(n_705),
.A2(n_736),
.B(n_724),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_773),
.B(n_778),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_719),
.B(n_713),
.Y(n_822)
);

OAI21x1_ASAP7_75t_SL g823 ( 
.A1(n_699),
.A2(n_714),
.B(n_713),
.Y(n_823)
);

AO21x2_ASAP7_75t_L g824 ( 
.A1(n_705),
.A2(n_724),
.B(n_731),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_731),
.Y(n_825)
);

NAND2x1p5_ASAP7_75t_L g826 ( 
.A(n_746),
.B(n_758),
.Y(n_826)
);

OA21x2_ASAP7_75t_L g827 ( 
.A1(n_746),
.A2(n_739),
.B(n_720),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_700),
.B(n_596),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_SL g829 ( 
.A(n_703),
.B(n_547),
.Y(n_829)
);

BUFx12f_ASAP7_75t_L g830 ( 
.A(n_762),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_689),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_727),
.A2(n_656),
.B1(n_633),
.B2(n_771),
.Y(n_832)
);

INVx1_ASAP7_75t_SL g833 ( 
.A(n_689),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_686),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_802),
.B(n_798),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_788),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_828),
.B(n_797),
.Y(n_837)
);

OR2x2_ASAP7_75t_SL g838 ( 
.A(n_806),
.B(n_786),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_781),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_795),
.B(n_781),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_802),
.B(n_798),
.Y(n_841)
);

OAI222xp33_ASAP7_75t_L g842 ( 
.A1(n_832),
.A2(n_803),
.B1(n_789),
.B2(n_821),
.C1(n_817),
.C2(n_805),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_812),
.B(n_826),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_812),
.B(n_826),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_794),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_801),
.Y(n_846)
);

BUFx3_ASAP7_75t_L g847 ( 
.A(n_823),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_804),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_793),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_803),
.A2(n_792),
.B1(n_787),
.B2(n_799),
.Y(n_850)
);

AO21x2_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_784),
.B(n_824),
.Y(n_851)
);

INVxp67_ASAP7_75t_L g852 ( 
.A(n_782),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_812),
.B(n_827),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_790),
.B(n_825),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_800),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_800),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_800),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_827),
.B(n_807),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_834),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_807),
.B(n_820),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_836),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_859),
.B(n_843),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_855),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_837),
.B(n_786),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_854),
.B(n_784),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_855),
.Y(n_867)
);

NOR2x1_ASAP7_75t_R g868 ( 
.A(n_847),
.B(n_819),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_844),
.B(n_813),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_850),
.A2(n_817),
.B1(n_822),
.B2(n_805),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_853),
.B(n_808),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_835),
.B(n_841),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_839),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_853),
.B(n_808),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_874),
.B(n_861),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_864),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_866),
.B(n_856),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_865),
.B(n_838),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_872),
.B(n_841),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_874),
.B(n_861),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_862),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_874),
.B(n_861),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_874),
.B(n_857),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_869),
.B(n_856),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_869),
.B(n_871),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_869),
.B(n_851),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_871),
.B(n_851),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_877),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_887),
.B(n_872),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_878),
.B(n_865),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_885),
.B(n_875),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_887),
.B(n_871),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_885),
.B(n_875),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_883),
.Y(n_894)
);

INVx2_ASAP7_75t_SL g895 ( 
.A(n_884),
.Y(n_895)
);

OR2x2_ASAP7_75t_L g896 ( 
.A(n_878),
.B(n_865),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_876),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_887),
.B(n_867),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_885),
.B(n_863),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_881),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_875),
.B(n_863),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_880),
.B(n_863),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_900),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_894),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_891),
.B(n_886),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_888),
.B(n_883),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_895),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_889),
.B(n_842),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_900),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_897),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_898),
.A2(n_868),
.B(n_842),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_889),
.B(n_879),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_890),
.B(n_880),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_898),
.B(n_882),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_899),
.B(n_882),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_897),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_899),
.B(n_882),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_890),
.A2(n_870),
.B1(n_879),
.B2(n_850),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_903),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_905),
.B(n_891),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_912),
.B(n_893),
.Y(n_921)
);

NOR3xp33_ASAP7_75t_L g922 ( 
.A(n_911),
.B(n_908),
.C(n_796),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_912),
.B(n_830),
.Y(n_923)
);

OAI211xp5_ASAP7_75t_SL g924 ( 
.A1(n_918),
.A2(n_870),
.B(n_833),
.C(n_852),
.Y(n_924)
);

INVxp33_ASAP7_75t_L g925 ( 
.A(n_907),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_908),
.A2(n_895),
.B1(n_886),
.B2(n_902),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_910),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_916),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_903),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_909),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_905),
.B(n_893),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_909),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_906),
.Y(n_933)
);

OAI322xp33_ASAP7_75t_SL g934 ( 
.A1(n_921),
.A2(n_917),
.A3(n_915),
.B1(n_914),
.B2(n_892),
.C1(n_904),
.C2(n_819),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_SL g935 ( 
.A1(n_922),
.A2(n_926),
.B1(n_923),
.B2(n_933),
.C(n_896),
.Y(n_935)
);

AOI221xp5_ASAP7_75t_L g936 ( 
.A1(n_926),
.A2(n_906),
.B1(n_901),
.B2(n_902),
.C(n_892),
.Y(n_936)
);

OAI322xp33_ASAP7_75t_SL g937 ( 
.A1(n_927),
.A2(n_845),
.A3(n_846),
.B1(n_848),
.B2(n_913),
.C1(n_858),
.C2(n_860),
.Y(n_937)
);

NAND3xp33_ASAP7_75t_SL g938 ( 
.A(n_925),
.B(n_831),
.C(n_814),
.Y(n_938)
);

AOI21xp33_ASAP7_75t_SL g939 ( 
.A1(n_933),
.A2(n_810),
.B(n_791),
.Y(n_939)
);

AOI222xp33_ASAP7_75t_SL g940 ( 
.A1(n_924),
.A2(n_852),
.B1(n_830),
.B2(n_811),
.C1(n_888),
.C2(n_849),
.Y(n_940)
);

NAND4xp25_ASAP7_75t_SL g941 ( 
.A(n_939),
.B(n_920),
.C(n_931),
.D(n_901),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_938),
.A2(n_868),
.B(n_933),
.Y(n_942)
);

AOI321xp33_ASAP7_75t_L g943 ( 
.A1(n_935),
.A2(n_906),
.A3(n_920),
.B1(n_931),
.B2(n_896),
.C(n_886),
.Y(n_943)
);

INVx2_ASAP7_75t_SL g944 ( 
.A(n_934),
.Y(n_944)
);

AOI211xp5_ASAP7_75t_SL g945 ( 
.A1(n_937),
.A2(n_868),
.B(n_840),
.C(n_873),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_940),
.A2(n_927),
.B1(n_928),
.B2(n_888),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_945),
.B(n_944),
.Y(n_947)
);

AOI221xp5_ASAP7_75t_L g948 ( 
.A1(n_941),
.A2(n_936),
.B1(n_928),
.B2(n_929),
.C(n_930),
.Y(n_948)
);

NAND4xp25_ASAP7_75t_L g949 ( 
.A(n_943),
.B(n_942),
.C(n_946),
.D(n_780),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_945),
.B(n_929),
.Y(n_950)
);

NAND5xp2_ASAP7_75t_L g951 ( 
.A(n_947),
.B(n_829),
.C(n_779),
.D(n_809),
.E(n_840),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_949),
.B(n_950),
.C(n_948),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_947),
.B(n_780),
.C(n_785),
.Y(n_953)
);

NAND4xp75_ASAP7_75t_L g954 ( 
.A(n_947),
.B(n_809),
.C(n_840),
.D(n_816),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_954),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_953),
.B(n_919),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_955),
.B(n_952),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_956),
.B(n_818),
.Y(n_958)
);

INVx5_ASAP7_75t_L g959 ( 
.A(n_957),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_SL g960 ( 
.A1(n_959),
.A2(n_957),
.B1(n_958),
.B2(n_818),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_960),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_961),
.A2(n_959),
.B(n_951),
.Y(n_962)
);

INVxp67_ASAP7_75t_L g963 ( 
.A(n_962),
.Y(n_963)
);

AOI22xp33_ASAP7_75t_L g964 ( 
.A1(n_963),
.A2(n_959),
.B1(n_956),
.B2(n_932),
.Y(n_964)
);


endmodule