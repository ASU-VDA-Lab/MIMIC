module fake_jpeg_291_n_206 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_206);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_47),
.B(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_55),
.Y(n_84)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_49),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_48),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_54),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_49),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_51),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_53),
.B1(n_68),
.B2(n_65),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_88),
.B1(n_51),
.B2(n_57),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_57),
.B1(n_65),
.B2(n_68),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_76),
.B(n_73),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_50),
.B(n_63),
.Y(n_114)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_77),
.A2(n_58),
.B1(n_62),
.B2(n_75),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_106),
.B1(n_50),
.B2(n_75),
.Y(n_108)
);

INVx5_ASAP7_75t_SL g98 ( 
.A(n_85),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_71),
.B1(n_1),
.B2(n_2),
.Y(n_121)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_105),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_59),
.C(n_56),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_60),
.C(n_52),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_59),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_60),
.B1(n_52),
.B2(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_89),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_110),
.B1(n_121),
.B2(n_101),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_126),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_62),
.B1(n_58),
.B2(n_54),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_96),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_61),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_5),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_90),
.A2(n_89),
.B1(n_71),
.B2(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_45),
.C(n_41),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_35),
.C(n_34),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_0),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_125),
.B(n_127),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_5),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_128),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_132),
.B1(n_137),
.B2(n_145),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_121),
.A2(n_99),
.B1(n_107),
.B2(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_135),
.Y(n_150)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_6),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_138),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_140),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_23),
.B(n_39),
.C(n_36),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_122),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_141),
.B(n_142),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_120),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_22),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_40),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_123),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_154),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_126),
.C(n_33),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_161),
.C(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_153),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_159),
.Y(n_180)
);

NAND2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_8),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_29),
.C(n_28),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_21),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_27),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_26),
.C(n_25),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_9),
.Y(n_177)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_24),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_168),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_179),
.Y(n_187)
);

AOI21xp33_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_140),
.B(n_12),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_161),
.B(n_155),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_172),
.B(n_177),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_173),
.Y(n_185)
);

AOI322xp5_ASAP7_75t_SL g176 ( 
.A1(n_152),
.A2(n_156),
.A3(n_163),
.B1(n_155),
.B2(n_151),
.C1(n_164),
.C2(n_167),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_176),
.B(n_181),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_178),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_182),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g184 ( 
.A(n_169),
.B(n_158),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_172),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_175),
.A2(n_12),
.B(n_13),
.Y(n_190)
);

AOI31xp67_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_191),
.A3(n_182),
.B(n_16),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_13),
.C(n_14),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_180),
.B1(n_171),
.B2(n_174),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_195),
.B1(n_188),
.B2(n_191),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_186),
.B(n_189),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_197),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_177),
.B(n_16),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_198),
.A2(n_194),
.B1(n_17),
.B2(n_18),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_202),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_203),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_200),
.B(n_15),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_19),
.Y(n_206)
);


endmodule