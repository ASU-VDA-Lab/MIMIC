module real_jpeg_30135_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_0),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_0),
.A2(n_26),
.B1(n_30),
.B2(n_108),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_0),
.A2(n_52),
.B1(n_53),
.B2(n_108),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_0),
.A2(n_57),
.B1(n_59),
.B2(n_108),
.Y(n_242)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_1),
.Y(n_93)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_36),
.B1(n_57),
.B2(n_59),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_36),
.B1(n_52),
.B2(n_53),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_3),
.A2(n_24),
.B1(n_52),
.B2(n_53),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_3),
.A2(n_24),
.B1(n_26),
.B2(n_30),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_3),
.A2(n_24),
.B1(n_57),
.B2(n_59),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_5),
.A2(n_47),
.B1(n_52),
.B2(n_53),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_5),
.A2(n_47),
.B1(n_57),
.B2(n_59),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_5),
.A2(n_26),
.B1(n_30),
.B2(n_47),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_7),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_7),
.A2(n_26),
.B1(n_30),
.B2(n_169),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_7),
.A2(n_52),
.B1(n_53),
.B2(n_169),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_7),
.A2(n_57),
.B1(n_59),
.B2(n_169),
.Y(n_255)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_9),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_9),
.B(n_25),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_9),
.B(n_30),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_30),
.B(n_207),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_167),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_9),
.A2(n_54),
.B(n_57),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_9),
.B(n_74),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_9),
.A2(n_93),
.B1(n_112),
.B2(n_255),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_10),
.A2(n_22),
.B1(n_23),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_10),
.A2(n_45),
.B1(n_52),
.B2(n_53),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_10),
.A2(n_26),
.B1(n_30),
.B2(n_45),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_10),
.A2(n_45),
.B1(n_57),
.B2(n_59),
.Y(n_182)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_12),
.A2(n_22),
.B1(n_23),
.B2(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_12),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_12),
.A2(n_26),
.B1(n_30),
.B2(n_134),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_134),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_12),
.A2(n_57),
.B1(n_59),
.B2(n_134),
.Y(n_247)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_14),
.A2(n_52),
.B1(n_53),
.B2(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_14),
.A2(n_26),
.B1(n_30),
.B2(n_65),
.Y(n_70)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_14),
.Y(n_206)
);

INVx11_ASAP7_75t_SL g58 ( 
.A(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_81),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_79),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_37),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_31),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_20),
.A2(n_43),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_21),
.A2(n_32),
.B(n_78),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_28),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_28),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g166 ( 
.A(n_22),
.B(n_167),
.CON(n_166),
.SN(n_166)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_25),
.A2(n_32),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_26),
.A2(n_33),
.B1(n_166),
.B2(n_180),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g203 ( 
.A1(n_26),
.A2(n_52),
.A3(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_28),
.B(n_30),
.Y(n_180)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_31),
.A2(n_44),
.B(n_48),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_32),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_80),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_71),
.C(n_76),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_39),
.A2(n_40),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_49),
.C(n_62),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_41),
.A2(n_42),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_43),
.A2(n_48),
.B1(n_107),
.B2(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_43),
.A2(n_48),
.B1(n_133),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_49),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_49),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_49),
.A2(n_62),
.B1(n_307),
.B2(n_321),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_56),
.B(n_60),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_56),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_50),
.A2(n_100),
.B(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_50),
.A2(n_60),
.B(n_116),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_50),
.A2(n_56),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_50),
.A2(n_140),
.B(n_215),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_50),
.A2(n_56),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_50),
.A2(n_56),
.B1(n_214),
.B2(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_53),
.B(n_205),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g233 ( 
.A1(n_53),
.A2(n_55),
.B(n_167),
.C(n_234),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_56)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_99),
.B(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_56),
.B(n_167),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_57),
.Y(n_59)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_59),
.B(n_260),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_61),
.B(n_118),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_62),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_63),
.A2(n_73),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_68),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_64),
.A2(n_69),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_64),
.A2(n_69),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_64),
.A2(n_69),
.B1(n_163),
.B2(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_64),
.A2(n_69),
.B1(n_191),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_74),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_71),
.A2(n_72),
.B1(n_76),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_73),
.A2(n_74),
.B(n_75),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_73),
.A2(n_75),
.B(n_130),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_73),
.A2(n_130),
.B(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_76),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_332),
.B(n_338),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_302),
.A3(n_324),
.B1(n_330),
.B2(n_331),
.C(n_340),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_152),
.B(n_301),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_135),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_85),
.B(n_135),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_109),
.C(n_120),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_86),
.A2(n_87),
.B1(n_109),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_103),
.C(n_105),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_98),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_89),
.B(n_98),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_90),
.A2(n_113),
.B(n_182),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_91),
.A2(n_97),
.B(n_125),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_91),
.A2(n_92),
.B1(n_246),
.B2(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_97),
.Y(n_96)
);

INVx11_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_93),
.A2(n_112),
.B1(n_123),
.B2(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_113),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_96),
.A2(n_112),
.B(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_97),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_104),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_109),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_119),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_111),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_115),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_111),
.A2(n_146),
.B(n_149),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_112),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_112),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_128),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_120),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_129),
.C(n_131),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_121),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_126),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_129),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_150),
.B2(n_151),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_138),
.B(n_145),
.C(n_151),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_141),
.B(n_144),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_143),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_144),
.B(n_304),
.C(n_314),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_144),
.A2(n_304),
.B1(n_305),
.B2(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_144),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_295),
.B(n_300),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_195),
.B(n_281),
.C(n_294),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_183),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_155),
.B(n_183),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_170),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_157),
.B(n_158),
.C(n_170),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_165),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_167),
.B(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_168),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_189),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_184),
.A2(n_185),
.B1(n_276),
.B2(n_278),
.Y(n_275)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_189),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_194),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_280),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_273),
.B(n_279),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_225),
.B(n_272),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_216),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_199),
.B(n_216),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_209),
.C(n_212),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_200),
.A2(n_201),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_203),
.Y(n_223)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_210),
.B1(n_212),
.B2(n_213),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_221),
.B2(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_223),
.C(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_266),
.B(n_271),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_243),
.B(n_265),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_235),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_228),
.B(n_235),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_230),
.B1(n_233),
.B2(n_250),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_233),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_251),
.B(n_264),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_245),
.B(n_249),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_257),
.B(n_263),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_274),
.B(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_282),
.B(n_283),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_284),
.A2(n_285),
.B1(n_292),
.B2(n_293),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_292),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_316),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_316),
.Y(n_331)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_305)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_309),
.C(n_311),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.B1(n_318),
.B2(n_322),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_322),
.C(n_323),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_315),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_323),
.Y(n_316)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule