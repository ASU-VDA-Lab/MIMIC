module fake_jpeg_3327_n_199 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_199);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_199;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_5),
.B(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVxp33_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx10_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_14),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_7),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_69),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_22),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_52),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_48),
.B1(n_47),
.B2(n_45),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_50),
.B1(n_65),
.B2(n_58),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g77 ( 
.A(n_61),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_70),
.Y(n_83)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_50),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_81),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_83),
.Y(n_112)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_86),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_74),
.A2(n_50),
.B1(n_65),
.B2(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_89),
.B(n_93),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_56),
.C(n_53),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_59),
.C(n_56),
.Y(n_110)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_91),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_57),
.Y(n_92)
);

OR2x2_ASAP7_75t_SL g94 ( 
.A(n_84),
.B(n_75),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_73),
.B1(n_76),
.B2(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_95),
.A2(n_83),
.B1(n_85),
.B2(n_81),
.Y(n_115)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g117 ( 
.A(n_99),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_79),
.B(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_101),
.B(n_1),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_89),
.B(n_66),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_63),
.C(n_51),
.Y(n_130)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_65),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_60),
.Y(n_121)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_108),
.B(n_83),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_109),
.A2(n_81),
.B1(n_90),
.B2(n_85),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_118),
.B1(n_95),
.B2(n_97),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_44),
.B1(n_43),
.B2(n_42),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_93),
.B(n_68),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_116),
.A2(n_100),
.B(n_99),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_64),
.B1(n_55),
.B2(n_78),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_41),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_123),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_94),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_4),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_5),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_117),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_111),
.C(n_106),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_136),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_116),
.B(n_103),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_38),
.B(n_37),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_129),
.Y(n_142)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_114),
.A2(n_110),
.B1(n_100),
.B2(n_107),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_26),
.B1(n_25),
.B2(n_28),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_51),
.B(n_63),
.C(n_24),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_121),
.B(n_122),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_149),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_119),
.B(n_23),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_147),
.B(n_153),
.C(n_154),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_8),
.B1(n_12),
.B2(n_13),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g149 ( 
.A(n_120),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_6),
.B(n_7),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_151),
.A2(n_128),
.B(n_10),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_128),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_152),
.B(n_16),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_40),
.C(n_39),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_170),
.B1(n_171),
.B2(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_155),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_133),
.B(n_146),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_137),
.A2(n_8),
.B(n_11),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_166),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_167),
.B(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_35),
.C(n_32),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_15),
.C(n_16),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_160),
.A2(n_138),
.B1(n_143),
.B2(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_177),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_165),
.B1(n_157),
.B2(n_170),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_171),
.Y(n_181)
);

OAI322xp33_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_145),
.A3(n_169),
.B1(n_162),
.B2(n_159),
.C1(n_157),
.C2(n_172),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_185),
.B(n_178),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_156),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_184),
.B(n_187),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_161),
.B(n_164),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_178),
.B(n_174),
.Y(n_189)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_192),
.C(n_186),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_191),
.A2(n_184),
.B(n_190),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_183),
.B(n_176),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_168),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_176),
.B(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_197),
.A2(n_17),
.A3(n_18),
.B1(n_19),
.B2(n_20),
.C1(n_196),
.C2(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_17),
.Y(n_199)
);


endmodule