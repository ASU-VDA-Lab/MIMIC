module fake_netlist_1_7993_n_1517 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_331, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1517);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_331;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1517;
wire n_1309;
wire n_1497;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1477;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1503;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1475;
wire n_1505;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1500;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_641;
wire n_379;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_822;
wire n_706;
wire n_823;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1499;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1510;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_1502;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1361;
wire n_1333;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1488;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_1468;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_1515;
wire n_897;
wire n_1188;
wire n_1496;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_1472;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_1514;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_1060;
wire n_721;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_1490;
wire n_867;
wire n_1070;
wire n_1270;
wire n_1474;
wire n_1512;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1507;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_1495;
wire n_606;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_1483;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1513;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_659;
wire n_432;
wire n_1329;
wire n_1509;
wire n_1185;
wire n_1511;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1508;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_1480;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_805;
wire n_729;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_1470;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1471;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_1473;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1478;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_1492;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_1489;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1516;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_1493;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1498;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_1501;
wire n_777;
wire n_1504;
wire n_351;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1479;
wire n_1360;
wire n_1486;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_1481;
wire n_798;
wire n_887;
wire n_471;
wire n_1476;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1491;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1485;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1482;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_1494;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_1506;
wire n_1469;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1484;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_445;
wire n_398;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_1487;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_819;
wire n_772;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g348 ( .A(n_102), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_188), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_345), .Y(n_350) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_77), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_61), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_202), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_323), .Y(n_354) );
BUFx2_ASAP7_75t_SL g355 ( .A(n_63), .Y(n_355) );
INVxp67_ASAP7_75t_L g356 ( .A(n_240), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_160), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_66), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_31), .B(n_179), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
CKINVDCx20_ASAP7_75t_R g361 ( .A(n_209), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_36), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_26), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_312), .B(n_200), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_220), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_118), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_4), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_159), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_22), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_12), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_19), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_186), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_265), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_327), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_151), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_147), .Y(n_376) );
CKINVDCx20_ASAP7_75t_R g377 ( .A(n_100), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_181), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_258), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_218), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_9), .Y(n_381) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_40), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_141), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_252), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_57), .Y(n_385) );
CKINVDCx5p33_ASAP7_75t_R g386 ( .A(n_342), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_42), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_76), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_170), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_68), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_50), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_290), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g394 ( .A(n_340), .Y(n_394) );
CKINVDCx14_ASAP7_75t_R g395 ( .A(n_231), .Y(n_395) );
INVxp33_ASAP7_75t_SL g396 ( .A(n_245), .Y(n_396) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_162), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_92), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_332), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_29), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_296), .Y(n_401) );
INVxp67_ASAP7_75t_L g402 ( .A(n_140), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_214), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_262), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_62), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_45), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_22), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_292), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_76), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_343), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_228), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_331), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_308), .Y(n_413) );
BUFx3_ASAP7_75t_L g414 ( .A(n_47), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_40), .Y(n_415) );
INVx2_ASAP7_75t_SL g416 ( .A(n_157), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_148), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_78), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_11), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_326), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_158), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_180), .Y(n_422) );
BUFx5_ASAP7_75t_L g423 ( .A(n_68), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_61), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_48), .Y(n_425) );
INVxp67_ASAP7_75t_SL g426 ( .A(n_208), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_125), .Y(n_427) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_96), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_301), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_203), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_72), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_167), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_289), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_45), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_196), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_310), .Y(n_436) );
CKINVDCx5p33_ASAP7_75t_R g437 ( .A(n_324), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_337), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_111), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_172), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_169), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_109), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g443 ( .A(n_201), .B(n_63), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_14), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_250), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_100), .Y(n_446) );
BUFx2_ASAP7_75t_SL g447 ( .A(n_269), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_293), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_318), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_42), .Y(n_450) );
BUFx3_ASAP7_75t_L g451 ( .A(n_234), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_53), .Y(n_452) );
INVxp33_ASAP7_75t_L g453 ( .A(n_119), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_316), .Y(n_454) );
CKINVDCx14_ASAP7_75t_R g455 ( .A(n_210), .Y(n_455) );
CKINVDCx14_ASAP7_75t_R g456 ( .A(n_69), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_216), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_38), .B(n_338), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_168), .Y(n_459) );
XOR2xp5_ASAP7_75t_L g460 ( .A(n_103), .B(n_50), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_5), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_256), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_212), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g464 ( .A(n_153), .Y(n_464) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_317), .Y(n_465) );
BUFx2_ASAP7_75t_SL g466 ( .A(n_103), .Y(n_466) );
CKINVDCx16_ASAP7_75t_R g467 ( .A(n_55), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_206), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_144), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_11), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_88), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_58), .Y(n_472) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_133), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_112), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_268), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_164), .Y(n_476) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_44), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_60), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_65), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_261), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_270), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_46), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_184), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_46), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_287), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_74), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_155), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_242), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_276), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_185), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_58), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_300), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_211), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_9), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_314), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_85), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_47), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_222), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_173), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_330), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_37), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_255), .Y(n_502) );
BUFx3_ASAP7_75t_L g503 ( .A(n_7), .Y(n_503) );
INVx2_ASAP7_75t_SL g504 ( .A(n_166), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_138), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_31), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_23), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_277), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_283), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_295), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_66), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_236), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_266), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_219), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_82), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_251), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_263), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_232), .Y(n_518) );
INVxp33_ASAP7_75t_SL g519 ( .A(n_150), .Y(n_519) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_285), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_335), .Y(n_521) );
BUFx10_ASAP7_75t_L g522 ( .A(n_152), .Y(n_522) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_225), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_92), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_416), .B(n_0), .Y(n_525) );
NOR2xp33_ASAP7_75t_R g526 ( .A(n_395), .B(n_113), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_400), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_400), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_423), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_408), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_451), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_408), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_400), .B(n_0), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_423), .Y(n_534) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_408), .Y(n_535) );
INVx4_ASAP7_75t_L g536 ( .A(n_522), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_397), .B(n_1), .Y(n_537) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_408), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_363), .B(n_1), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_394), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_423), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_456), .Y(n_542) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_490), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_456), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_363), .B(n_2), .Y(n_545) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_374), .A2(n_115), .B(n_114), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_423), .Y(n_547) );
INVx6_ASAP7_75t_L g548 ( .A(n_522), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_420), .B(n_2), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_423), .Y(n_550) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_352), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_551) );
NAND2xp33_ASAP7_75t_L g552 ( .A(n_423), .B(n_347), .Y(n_552) );
BUFx8_ASAP7_75t_L g553 ( .A(n_423), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_453), .B(n_3), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_385), .B(n_6), .Y(n_555) );
INVx4_ASAP7_75t_L g556 ( .A(n_522), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_362), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_504), .B(n_467), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_385), .B(n_6), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_361), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_362), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_387), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_387), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_409), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_367), .B(n_7), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_542), .B(n_453), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_536), .B(n_370), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_542), .B(n_395), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_536), .B(n_356), .Y(n_569) );
AO22x2_ASAP7_75t_L g570 ( .A1(n_533), .A2(n_460), .B1(n_466), .B2(n_355), .Y(n_570) );
INVx4_ASAP7_75t_L g571 ( .A(n_533), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_533), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_536), .B(n_370), .Y(n_573) );
OR2x2_ASAP7_75t_SL g574 ( .A(n_558), .B(n_359), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_536), .B(n_368), .Y(n_575) );
AND2x6_ASAP7_75t_L g576 ( .A(n_533), .B(n_451), .Y(n_576) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_530), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_556), .B(n_391), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_556), .B(n_455), .Y(n_579) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_556), .Y(n_580) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_556), .B(n_402), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_553), .B(n_378), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_553), .B(n_378), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_529), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_553), .B(n_461), .C(n_391), .Y(n_585) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_539), .B(n_458), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_529), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_548), .B(n_470), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_539), .B(n_364), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_541), .Y(n_590) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_548), .B(n_493), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_548), .B(n_470), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_541), .Y(n_593) );
BUFx2_ASAP7_75t_L g594 ( .A(n_553), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_539), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_554), .A2(n_396), .B1(n_519), .B2(n_491), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_539), .B(n_414), .Y(n_597) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_530), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_545), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_554), .Y(n_601) );
AO22x2_ASAP7_75t_L g602 ( .A1(n_545), .A2(n_477), .B1(n_428), .B2(n_418), .Y(n_602) );
BUFx3_ASAP7_75t_L g603 ( .A(n_531), .Y(n_603) );
INVx4_ASAP7_75t_L g604 ( .A(n_545), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_555), .Y(n_605) );
NAND2xp33_ASAP7_75t_L g606 ( .A(n_526), .B(n_490), .Y(n_606) );
BUFx2_ASAP7_75t_L g607 ( .A(n_544), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g608 ( .A(n_540), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_548), .B(n_455), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_534), .Y(n_610) );
AND2x6_ASAP7_75t_L g611 ( .A(n_555), .B(n_349), .Y(n_611) );
CKINVDCx16_ASAP7_75t_R g612 ( .A(n_555), .Y(n_612) );
INVx4_ASAP7_75t_L g613 ( .A(n_555), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
OR2x6_ASAP7_75t_L g615 ( .A(n_570), .B(n_559), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_567), .B(n_537), .Y(n_616) );
INVx4_ASAP7_75t_L g617 ( .A(n_594), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_580), .B(n_549), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_602), .A2(n_611), .B1(n_586), .B2(n_599), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_603), .Y(n_620) );
AND2x4_ASAP7_75t_L g621 ( .A(n_594), .B(n_559), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_608), .Y(n_622) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_611), .Y(n_623) );
INVx2_ASAP7_75t_SL g624 ( .A(n_568), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g625 ( .A(n_612), .B(n_559), .Y(n_625) );
INVx2_ASAP7_75t_SL g626 ( .A(n_568), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_566), .B(n_531), .Y(n_627) );
AND2x4_ASAP7_75t_L g628 ( .A(n_601), .B(n_559), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_608), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_571), .B(n_547), .Y(n_630) );
INVx3_ASAP7_75t_L g631 ( .A(n_571), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_603), .Y(n_632) );
INVx2_ASAP7_75t_SL g633 ( .A(n_566), .Y(n_633) );
AOI22xp5_ASAP7_75t_L g634 ( .A1(n_586), .A2(n_525), .B1(n_441), .B2(n_459), .Y(n_634) );
INVx2_ASAP7_75t_SL g635 ( .A(n_609), .Y(n_635) );
AND2x4_ASAP7_75t_L g636 ( .A(n_601), .B(n_565), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g637 ( .A(n_571), .B(n_547), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_579), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_579), .B(n_531), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_573), .B(n_527), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_604), .B(n_550), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_578), .B(n_527), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_602), .Y(n_644) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_611), .Y(n_645) );
NAND3xp33_ASAP7_75t_L g646 ( .A(n_596), .B(n_552), .C(n_551), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_602), .Y(n_647) );
AOI22xp33_ASAP7_75t_L g648 ( .A1(n_611), .A2(n_550), .B1(n_528), .B2(n_557), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_611), .A2(n_441), .B1(n_459), .B2(n_361), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_609), .B(n_464), .Y(n_650) );
NOR3xp33_ASAP7_75t_SL g651 ( .A(n_585), .B(n_560), .C(n_491), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g652 ( .A(n_607), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_604), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_589), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g655 ( .A(n_607), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g656 ( .A(n_613), .B(n_350), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_588), .B(n_464), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_569), .B(n_528), .Y(n_658) );
AND2x6_ASAP7_75t_SL g659 ( .A(n_592), .B(n_348), .Y(n_659) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_589), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_613), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_575), .B(n_386), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_597), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_589), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_613), .B(n_499), .Y(n_665) );
BUFx3_ASAP7_75t_L g666 ( .A(n_576), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_597), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_572), .B(n_353), .Y(n_668) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_576), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_595), .B(n_354), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_597), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_600), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_605), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_576), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_576), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_581), .B(n_386), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_591), .B(n_393), .Y(n_677) );
INVx4_ASAP7_75t_L g678 ( .A(n_576), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_610), .B(n_357), .Y(n_679) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_610), .B(n_360), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_611), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_576), .A2(n_561), .B1(n_562), .B2(n_557), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_574), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_574), .Y(n_684) );
BUFx3_ASAP7_75t_L g685 ( .A(n_584), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_582), .B(n_393), .Y(n_686) );
BUFx2_ASAP7_75t_R g687 ( .A(n_583), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_614), .B(n_436), .Y(n_688) );
OR2x6_ASAP7_75t_L g689 ( .A(n_570), .B(n_447), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_614), .B(n_436), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_590), .B(n_437), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_570), .B(n_499), .C(n_369), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_590), .Y(n_693) );
OAI22xp5_ASAP7_75t_SL g694 ( .A1(n_570), .A2(n_352), .B1(n_377), .B2(n_369), .Y(n_694) );
BUFx2_ASAP7_75t_L g695 ( .A(n_593), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_593), .Y(n_696) );
INVx4_ASAP7_75t_L g697 ( .A(n_587), .Y(n_697) );
AO22x1_ASAP7_75t_L g698 ( .A1(n_587), .A2(n_396), .B1(n_519), .B2(n_439), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_606), .A2(n_546), .B(n_376), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_577), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_577), .B(n_564), .Y(n_701) );
NAND2xp5_ASAP7_75t_SL g702 ( .A(n_577), .B(n_365), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_577), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_577), .B(n_437), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_598), .B(n_439), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_598), .B(n_469), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_598), .B(n_561), .Y(n_707) );
AOI21xp5_ASAP7_75t_L g708 ( .A1(n_630), .A2(n_546), .B(n_445), .Y(n_708) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_623), .Y(n_709) );
INVx4_ASAP7_75t_L g710 ( .A(n_617), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_636), .B(n_351), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_695), .Y(n_712) );
BUFx3_ASAP7_75t_L g713 ( .A(n_652), .Y(n_713) );
INVx4_ASAP7_75t_L g714 ( .A(n_617), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_667), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_671), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_630), .A2(n_546), .B(n_465), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_685), .Y(n_718) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_637), .A2(n_546), .B(n_523), .Y(n_719) );
OAI22xp5_ASAP7_75t_SL g720 ( .A1(n_694), .A2(n_407), .B1(n_377), .B2(n_415), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_636), .B(n_407), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_633), .B(n_515), .Y(n_722) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_623), .Y(n_723) );
INVx3_ASAP7_75t_L g724 ( .A(n_685), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_619), .A2(n_473), .B1(n_475), .B2(n_469), .Y(n_725) );
AO21x1_ASAP7_75t_L g726 ( .A1(n_699), .A2(n_372), .B(n_366), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_619), .A2(n_475), .B1(n_483), .B2(n_473), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_628), .B(n_483), .Y(n_728) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_644), .A2(n_492), .B1(n_488), .B2(n_371), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_622), .Y(n_730) );
AND2x4_ASAP7_75t_L g731 ( .A(n_624), .B(n_358), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_638), .B(n_488), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_657), .B(n_414), .Y(n_733) );
NAND2x1p5_ASAP7_75t_L g734 ( .A(n_664), .B(n_503), .Y(n_734) );
INVxp67_ASAP7_75t_L g735 ( .A(n_665), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_638), .B(n_492), .Y(n_736) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_623), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_653), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_683), .B(n_381), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_637), .A2(n_426), .B(n_375), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_616), .B(n_618), .Y(n_741) );
BUFx12f_ASAP7_75t_L g742 ( .A(n_629), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_663), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_616), .B(n_627), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g745 ( .A(n_684), .B(n_388), .Y(n_745) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_644), .A2(n_398), .B1(n_405), .B2(n_392), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_657), .B(n_503), .Y(n_747) );
BUFx2_ASAP7_75t_L g748 ( .A(n_665), .Y(n_748) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_615), .A2(n_419), .B1(n_424), .B2(n_406), .Y(n_749) );
BUFx6f_ASAP7_75t_L g750 ( .A(n_623), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_654), .Y(n_751) );
AND2x4_ASAP7_75t_L g752 ( .A(n_626), .B(n_442), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_641), .A2(n_446), .B(n_450), .C(n_444), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g754 ( .A(n_655), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_672), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_654), .A2(n_471), .B1(n_472), .B2(n_452), .Y(n_756) );
BUFx3_ASAP7_75t_L g757 ( .A(n_615), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_661), .Y(n_758) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_642), .A2(n_379), .B(n_373), .Y(n_759) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_660), .Y(n_760) );
A2O1A1Ixp33_ASAP7_75t_L g761 ( .A1(n_673), .A2(n_478), .B(n_482), .C(n_479), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g762 ( .A(n_660), .B(n_484), .Y(n_762) );
O2A1O1Ixp33_ASAP7_75t_L g763 ( .A1(n_647), .A2(n_494), .B(n_496), .C(n_486), .Y(n_763) );
A2O1A1Ixp33_ASAP7_75t_SL g764 ( .A1(n_682), .A2(n_563), .B(n_564), .C(n_562), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_693), .Y(n_765) );
INVx3_ASAP7_75t_L g766 ( .A(n_697), .Y(n_766) );
OR2x6_ASAP7_75t_L g767 ( .A(n_689), .B(n_409), .Y(n_767) );
INVx2_ASAP7_75t_L g768 ( .A(n_631), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_634), .A2(n_506), .B1(n_507), .B2(n_501), .C(n_497), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g770 ( .A(n_650), .B(n_511), .Y(n_770) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_645), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_642), .A2(n_383), .B(n_380), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_621), .B(n_524), .Y(n_773) );
O2A1O1Ixp33_ASAP7_75t_L g774 ( .A1(n_625), .A2(n_425), .B(n_431), .C(n_418), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_696), .Y(n_775) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_692), .A2(n_646), .B1(n_650), .B2(n_625), .C(n_635), .Y(n_776) );
OAI21xp33_ASAP7_75t_SL g777 ( .A1(n_615), .A2(n_563), .B(n_443), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_640), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_621), .B(n_425), .Y(n_779) );
NOR2x1_ASAP7_75t_L g780 ( .A(n_666), .B(n_678), .Y(n_780) );
BUFx6f_ASAP7_75t_L g781 ( .A(n_645), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g782 ( .A1(n_649), .A2(n_431), .B1(n_434), .B2(n_382), .Y(n_782) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_689), .Y(n_783) );
OR2x6_ASAP7_75t_SL g784 ( .A(n_687), .B(n_401), .Y(n_784) );
HB1xp67_ASAP7_75t_L g785 ( .A(n_689), .Y(n_785) );
INVx1_ASAP7_75t_SL g786 ( .A(n_645), .Y(n_786) );
INVx2_ASAP7_75t_SL g787 ( .A(n_698), .Y(n_787) );
INVx3_ASAP7_75t_L g788 ( .A(n_631), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_643), .Y(n_789) );
BUFx6f_ASAP7_75t_L g790 ( .A(n_645), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g791 ( .A1(n_656), .A2(n_389), .B(n_384), .Y(n_791) );
BUFx2_ASAP7_75t_L g792 ( .A(n_659), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_670), .Y(n_793) );
INVx5_ASAP7_75t_L g794 ( .A(n_678), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_668), .Y(n_795) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_666), .Y(n_796) );
A2O1A1Ixp33_ASAP7_75t_L g797 ( .A1(n_658), .A2(n_434), .B(n_399), .C(n_403), .Y(n_797) );
INVx3_ASAP7_75t_L g798 ( .A(n_620), .Y(n_798) );
AOI21xp5_ASAP7_75t_L g799 ( .A1(n_656), .A2(n_410), .B(n_390), .Y(n_799) );
AOI21x1_ASAP7_75t_L g800 ( .A1(n_702), .A2(n_412), .B(n_411), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g801 ( .A1(n_639), .A2(n_417), .B(n_413), .Y(n_801) );
NOR3xp33_ASAP7_75t_L g802 ( .A(n_686), .B(n_480), .C(n_422), .Y(n_802) );
AOI21xp5_ASAP7_75t_L g803 ( .A1(n_688), .A2(n_427), .B(n_421), .Y(n_803) );
BUFx2_ASAP7_75t_L g804 ( .A(n_669), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g805 ( .A1(n_681), .A2(n_382), .B1(n_430), .B2(n_429), .Y(n_805) );
O2A1O1Ixp33_ASAP7_75t_L g806 ( .A1(n_679), .A2(n_435), .B(n_438), .C(n_432), .Y(n_806) );
INVx2_ASAP7_75t_L g807 ( .A(n_701), .Y(n_807) );
BUFx6f_ASAP7_75t_L g808 ( .A(n_701), .Y(n_808) );
INVx4_ASAP7_75t_L g809 ( .A(n_669), .Y(n_809) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_707), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_707), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g812 ( .A1(n_690), .A2(n_457), .B(n_454), .Y(n_812) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_651), .Y(n_813) );
O2A1O1Ixp33_ASAP7_75t_L g814 ( .A1(n_679), .A2(n_463), .B(n_468), .C(n_462), .Y(n_814) );
INVx3_ASAP7_75t_L g815 ( .A(n_632), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_682), .A2(n_476), .B1(n_481), .B2(n_474), .Y(n_816) );
INVx1_ASAP7_75t_SL g817 ( .A(n_691), .Y(n_817) );
OR2x2_ASAP7_75t_L g818 ( .A(n_677), .B(n_8), .Y(n_818) );
OR2x6_ASAP7_75t_L g819 ( .A(n_681), .B(n_382), .Y(n_819) );
BUFx2_ASAP7_75t_L g820 ( .A(n_651), .Y(n_820) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_703), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g822 ( .A1(n_674), .A2(n_487), .B(n_485), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_648), .B(n_404), .Y(n_823) );
OAI21xp33_ASAP7_75t_L g824 ( .A1(n_648), .A2(n_495), .B(n_489), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_704), .Y(n_825) );
OAI21xp33_ASAP7_75t_L g826 ( .A1(n_662), .A2(n_676), .B(n_680), .Y(n_826) );
INVx2_ASAP7_75t_SL g827 ( .A(n_680), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_705), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_706), .Y(n_829) );
AOI21xp5_ASAP7_75t_L g830 ( .A1(n_675), .A2(n_505), .B(n_500), .Y(n_830) );
OR2x6_ASAP7_75t_L g831 ( .A(n_702), .B(n_382), .Y(n_831) );
AND2x2_ASAP7_75t_L g832 ( .A(n_703), .B(n_8), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_700), .B(n_433), .Y(n_833) );
NOR2xp33_ASAP7_75t_L g834 ( .A(n_703), .B(n_440), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_703), .A2(n_510), .B(n_508), .Y(n_835) );
INVx3_ASAP7_75t_L g836 ( .A(n_617), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_633), .B(n_448), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_636), .B(n_513), .Y(n_838) );
INVx1_ASAP7_75t_SL g839 ( .A(n_654), .Y(n_839) );
OR2x2_ASAP7_75t_L g840 ( .A(n_622), .B(n_10), .Y(n_840) );
INVx1_ASAP7_75t_SL g841 ( .A(n_654), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_633), .B(n_514), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_685), .Y(n_843) );
NOR2xp33_ASAP7_75t_R g844 ( .A(n_622), .B(n_10), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_695), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_695), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_665), .Y(n_847) );
OAI21x1_ASAP7_75t_L g848 ( .A1(n_708), .A2(n_376), .B(n_374), .Y(n_848) );
NAND2x1p5_ASAP7_75t_L g849 ( .A(n_710), .B(n_516), .Y(n_849) );
INVx2_ASAP7_75t_SL g850 ( .A(n_713), .Y(n_850) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_839), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_821), .Y(n_852) );
INVx2_ASAP7_75t_L g853 ( .A(n_821), .Y(n_853) );
BUFx2_ASAP7_75t_L g854 ( .A(n_841), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_712), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_726), .A2(n_498), .B(n_449), .Y(n_856) );
OAI21x1_ASAP7_75t_L g857 ( .A1(n_717), .A2(n_498), .B(n_449), .Y(n_857) );
OAI21x1_ASAP7_75t_L g858 ( .A1(n_719), .A2(n_509), .B(n_502), .Y(n_858) );
OAI21x1_ASAP7_75t_L g859 ( .A1(n_800), .A2(n_509), .B(n_502), .Y(n_859) );
OAI21x1_ASAP7_75t_L g860 ( .A1(n_835), .A2(n_518), .B(n_512), .Y(n_860) );
NAND2xp5_ASAP7_75t_SL g861 ( .A(n_709), .B(n_517), .Y(n_861) );
OAI21x1_ASAP7_75t_L g862 ( .A1(n_822), .A2(n_518), .B(n_512), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_778), .A2(n_521), .B1(n_520), .B2(n_490), .Y(n_863) );
OA21x2_ASAP7_75t_L g864 ( .A1(n_826), .A2(n_520), .B(n_490), .Y(n_864) );
AND2x4_ASAP7_75t_L g865 ( .A(n_789), .B(n_12), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_741), .B(n_13), .Y(n_866) );
INVx1_ASAP7_75t_L g867 ( .A(n_845), .Y(n_867) );
OAI21x1_ASAP7_75t_L g868 ( .A1(n_825), .A2(n_520), .B(n_117), .Y(n_868) );
BUFx2_ASAP7_75t_R g869 ( .A(n_784), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_821), .Y(n_870) );
OR2x6_ASAP7_75t_L g871 ( .A(n_710), .B(n_520), .Y(n_871) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_841), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g873 ( .A1(n_749), .A2(n_532), .B1(n_535), .B2(n_530), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g874 ( .A1(n_744), .A2(n_532), .B1(n_535), .B2(n_530), .Y(n_874) );
OAI21x1_ASAP7_75t_L g875 ( .A1(n_830), .A2(n_120), .B(n_116), .Y(n_875) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_751), .Y(n_876) );
OR2x2_ASAP7_75t_L g877 ( .A(n_721), .B(n_13), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_846), .Y(n_878) );
AND2x4_ASAP7_75t_L g879 ( .A(n_714), .B(n_14), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_776), .A2(n_532), .B1(n_535), .B2(n_530), .Y(n_880) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_828), .A2(n_122), .B(n_121), .Y(n_881) );
AO21x2_ASAP7_75t_L g882 ( .A1(n_826), .A2(n_535), .B(n_532), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_760), .B(n_15), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_755), .Y(n_884) );
OAI21x1_ASAP7_75t_SL g885 ( .A1(n_714), .A2(n_15), .B(n_16), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g886 ( .A(n_742), .Y(n_886) );
AO21x2_ASAP7_75t_L g887 ( .A1(n_764), .A2(n_535), .B(n_532), .Y(n_887) );
OAI21x1_ASAP7_75t_L g888 ( .A1(n_832), .A2(n_124), .B(n_123), .Y(n_888) );
INVx2_ASAP7_75t_L g889 ( .A(n_765), .Y(n_889) );
OR2x6_ASAP7_75t_L g890 ( .A(n_767), .B(n_16), .Y(n_890) );
AO21x2_ASAP7_75t_L g891 ( .A1(n_797), .A2(n_543), .B(n_538), .Y(n_891) );
OAI21x1_ASAP7_75t_L g892 ( .A1(n_801), .A2(n_127), .B(n_126), .Y(n_892) );
OAI21x1_ASAP7_75t_L g893 ( .A1(n_803), .A2(n_129), .B(n_128), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_775), .Y(n_894) );
OR2x6_ASAP7_75t_L g895 ( .A(n_767), .B(n_757), .Y(n_895) );
INVx3_ASAP7_75t_L g896 ( .A(n_766), .Y(n_896) );
INVx2_ASAP7_75t_L g897 ( .A(n_709), .Y(n_897) );
INVx2_ASAP7_75t_L g898 ( .A(n_709), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_817), .B(n_17), .Y(n_899) );
AND2x2_ASAP7_75t_L g900 ( .A(n_748), .B(n_17), .Y(n_900) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_829), .A2(n_543), .B(n_538), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_767), .A2(n_543), .B1(n_538), .B2(n_598), .Y(n_902) );
NAND2x1p5_ASAP7_75t_L g903 ( .A(n_836), .B(n_538), .Y(n_903) );
OR2x6_ASAP7_75t_L g904 ( .A(n_819), .B(n_18), .Y(n_904) );
INVx1_ASAP7_75t_L g905 ( .A(n_779), .Y(n_905) );
NAND2x1p5_ASAP7_75t_L g906 ( .A(n_836), .B(n_538), .Y(n_906) );
O2A1O1Ixp33_ASAP7_75t_SL g907 ( .A1(n_783), .A2(n_131), .B(n_132), .C(n_130), .Y(n_907) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_833), .A2(n_598), .B(n_543), .Y(n_908) );
OAI21x1_ASAP7_75t_L g909 ( .A1(n_812), .A2(n_135), .B(n_134), .Y(n_909) );
INVx2_ASAP7_75t_SL g910 ( .A(n_734), .Y(n_910) );
OAI21x1_ASAP7_75t_L g911 ( .A1(n_759), .A2(n_137), .B(n_136), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_817), .B(n_18), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_746), .B(n_19), .Y(n_913) );
BUFx8_ASAP7_75t_SL g914 ( .A(n_754), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_723), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_743), .Y(n_916) );
INVx6_ASAP7_75t_L g917 ( .A(n_808), .Y(n_917) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_723), .Y(n_918) );
OAI21x1_ASAP7_75t_L g919 ( .A1(n_798), .A2(n_815), .B(n_780), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_723), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_731), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_746), .B(n_20), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_731), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_815), .A2(n_142), .B(n_139), .Y(n_924) );
INVx1_ASAP7_75t_L g925 ( .A(n_752), .Y(n_925) );
AND2x2_ASAP7_75t_L g926 ( .A(n_847), .B(n_20), .Y(n_926) );
INVx1_ASAP7_75t_L g927 ( .A(n_752), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_737), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_838), .B(n_21), .Y(n_929) );
INVx2_ASAP7_75t_SL g930 ( .A(n_730), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_715), .Y(n_931) );
OR2x2_ASAP7_75t_L g932 ( .A(n_711), .B(n_21), .Y(n_932) );
INVx1_ASAP7_75t_L g933 ( .A(n_716), .Y(n_933) );
INVx2_ASAP7_75t_L g934 ( .A(n_737), .Y(n_934) );
NOR2xp67_ASAP7_75t_L g935 ( .A(n_777), .B(n_24), .Y(n_935) );
OR2x6_ASAP7_75t_L g936 ( .A(n_819), .B(n_24), .Y(n_936) );
AO21x2_ASAP7_75t_L g937 ( .A1(n_749), .A2(n_543), .B(n_143), .Y(n_937) );
OA21x2_ASAP7_75t_L g938 ( .A1(n_824), .A2(n_146), .B(n_145), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_737), .Y(n_939) );
O2A1O1Ixp33_ASAP7_75t_SL g940 ( .A1(n_785), .A2(n_191), .B(n_341), .C(n_339), .Y(n_940) );
O2A1O1Ixp33_ASAP7_75t_L g941 ( .A1(n_761), .A2(n_25), .B(n_26), .C(n_27), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_735), .B(n_25), .Y(n_942) );
OR2x2_ASAP7_75t_L g943 ( .A(n_720), .B(n_27), .Y(n_943) );
AO31x2_ASAP7_75t_L g944 ( .A1(n_739), .A2(n_28), .A3(n_29), .B(n_30), .Y(n_944) );
OA21x2_ASAP7_75t_L g945 ( .A1(n_824), .A2(n_154), .B(n_149), .Y(n_945) );
OAI21x1_ASAP7_75t_L g946 ( .A1(n_780), .A2(n_161), .B(n_156), .Y(n_946) );
CKINVDCx16_ASAP7_75t_R g947 ( .A(n_844), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_733), .Y(n_948) );
BUFx6f_ASAP7_75t_L g949 ( .A(n_750), .Y(n_949) );
AND2x4_ASAP7_75t_L g950 ( .A(n_794), .B(n_28), .Y(n_950) );
BUFx8_ASAP7_75t_L g951 ( .A(n_792), .Y(n_951) );
INVx2_ASAP7_75t_L g952 ( .A(n_750), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_747), .Y(n_953) );
INVx3_ASAP7_75t_L g954 ( .A(n_766), .Y(n_954) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_773), .B(n_30), .Y(n_955) );
BUFx2_ASAP7_75t_SL g956 ( .A(n_794), .Y(n_956) );
BUFx2_ASAP7_75t_SL g957 ( .A(n_794), .Y(n_957) );
OAI21x1_ASAP7_75t_L g958 ( .A1(n_772), .A2(n_165), .B(n_163), .Y(n_958) );
AO21x2_ASAP7_75t_L g959 ( .A1(n_791), .A2(n_174), .B(n_171), .Y(n_959) );
NOR2x1p5_ASAP7_75t_L g960 ( .A(n_840), .B(n_32), .Y(n_960) );
OAI21xp5_ASAP7_75t_L g961 ( .A1(n_793), .A2(n_176), .B(n_175), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_795), .Y(n_962) );
OA21x2_ASAP7_75t_L g963 ( .A1(n_799), .A2(n_178), .B(n_177), .Y(n_963) );
OA21x2_ASAP7_75t_L g964 ( .A1(n_740), .A2(n_183), .B(n_182), .Y(n_964) );
A2O1A1Ixp33_ASAP7_75t_L g965 ( .A1(n_777), .A2(n_32), .B(n_33), .C(n_34), .Y(n_965) );
AND2x2_ASAP7_75t_L g966 ( .A(n_722), .B(n_33), .Y(n_966) );
OAI21x1_ASAP7_75t_L g967 ( .A1(n_774), .A2(n_189), .B(n_187), .Y(n_967) );
OAI21x1_ASAP7_75t_L g968 ( .A1(n_724), .A2(n_192), .B(n_190), .Y(n_968) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_724), .Y(n_969) );
OAI21x1_ASAP7_75t_L g970 ( .A1(n_806), .A2(n_194), .B(n_193), .Y(n_970) );
NOR2x1_ASAP7_75t_R g971 ( .A(n_820), .B(n_34), .Y(n_971) );
OAI221xp5_ASAP7_75t_L g972 ( .A1(n_769), .A2(n_35), .B1(n_36), .B2(n_37), .C(n_38), .Y(n_972) );
OAI21x1_ASAP7_75t_L g973 ( .A1(n_814), .A2(n_197), .B(n_195), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_782), .A2(n_35), .B1(n_39), .B2(n_41), .Y(n_974) );
BUFx6f_ASAP7_75t_L g975 ( .A(n_750), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_818), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_816), .A2(n_819), .B1(n_787), .B2(n_718), .Y(n_977) );
OAI21xp5_ASAP7_75t_L g978 ( .A1(n_827), .A2(n_199), .B(n_198), .Y(n_978) );
HB1xp67_ASAP7_75t_L g979 ( .A(n_804), .Y(n_979) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_843), .Y(n_980) );
OAI21x1_ASAP7_75t_L g981 ( .A1(n_753), .A2(n_205), .B(n_204), .Y(n_981) );
AOI21xp33_ASAP7_75t_L g982 ( .A1(n_770), .A2(n_39), .B(n_41), .Y(n_982) );
AO32x2_ASAP7_75t_L g983 ( .A1(n_729), .A2(n_43), .A3(n_44), .B1(n_48), .B2(n_49), .Y(n_983) );
AOI221xp5_ASAP7_75t_L g984 ( .A1(n_756), .A2(n_43), .B1(n_49), .B2(n_51), .C(n_52), .Y(n_984) );
OAI21x1_ASAP7_75t_L g985 ( .A1(n_788), .A2(n_805), .B(n_768), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_762), .B(n_51), .Y(n_986) );
AOI21xp5_ASAP7_75t_L g987 ( .A1(n_823), .A2(n_230), .B(n_336), .Y(n_987) );
INVx2_ASAP7_75t_L g988 ( .A(n_771), .Y(n_988) );
NOR2x1_ASAP7_75t_R g989 ( .A(n_720), .B(n_52), .Y(n_989) );
INVx5_ASAP7_75t_L g990 ( .A(n_771), .Y(n_990) );
OR2x6_ASAP7_75t_L g991 ( .A(n_831), .B(n_771), .Y(n_991) );
OAI21x1_ASAP7_75t_L g992 ( .A1(n_788), .A2(n_229), .B(n_334), .Y(n_992) );
BUFx2_ASAP7_75t_L g993 ( .A(n_808), .Y(n_993) );
BUFx3_ASAP7_75t_L g994 ( .A(n_781), .Y(n_994) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_763), .A2(n_53), .B(n_54), .C(n_55), .Y(n_995) );
A2O1A1Ixp33_ASAP7_75t_L g996 ( .A1(n_745), .A2(n_54), .B(n_56), .C(n_57), .Y(n_996) );
OA21x2_ASAP7_75t_L g997 ( .A1(n_816), .A2(n_235), .B(n_333), .Y(n_997) );
AND2x4_ASAP7_75t_L g998 ( .A(n_809), .B(n_56), .Y(n_998) );
AO21x2_ASAP7_75t_L g999 ( .A1(n_802), .A2(n_237), .B(n_329), .Y(n_999) );
AOI21xp33_ASAP7_75t_L g1000 ( .A1(n_837), .A2(n_59), .B(n_60), .Y(n_1000) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_842), .A2(n_59), .B1(n_62), .B2(n_64), .Y(n_1001) );
BUFx3_ASAP7_75t_L g1002 ( .A(n_781), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_807), .Y(n_1003) );
BUFx6f_ASAP7_75t_L g1004 ( .A(n_781), .Y(n_1004) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_813), .Y(n_1005) );
BUFx10_ASAP7_75t_L g1006 ( .A(n_808), .Y(n_1006) );
OAI21x1_ASAP7_75t_L g1007 ( .A1(n_738), .A2(n_233), .B(n_325), .Y(n_1007) );
OAI21x1_ASAP7_75t_SL g1008 ( .A1(n_809), .A2(n_64), .B(n_65), .Y(n_1008) );
BUFx3_ASAP7_75t_L g1009 ( .A(n_914), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1010 ( .A1(n_865), .A2(n_725), .B1(n_727), .B2(n_732), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1011 ( .A1(n_908), .A2(n_786), .B(n_834), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_889), .Y(n_1012) );
OAI21x1_ASAP7_75t_L g1013 ( .A1(n_857), .A2(n_758), .B(n_811), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1014 ( .A1(n_865), .A2(n_831), .B1(n_736), .B2(n_786), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_865), .A2(n_728), .B1(n_810), .B2(n_831), .Y(n_1015) );
BUFx6f_ASAP7_75t_L g1016 ( .A(n_918), .Y(n_1016) );
OAI22xp5_ASAP7_75t_L g1017 ( .A1(n_890), .A2(n_810), .B1(n_796), .B2(n_790), .Y(n_1017) );
OR2x2_ASAP7_75t_L g1018 ( .A(n_854), .B(n_810), .Y(n_1018) );
AO31x2_ASAP7_75t_L g1019 ( .A1(n_965), .A2(n_790), .A3(n_69), .B(n_70), .Y(n_1019) );
INVx2_ASAP7_75t_L g1020 ( .A(n_889), .Y(n_1020) );
OAI22xp5_ASAP7_75t_L g1021 ( .A1(n_890), .A2(n_796), .B1(n_790), .B2(n_71), .Y(n_1021) );
AOI222xp33_ASAP7_75t_L g1022 ( .A1(n_989), .A2(n_796), .B1(n_70), .B2(n_71), .C1(n_72), .C2(n_73), .Y(n_1022) );
AOI22xp33_ASAP7_75t_L g1023 ( .A1(n_890), .A2(n_67), .B1(n_73), .B2(n_74), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_855), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g1025 ( .A1(n_904), .A2(n_67), .B1(n_75), .B2(n_77), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_904), .A2(n_75), .B1(n_78), .B2(n_79), .Y(n_1026) );
CKINVDCx16_ASAP7_75t_R g1027 ( .A(n_947), .Y(n_1027) );
INVx2_ASAP7_75t_L g1028 ( .A(n_894), .Y(n_1028) );
OAI22xp5_ASAP7_75t_SL g1029 ( .A1(n_943), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_851), .B(n_80), .Y(n_1030) );
CKINVDCx6p67_ASAP7_75t_R g1031 ( .A(n_904), .Y(n_1031) );
OAI31xp33_ASAP7_75t_L g1032 ( .A1(n_972), .A2(n_81), .A3(n_82), .B(n_83), .Y(n_1032) );
AOI222xp33_ASAP7_75t_L g1033 ( .A1(n_971), .A2(n_83), .B1(n_84), .B2(n_85), .C1(n_86), .C2(n_87), .Y(n_1033) );
NAND2xp5_ASAP7_75t_L g1034 ( .A(n_851), .B(n_84), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_872), .B(n_866), .Y(n_1035) );
OAI221xp5_ASAP7_75t_L g1036 ( .A1(n_976), .A2(n_86), .B1(n_87), .B2(n_88), .C(n_89), .Y(n_1036) );
AOI22xp33_ASAP7_75t_SL g1037 ( .A1(n_879), .A2(n_89), .B1(n_90), .B2(n_91), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_894), .Y(n_1038) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_936), .A2(n_90), .B1(n_91), .B2(n_93), .Y(n_1039) );
OAI21xp33_ASAP7_75t_SL g1040 ( .A1(n_936), .A2(n_93), .B(n_94), .Y(n_1040) );
OAI21x1_ASAP7_75t_L g1041 ( .A1(n_857), .A2(n_259), .B(n_322), .Y(n_1041) );
OAI222xp33_ASAP7_75t_L g1042 ( .A1(n_936), .A2(n_94), .B1(n_95), .B2(n_96), .C1(n_97), .C2(n_98), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_872), .B(n_95), .Y(n_1043) );
O2A1O1Ixp33_ASAP7_75t_L g1044 ( .A1(n_965), .A2(n_97), .B(n_98), .C(n_99), .Y(n_1044) );
OAI22xp5_ASAP7_75t_L g1045 ( .A1(n_977), .A2(n_99), .B1(n_101), .B2(n_102), .Y(n_1045) );
INVx1_ASAP7_75t_L g1046 ( .A(n_867), .Y(n_1046) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_948), .A2(n_101), .B1(n_104), .B2(n_105), .C(n_106), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1048 ( .A1(n_895), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_1048) );
INVx1_ASAP7_75t_L g1049 ( .A(n_878), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_876), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_884), .B(n_107), .Y(n_1051) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_953), .A2(n_107), .B1(n_108), .B2(n_109), .C(n_110), .Y(n_1052) );
OAI22xp33_ASAP7_75t_L g1053 ( .A1(n_895), .A2(n_108), .B1(n_110), .B2(n_207), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1054 ( .A(n_905), .B(n_921), .Y(n_1054) );
AO31x2_ASAP7_75t_L g1055 ( .A1(n_874), .A2(n_213), .A3(n_215), .B(n_217), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_916), .Y(n_1056) );
OA21x2_ASAP7_75t_L g1057 ( .A1(n_858), .A2(n_221), .B(n_223), .Y(n_1057) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_923), .A2(n_224), .B1(n_226), .B2(n_227), .C(n_238), .Y(n_1058) );
NOR2xp33_ASAP7_75t_L g1059 ( .A(n_877), .B(n_239), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1060 ( .A(n_914), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_925), .B(n_346), .Y(n_1061) );
OAI222xp33_ASAP7_75t_L g1062 ( .A1(n_1001), .A2(n_241), .B1(n_243), .B2(n_244), .C1(n_246), .C2(n_247), .Y(n_1062) );
INVx1_ASAP7_75t_L g1063 ( .A(n_931), .Y(n_1063) );
OAI21x1_ASAP7_75t_L g1064 ( .A1(n_858), .A2(n_248), .B(n_249), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_960), .A2(n_253), .B1(n_254), .B2(n_257), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_879), .A2(n_260), .B1(n_264), .B2(n_267), .Y(n_1066) );
OAI211xp5_ASAP7_75t_L g1067 ( .A1(n_1001), .A2(n_271), .B(n_272), .C(n_273), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1068 ( .A(n_895), .B(n_274), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_927), .B(n_321), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1070 ( .A1(n_998), .A2(n_275), .B1(n_278), .B2(n_279), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_933), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_966), .B(n_320), .Y(n_1072) );
INVx1_ASAP7_75t_L g1073 ( .A(n_962), .Y(n_1073) );
O2A1O1Ixp33_ASAP7_75t_L g1074 ( .A1(n_1000), .A2(n_280), .B(n_281), .C(n_282), .Y(n_1074) );
AOI21xp5_ASAP7_75t_L g1075 ( .A1(n_848), .A2(n_284), .B(n_286), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_979), .B(n_876), .Y(n_1076) );
AOI21xp5_ASAP7_75t_L g1077 ( .A1(n_901), .A2(n_288), .B(n_291), .Y(n_1077) );
AOI21xp5_ASAP7_75t_L g1078 ( .A1(n_856), .A2(n_294), .B(n_297), .Y(n_1078) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1003), .Y(n_1079) );
AOI21xp5_ASAP7_75t_L g1080 ( .A1(n_856), .A2(n_298), .B(n_299), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_979), .B(n_302), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_871), .Y(n_1082) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_932), .A2(n_303), .B1(n_304), .B2(n_305), .C(n_306), .Y(n_1083) );
A2O1A1Ixp33_ASAP7_75t_L g1084 ( .A1(n_935), .A2(n_307), .B(n_309), .C(n_311), .Y(n_1084) );
OAI211xp5_ASAP7_75t_L g1085 ( .A1(n_984), .A2(n_313), .B(n_315), .C(n_319), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_879), .A2(n_986), .B1(n_922), .B2(n_913), .Y(n_1086) );
AOI21xp5_ASAP7_75t_L g1087 ( .A1(n_882), .A2(n_861), .B(n_859), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_900), .B(n_926), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_998), .A2(n_899), .B1(n_912), .B2(n_950), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1090 ( .A1(n_871), .A2(n_849), .B1(n_991), .B2(n_998), .Y(n_1090) );
AOI21xp5_ASAP7_75t_L g1091 ( .A1(n_882), .A2(n_861), .B(n_859), .Y(n_1091) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_871), .A2(n_849), .B1(n_991), .B2(n_929), .Y(n_1092) );
OA21x2_ASAP7_75t_L g1093 ( .A1(n_868), .A2(n_985), .B(n_888), .Y(n_1093) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_942), .A2(n_955), .B1(n_995), .B2(n_883), .C(n_850), .Y(n_1094) );
INVx3_ASAP7_75t_L g1095 ( .A(n_991), .Y(n_1095) );
INVx1_ASAP7_75t_L g1096 ( .A(n_944), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1097 ( .A1(n_950), .A2(n_930), .B1(n_982), .B2(n_1005), .Y(n_1097) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_950), .A2(n_1005), .B1(n_980), .B2(n_910), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_980), .A2(n_974), .B1(n_993), .B2(n_917), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_974), .A2(n_996), .B1(n_969), .B2(n_880), .Y(n_1100) );
INVx2_ASAP7_75t_SL g1101 ( .A(n_1006), .Y(n_1101) );
OAI211xp5_ASAP7_75t_L g1102 ( .A1(n_996), .A2(n_941), .B(n_863), .C(n_880), .Y(n_1102) );
INVx1_ASAP7_75t_L g1103 ( .A(n_944), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_944), .Y(n_1104) );
AOI222xp33_ASAP7_75t_L g1105 ( .A1(n_951), .A2(n_869), .B1(n_885), .B2(n_1008), .C1(n_886), .C2(n_969), .Y(n_1105) );
AOI221xp5_ASAP7_75t_L g1106 ( .A1(n_873), .A2(n_863), .B1(n_886), .B2(n_907), .C(n_940), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1107 ( .A(n_1006), .B(n_983), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1108 ( .A1(n_997), .A2(n_873), .B1(n_902), .B2(n_978), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_944), .Y(n_1109) );
INVx2_ASAP7_75t_L g1110 ( .A(n_891), .Y(n_1110) );
NOR2x1_ASAP7_75t_SL g1111 ( .A(n_956), .B(n_957), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1112 ( .A1(n_907), .A2(n_940), .B1(n_896), .B2(n_954), .C(n_987), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_951), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1114 ( .A1(n_917), .A2(n_951), .B1(n_896), .B2(n_954), .Y(n_1114) );
BUFx5_ASAP7_75t_L g1115 ( .A(n_994), .Y(n_1115) );
AND2x4_ASAP7_75t_L g1116 ( .A(n_990), .B(n_1002), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1117 ( .A1(n_864), .A2(n_887), .B(n_853), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_917), .A2(n_891), .B1(n_999), .B2(n_997), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_983), .B(n_903), .Y(n_1119) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_983), .B(n_903), .Y(n_1120) );
OAI22xp5_ASAP7_75t_L g1121 ( .A1(n_902), .A2(n_997), .B1(n_906), .B2(n_990), .Y(n_1121) );
OA21x2_ASAP7_75t_L g1122 ( .A1(n_888), .A2(n_862), .B(n_860), .Y(n_1122) );
NAND3xp33_ASAP7_75t_L g1123 ( .A(n_961), .B(n_964), .C(n_963), .Y(n_1123) );
OR2x4_ASAP7_75t_L g1124 ( .A(n_918), .B(n_975), .Y(n_1124) );
INVx6_ASAP7_75t_L g1125 ( .A(n_990), .Y(n_1125) );
AOI21xp5_ASAP7_75t_L g1126 ( .A1(n_864), .A2(n_887), .B(n_853), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_906), .B(n_919), .Y(n_1127) );
INVx2_ASAP7_75t_L g1128 ( .A(n_860), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1129 ( .A1(n_964), .A2(n_963), .B1(n_938), .B2(n_945), .C(n_928), .Y(n_1129) );
INVx1_ASAP7_75t_L g1130 ( .A(n_983), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1131 ( .A1(n_990), .A2(n_945), .B1(n_938), .B2(n_1002), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_981), .A2(n_999), .B1(n_937), .B2(n_973), .Y(n_1132) );
INVx1_ASAP7_75t_L g1133 ( .A(n_893), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1134 ( .A1(n_864), .A2(n_852), .B(n_870), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_981), .B(n_937), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_862), .B(n_920), .Y(n_1136) );
INVx2_ASAP7_75t_L g1137 ( .A(n_911), .Y(n_1137) );
AOI21xp5_ASAP7_75t_L g1138 ( .A1(n_852), .A2(n_870), .B(n_988), .Y(n_1138) );
INVxp67_ASAP7_75t_SL g1139 ( .A(n_918), .Y(n_1139) );
AOI22xp33_ASAP7_75t_SL g1140 ( .A1(n_970), .A2(n_973), .B1(n_893), .B2(n_909), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1141 ( .A1(n_994), .A2(n_949), .B1(n_1004), .B2(n_918), .Y(n_1141) );
OAI211xp5_ASAP7_75t_L g1142 ( .A1(n_909), .A2(n_892), .B(n_946), .C(n_958), .Y(n_1142) );
OAI22xp33_ASAP7_75t_L g1143 ( .A1(n_949), .A2(n_975), .B1(n_1004), .B2(n_915), .Y(n_1143) );
OAI22xp5_ASAP7_75t_L g1144 ( .A1(n_949), .A2(n_975), .B1(n_1004), .B2(n_915), .Y(n_1144) );
O2A1O1Ixp33_ASAP7_75t_L g1145 ( .A1(n_959), .A2(n_952), .B(n_988), .C(n_928), .Y(n_1145) );
BUFx12f_ASAP7_75t_L g1146 ( .A(n_949), .Y(n_1146) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_975), .A2(n_1004), .B1(n_952), .B2(n_897), .Y(n_1147) );
AOI21xp5_ASAP7_75t_L g1148 ( .A1(n_897), .A2(n_920), .B(n_939), .Y(n_1148) );
INVx2_ASAP7_75t_L g1149 ( .A(n_911), .Y(n_1149) );
A2O1A1Ixp33_ASAP7_75t_L g1150 ( .A1(n_970), .A2(n_967), .B(n_892), .C(n_875), .Y(n_1150) );
AOI222xp33_ASAP7_75t_L g1151 ( .A1(n_875), .A2(n_898), .B1(n_934), .B2(n_939), .C1(n_958), .C2(n_967), .Y(n_1151) );
OAI211xp5_ASAP7_75t_L g1152 ( .A1(n_881), .A2(n_992), .B(n_968), .C(n_924), .Y(n_1152) );
AOI22xp33_ASAP7_75t_L g1153 ( .A1(n_959), .A2(n_898), .B1(n_934), .B2(n_1007), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_855), .Y(n_1154) );
AOI21xp5_ASAP7_75t_L g1155 ( .A1(n_908), .A2(n_717), .B(n_708), .Y(n_1155) );
AOI21xp5_ASAP7_75t_L g1156 ( .A1(n_908), .A2(n_717), .B(n_708), .Y(n_1156) );
OR2x6_ASAP7_75t_L g1157 ( .A(n_890), .B(n_904), .Y(n_1157) );
AOI21xp5_ASAP7_75t_L g1158 ( .A1(n_908), .A2(n_717), .B(n_708), .Y(n_1158) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_865), .A2(n_767), .B1(n_890), .B2(n_619), .Y(n_1159) );
INVx2_ASAP7_75t_L g1160 ( .A(n_1012), .Y(n_1160) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1157), .B(n_1020), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1028), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1038), .Y(n_1163) );
INVx4_ASAP7_75t_L g1164 ( .A(n_1157), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1050), .Y(n_1165) );
NAND2xp5_ASAP7_75t_L g1166 ( .A(n_1056), .B(n_1024), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1013), .Y(n_1167) );
AND2x4_ASAP7_75t_L g1168 ( .A(n_1157), .B(n_1095), .Y(n_1168) );
OA21x2_ASAP7_75t_L g1169 ( .A1(n_1123), .A2(n_1126), .B(n_1117), .Y(n_1169) );
NOR2xp67_ASAP7_75t_L g1170 ( .A(n_1113), .B(n_1090), .Y(n_1170) );
INVx2_ASAP7_75t_L g1171 ( .A(n_1128), .Y(n_1171) );
AO31x2_ASAP7_75t_L g1172 ( .A1(n_1096), .A2(n_1104), .A3(n_1109), .B(n_1103), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1046), .Y(n_1173) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1049), .Y(n_1174) );
INVx2_ASAP7_75t_L g1175 ( .A(n_1093), .Y(n_1175) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1154), .Y(n_1176) );
HB1xp67_ASAP7_75t_L g1177 ( .A(n_1076), .Y(n_1177) );
BUFx6f_ASAP7_75t_L g1178 ( .A(n_1016), .Y(n_1178) );
INVx1_ASAP7_75t_L g1179 ( .A(n_1063), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1180 ( .A(n_1159), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1159), .B(n_1035), .Y(n_1181) );
AND2x4_ASAP7_75t_L g1182 ( .A(n_1095), .B(n_1116), .Y(n_1182) );
NOR2xp33_ASAP7_75t_L g1183 ( .A(n_1031), .B(n_1088), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1071), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1185 ( .A(n_1130), .B(n_1018), .Y(n_1185) );
OR2x2_ASAP7_75t_L g1186 ( .A(n_1086), .B(n_1073), .Y(n_1186) );
BUFx2_ASAP7_75t_L g1187 ( .A(n_1124), .Y(n_1187) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_1124), .Y(n_1188) );
INVx2_ASAP7_75t_SL g1189 ( .A(n_1125), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g1190 ( .A(n_1016), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1019), .Y(n_1191) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1093), .Y(n_1192) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1110), .Y(n_1193) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1019), .Y(n_1194) );
BUFx2_ASAP7_75t_L g1195 ( .A(n_1127), .Y(n_1195) );
INVx2_ASAP7_75t_SL g1196 ( .A(n_1146), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_1089), .A2(n_1015), .B1(n_1021), .B2(n_1014), .Y(n_1197) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1016), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1136), .Y(n_1199) );
AOI22xp33_ASAP7_75t_SL g1200 ( .A1(n_1025), .A2(n_1039), .B1(n_1029), .B2(n_1021), .Y(n_1200) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1019), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1079), .B(n_1030), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1025), .B(n_1039), .Y(n_1203) );
INVxp67_ASAP7_75t_SL g1204 ( .A(n_1014), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1119), .Y(n_1205) );
INVxp67_ASAP7_75t_SL g1206 ( .A(n_1082), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1068), .B(n_1081), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1068), .B(n_1037), .Y(n_1208) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_1111), .Y(n_1209) );
BUFx6f_ASAP7_75t_L g1210 ( .A(n_1116), .Y(n_1210) );
INVx2_ASAP7_75t_L g1211 ( .A(n_1122), .Y(n_1211) );
AO31x2_ASAP7_75t_L g1212 ( .A1(n_1150), .A2(n_1131), .A3(n_1133), .B(n_1108), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1022), .B(n_1054), .Y(n_1213) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1051), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1022), .B(n_1040), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1216 ( .A(n_1097), .B(n_1098), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1032), .B(n_1033), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1032), .B(n_1033), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1120), .B(n_1045), .Y(n_1219) );
BUFx3_ASAP7_75t_L g1220 ( .A(n_1101), .Y(n_1220) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1114), .B(n_1034), .Y(n_1221) );
AND2x4_ASAP7_75t_L g1222 ( .A(n_1139), .B(n_1107), .Y(n_1222) );
AO31x2_ASAP7_75t_L g1223 ( .A1(n_1131), .A2(n_1108), .A3(n_1149), .B(n_1137), .Y(n_1223) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1045), .B(n_1023), .Y(n_1224) );
INVx2_ASAP7_75t_L g1225 ( .A(n_1041), .Y(n_1225) );
INVx3_ASAP7_75t_L g1226 ( .A(n_1115), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1043), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_1092), .Y(n_1228) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1017), .Y(n_1229) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1064), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1105), .B(n_1070), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1105), .B(n_1070), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1059), .B(n_1099), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1047), .B(n_1052), .Y(n_1234) );
OR2x2_ASAP7_75t_L g1235 ( .A(n_1100), .B(n_1094), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1036), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1026), .B(n_1048), .Y(n_1237) );
INVx2_ASAP7_75t_SL g1238 ( .A(n_1115), .Y(n_1238) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1053), .Y(n_1239) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1057), .Y(n_1240) );
AOI21xp33_ASAP7_75t_L g1241 ( .A1(n_1102), .A2(n_1100), .B(n_1145), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1010), .B(n_1044), .Y(n_1242) );
INVx2_ASAP7_75t_L g1243 ( .A(n_1057), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1115), .B(n_1065), .Y(n_1244) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_1009), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1147), .B(n_1072), .Y(n_1246) );
INVx4_ASAP7_75t_R g1247 ( .A(n_1060), .Y(n_1247) );
INVx2_ASAP7_75t_L g1248 ( .A(n_1115), .Y(n_1248) );
BUFx2_ASAP7_75t_L g1249 ( .A(n_1115), .Y(n_1249) );
AND2x4_ASAP7_75t_SL g1250 ( .A(n_1066), .B(n_1027), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1055), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1061), .B(n_1069), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1253 ( .A1(n_1106), .A2(n_1083), .B1(n_1058), .B2(n_1121), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_1138), .B(n_1148), .Y(n_1254) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1055), .Y(n_1255) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_1147), .Y(n_1256) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1055), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1118), .B(n_1135), .Y(n_1258) );
NAND2xp5_ASAP7_75t_L g1259 ( .A(n_1085), .B(n_1112), .Y(n_1259) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1129), .Y(n_1260) );
AND2x4_ASAP7_75t_L g1261 ( .A(n_1078), .B(n_1080), .Y(n_1261) );
AO31x2_ASAP7_75t_L g1262 ( .A1(n_1087), .A2(n_1091), .A3(n_1134), .B(n_1158), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1132), .B(n_1067), .Y(n_1263) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1144), .Y(n_1264) );
AND2x4_ASAP7_75t_L g1265 ( .A(n_1084), .B(n_1075), .Y(n_1265) );
INVx2_ASAP7_75t_L g1266 ( .A(n_1141), .Y(n_1266) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1123), .Y(n_1267) );
HB1xp67_ASAP7_75t_L g1268 ( .A(n_1042), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1142), .Y(n_1269) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_1143), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1151), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1140), .B(n_1153), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1273 ( .A(n_1074), .B(n_1077), .Y(n_1273) );
INVx2_ASAP7_75t_SL g1274 ( .A(n_1062), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1156), .B(n_1155), .Y(n_1275) );
INVxp67_ASAP7_75t_L g1276 ( .A(n_1011), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1177), .B(n_1152), .Y(n_1277) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1211), .Y(n_1278) );
INVx2_ASAP7_75t_SL g1279 ( .A(n_1209), .Y(n_1279) );
NAND4xp25_ASAP7_75t_L g1280 ( .A(n_1200), .B(n_1231), .C(n_1232), .D(n_1218), .Y(n_1280) );
BUFx3_ASAP7_75t_L g1281 ( .A(n_1196), .Y(n_1281) );
OAI22xp5_ASAP7_75t_SL g1282 ( .A1(n_1164), .A2(n_1183), .B1(n_1217), .B2(n_1196), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1205), .B(n_1195), .Y(n_1283) );
INVx3_ASAP7_75t_L g1284 ( .A(n_1226), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1165), .B(n_1181), .Y(n_1285) );
BUFx3_ASAP7_75t_L g1286 ( .A(n_1210), .Y(n_1286) );
INVx2_ASAP7_75t_L g1287 ( .A(n_1211), .Y(n_1287) );
HB1xp67_ASAP7_75t_L g1288 ( .A(n_1195), .Y(n_1288) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1173), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1202), .B(n_1207), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1291 ( .A(n_1181), .B(n_1184), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1174), .Y(n_1292) );
INVx3_ASAP7_75t_L g1293 ( .A(n_1226), .Y(n_1293) );
NAND4xp25_ASAP7_75t_L g1294 ( .A(n_1231), .B(n_1232), .C(n_1235), .D(n_1203), .Y(n_1294) );
OAI221xp5_ASAP7_75t_L g1295 ( .A1(n_1216), .A2(n_1236), .B1(n_1268), .B2(n_1221), .C(n_1237), .Y(n_1295) );
HB1xp67_ASAP7_75t_L g1296 ( .A(n_1199), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1207), .B(n_1203), .Y(n_1297) );
INVx1_ASAP7_75t_SL g1298 ( .A(n_1220), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1205), .B(n_1180), .Y(n_1299) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1176), .Y(n_1300) );
OAI22xp5_ASAP7_75t_L g1301 ( .A1(n_1208), .A2(n_1213), .B1(n_1274), .B2(n_1215), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1186), .B(n_1161), .Y(n_1302) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1179), .Y(n_1303) );
BUFx2_ASAP7_75t_L g1304 ( .A(n_1188), .Y(n_1304) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1166), .Y(n_1305) );
NOR2x1_ASAP7_75t_L g1306 ( .A(n_1164), .B(n_1170), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1162), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1308 ( .A1(n_1227), .A2(n_1214), .B1(n_1215), .B2(n_1241), .C(n_1239), .Y(n_1308) );
NOR2xp33_ASAP7_75t_L g1309 ( .A(n_1208), .B(n_1235), .Y(n_1309) );
NAND2x1p5_ASAP7_75t_L g1310 ( .A(n_1164), .B(n_1220), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1311 ( .A(n_1245), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1199), .Y(n_1312) );
OAI31xp33_ASAP7_75t_L g1313 ( .A1(n_1197), .A2(n_1224), .A3(n_1250), .B(n_1274), .Y(n_1313) );
BUFx2_ASAP7_75t_L g1314 ( .A(n_1187), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1315 ( .A1(n_1224), .A2(n_1242), .B1(n_1228), .B2(n_1250), .Y(n_1315) );
NOR2xp33_ASAP7_75t_L g1316 ( .A(n_1233), .B(n_1168), .Y(n_1316) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1163), .B(n_1206), .Y(n_1317) );
OR2x6_ASAP7_75t_L g1318 ( .A(n_1187), .B(n_1249), .Y(n_1318) );
AOI22xp5_ASAP7_75t_L g1319 ( .A1(n_1234), .A2(n_1168), .B1(n_1252), .B2(n_1253), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1320 ( .A(n_1163), .B(n_1189), .Y(n_1320) );
AOI22xp5_ASAP7_75t_L g1321 ( .A1(n_1168), .A2(n_1252), .B1(n_1219), .B2(n_1204), .Y(n_1321) );
INVx4_ASAP7_75t_L g1322 ( .A(n_1210), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1271), .B(n_1160), .Y(n_1323) );
OR2x2_ASAP7_75t_L g1324 ( .A(n_1185), .B(n_1160), .Y(n_1324) );
HB1xp67_ASAP7_75t_L g1325 ( .A(n_1193), .Y(n_1325) );
AND2x2_ASAP7_75t_L g1326 ( .A(n_1258), .B(n_1275), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1210), .B(n_1182), .Y(n_1327) );
OR2x6_ASAP7_75t_L g1328 ( .A(n_1249), .B(n_1256), .Y(n_1328) );
NAND4xp75_ASAP7_75t_L g1329 ( .A(n_1275), .B(n_1244), .C(n_1247), .D(n_1269), .Y(n_1329) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1172), .Y(n_1330) );
INVx2_ASAP7_75t_SL g1331 ( .A(n_1238), .Y(n_1331) );
AND2x4_ASAP7_75t_L g1332 ( .A(n_1222), .B(n_1226), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1333 ( .A(n_1182), .B(n_1238), .Y(n_1333) );
AOI22xp5_ASAP7_75t_L g1334 ( .A1(n_1182), .A2(n_1244), .B1(n_1229), .B2(n_1259), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1222), .B(n_1258), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1336 ( .A(n_1222), .B(n_1272), .Y(n_1336) );
INVx2_ASAP7_75t_L g1337 ( .A(n_1175), .Y(n_1337) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1172), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1172), .Y(n_1339) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1192), .Y(n_1340) );
NAND2xp5_ASAP7_75t_SL g1341 ( .A(n_1248), .B(n_1270), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1272), .B(n_1194), .Y(n_1342) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1191), .B(n_1201), .Y(n_1343) );
INVx3_ASAP7_75t_L g1344 ( .A(n_1178), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1191), .B(n_1201), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1194), .B(n_1260), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1269), .B(n_1260), .Y(n_1347) );
OR2x2_ASAP7_75t_SL g1348 ( .A(n_1251), .B(n_1263), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1256), .B(n_1198), .Y(n_1349) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_1246), .A2(n_1270), .B1(n_1255), .B2(n_1265), .Y(n_1350) );
NAND2xp5_ASAP7_75t_SL g1351 ( .A(n_1255), .B(n_1257), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1246), .B(n_1193), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1326), .B(n_1212), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1326), .B(n_1267), .Y(n_1354) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1343), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1356 ( .A(n_1305), .B(n_1276), .Y(n_1356) );
NAND3xp33_ASAP7_75t_L g1357 ( .A(n_1308), .B(n_1255), .C(n_1251), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1342), .B(n_1335), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1309), .B(n_1171), .Y(n_1359) );
NAND4xp25_ASAP7_75t_L g1360 ( .A(n_1280), .B(n_1265), .C(n_1254), .D(n_1273), .Y(n_1360) );
INVx2_ASAP7_75t_L g1361 ( .A(n_1278), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1362 ( .A(n_1332), .B(n_1212), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1345), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1342), .B(n_1212), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1297), .B(n_1212), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1336), .B(n_1171), .Y(n_1366) );
INVx1_ASAP7_75t_SL g1367 ( .A(n_1281), .Y(n_1367) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1307), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1330), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1309), .B(n_1266), .Y(n_1370) );
AND2x4_ASAP7_75t_L g1371 ( .A(n_1332), .B(n_1192), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1302), .B(n_1223), .Y(n_1372) );
OR2x6_ASAP7_75t_L g1373 ( .A(n_1328), .B(n_1240), .Y(n_1373) );
AND2x4_ASAP7_75t_L g1374 ( .A(n_1332), .B(n_1223), .Y(n_1374) );
INVx2_ASAP7_75t_L g1375 ( .A(n_1287), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1285), .B(n_1288), .Y(n_1376) );
NOR2x1p5_ASAP7_75t_SL g1377 ( .A(n_1329), .B(n_1240), .Y(n_1377) );
AOI22xp33_ASAP7_75t_L g1378 ( .A1(n_1294), .A2(n_1265), .B1(n_1261), .B2(n_1264), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1323), .B(n_1223), .Y(n_1379) );
INVx1_ASAP7_75t_SL g1380 ( .A(n_1281), .Y(n_1380) );
AND2x4_ASAP7_75t_L g1381 ( .A(n_1328), .B(n_1262), .Y(n_1381) );
BUFx2_ASAP7_75t_L g1382 ( .A(n_1318), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1290), .B(n_1264), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1338), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1346), .B(n_1262), .Y(n_1385) );
AND2x2_ASAP7_75t_SL g1386 ( .A(n_1288), .B(n_1243), .Y(n_1386) );
INVx1_ASAP7_75t_SL g1387 ( .A(n_1298), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1311), .B(n_1178), .Y(n_1388) );
CKINVDCx16_ASAP7_75t_R g1389 ( .A(n_1282), .Y(n_1389) );
AND2x4_ASAP7_75t_L g1390 ( .A(n_1328), .B(n_1262), .Y(n_1390) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_1311), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1299), .B(n_1262), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1299), .B(n_1262), .Y(n_1393) );
AND2x4_ASAP7_75t_SL g1394 ( .A(n_1279), .B(n_1190), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1395 ( .A(n_1296), .B(n_1169), .Y(n_1395) );
OR2x2_ASAP7_75t_L g1396 ( .A(n_1352), .B(n_1291), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1296), .B(n_1169), .Y(n_1397) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1312), .B(n_1169), .Y(n_1398) );
OAI33xp33_ASAP7_75t_L g1399 ( .A1(n_1301), .A2(n_1243), .A3(n_1225), .B1(n_1230), .B2(n_1167), .B3(n_1261), .Y(n_1399) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_1328), .B(n_1225), .Y(n_1400) );
OAI211xp5_ASAP7_75t_SL g1401 ( .A1(n_1295), .A2(n_1230), .B(n_1261), .C(n_1190), .Y(n_1401) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1289), .B(n_1190), .Y(n_1402) );
INVx1_ASAP7_75t_SL g1403 ( .A(n_1304), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1404 ( .A(n_1325), .B(n_1190), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1339), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1406 ( .A(n_1354), .B(n_1277), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1358), .B(n_1349), .Y(n_1407) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1369), .Y(n_1408) );
AND2x4_ASAP7_75t_L g1409 ( .A(n_1374), .B(n_1318), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1358), .B(n_1392), .Y(n_1410) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1361), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1369), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1384), .Y(n_1413) );
INVx2_ASAP7_75t_SL g1414 ( .A(n_1394), .Y(n_1414) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1376), .Y(n_1415) );
OAI21xp5_ASAP7_75t_L g1416 ( .A1(n_1401), .A2(n_1313), .B(n_1347), .Y(n_1416) );
OR2x2_ASAP7_75t_L g1417 ( .A(n_1354), .B(n_1283), .Y(n_1417) );
INVx1_ASAP7_75t_SL g1418 ( .A(n_1391), .Y(n_1418) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1384), .Y(n_1419) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1405), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1405), .Y(n_1421) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1387), .B(n_1319), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1393), .B(n_1283), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1393), .B(n_1321), .Y(n_1424) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1368), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1353), .B(n_1350), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1427 ( .A(n_1364), .B(n_1337), .Y(n_1427) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1396), .B(n_1303), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1429 ( .A(n_1383), .B(n_1300), .Y(n_1429) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1368), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1372), .B(n_1324), .Y(n_1431) );
AND2x4_ASAP7_75t_L g1432 ( .A(n_1374), .B(n_1318), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1355), .B(n_1292), .Y(n_1433) );
AOI221x1_ASAP7_75t_L g1434 ( .A1(n_1360), .A2(n_1317), .B1(n_1284), .B2(n_1293), .C(n_1344), .Y(n_1434) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1363), .Y(n_1435) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_1360), .A2(n_1315), .B1(n_1316), .B2(n_1334), .Y(n_1436) );
AOI221x1_ASAP7_75t_L g1437 ( .A1(n_1357), .A2(n_1284), .B1(n_1293), .B2(n_1344), .C(n_1320), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1364), .B(n_1365), .Y(n_1438) );
NOR2xp67_ASAP7_75t_L g1439 ( .A(n_1357), .B(n_1331), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1365), .B(n_1340), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1363), .B(n_1315), .Y(n_1441) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1375), .Y(n_1442) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1356), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_1436), .A2(n_1378), .B1(n_1362), .B2(n_1316), .Y(n_1444) );
INVx1_ASAP7_75t_SL g1445 ( .A(n_1418), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1425), .Y(n_1446) );
INVxp33_ASAP7_75t_L g1447 ( .A(n_1439), .Y(n_1447) );
OAI31xp33_ASAP7_75t_L g1448 ( .A1(n_1422), .A2(n_1380), .A3(n_1367), .B(n_1403), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1449 ( .A1(n_1443), .A2(n_1399), .B1(n_1389), .B2(n_1370), .C(n_1359), .Y(n_1449) );
NOR2xp67_ASAP7_75t_L g1450 ( .A(n_1410), .B(n_1381), .Y(n_1450) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1435), .Y(n_1451) );
INVx2_ASAP7_75t_SL g1452 ( .A(n_1414), .Y(n_1452) );
NAND3xp33_ASAP7_75t_L g1453 ( .A(n_1434), .B(n_1390), .C(n_1381), .Y(n_1453) );
NAND2xp33_ASAP7_75t_L g1454 ( .A(n_1414), .B(n_1306), .Y(n_1454) );
A2O1A1Ixp33_ASAP7_75t_L g1455 ( .A1(n_1416), .A2(n_1377), .B(n_1382), .C(n_1388), .Y(n_1455) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_1441), .A2(n_1348), .B1(n_1310), .B2(n_1382), .Y(n_1456) );
AOI22xp33_ASAP7_75t_SL g1457 ( .A1(n_1409), .A2(n_1314), .B1(n_1381), .B2(n_1390), .Y(n_1457) );
OAI22xp5_ASAP7_75t_L g1458 ( .A1(n_1417), .A2(n_1310), .B1(n_1318), .B2(n_1373), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1435), .Y(n_1459) );
INVx2_ASAP7_75t_L g1460 ( .A(n_1411), .Y(n_1460) );
INVx2_ASAP7_75t_L g1461 ( .A(n_1411), .Y(n_1461) );
OAI21xp5_ASAP7_75t_L g1462 ( .A1(n_1437), .A2(n_1331), .B(n_1386), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1463 ( .A1(n_1431), .A2(n_1373), .B1(n_1333), .B2(n_1386), .Y(n_1463) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1438), .B(n_1379), .Y(n_1464) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1425), .Y(n_1465) );
INVx1_ASAP7_75t_L g1466 ( .A(n_1408), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1438), .B(n_1379), .Y(n_1467) );
NAND2xp5_ASAP7_75t_L g1468 ( .A(n_1415), .B(n_1385), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1469 ( .A(n_1450), .B(n_1407), .Y(n_1469) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1446), .Y(n_1470) );
OAI21xp5_ASAP7_75t_L g1471 ( .A1(n_1455), .A2(n_1437), .B(n_1428), .Y(n_1471) );
AOI22xp33_ASAP7_75t_L g1472 ( .A1(n_1444), .A2(n_1426), .B1(n_1424), .B2(n_1362), .Y(n_1472) );
INVx2_ASAP7_75t_SL g1473 ( .A(n_1452), .Y(n_1473) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1449), .B(n_1423), .Y(n_1474) );
NAND3xp33_ASAP7_75t_L g1475 ( .A(n_1448), .B(n_1433), .C(n_1429), .Y(n_1475) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1446), .Y(n_1476) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1466), .Y(n_1477) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1445), .B(n_1406), .Y(n_1478) );
INVx2_ASAP7_75t_L g1479 ( .A(n_1460), .Y(n_1479) );
XNOR2xp5_ASAP7_75t_L g1480 ( .A(n_1457), .B(n_1407), .Y(n_1480) );
AND2x2_ASAP7_75t_L g1481 ( .A(n_1464), .B(n_1440), .Y(n_1481) );
OAI21xp5_ASAP7_75t_L g1482 ( .A1(n_1455), .A2(n_1386), .B(n_1381), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1483 ( .A(n_1467), .B(n_1440), .Y(n_1483) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1466), .Y(n_1484) );
NAND2xp5_ASAP7_75t_L g1485 ( .A(n_1468), .B(n_1427), .Y(n_1485) );
AOI31xp33_ASAP7_75t_L g1486 ( .A1(n_1447), .A2(n_1432), .A3(n_1409), .B(n_1431), .Y(n_1486) );
INVx2_ASAP7_75t_SL g1487 ( .A(n_1452), .Y(n_1487) );
OAI21xp33_ASAP7_75t_L g1488 ( .A1(n_1474), .A2(n_1447), .B(n_1453), .Y(n_1488) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1469), .B(n_1427), .Y(n_1489) );
AOI22xp5_ASAP7_75t_L g1490 ( .A1(n_1472), .A2(n_1456), .B1(n_1463), .B2(n_1458), .Y(n_1490) );
AOI21xp33_ASAP7_75t_L g1491 ( .A1(n_1471), .A2(n_1454), .B(n_1462), .Y(n_1491) );
INVx2_ASAP7_75t_SL g1492 ( .A(n_1473), .Y(n_1492) );
AOI22xp5_ASAP7_75t_L g1493 ( .A1(n_1480), .A2(n_1362), .B1(n_1454), .B2(n_1390), .Y(n_1493) );
NOR2x1_ASAP7_75t_L g1494 ( .A(n_1486), .B(n_1284), .Y(n_1494) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_1486), .A2(n_1373), .B1(n_1390), .B2(n_1459), .Y(n_1495) );
AOI21xp5_ASAP7_75t_L g1496 ( .A1(n_1480), .A2(n_1451), .B(n_1465), .Y(n_1496) );
O2A1O1Ixp33_ASAP7_75t_L g1497 ( .A1(n_1475), .A2(n_1341), .B(n_1430), .C(n_1461), .Y(n_1497) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_1488), .A2(n_1475), .B1(n_1478), .B2(n_1482), .C(n_1473), .Y(n_1498) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_1491), .A2(n_1487), .B1(n_1476), .B2(n_1484), .C(n_1470), .Y(n_1499) );
AOI21xp5_ASAP7_75t_L g1500 ( .A1(n_1496), .A2(n_1479), .B(n_1484), .Y(n_1500) );
A2O1A1Ixp33_ASAP7_75t_L g1501 ( .A1(n_1494), .A2(n_1377), .B(n_1483), .C(n_1481), .Y(n_1501) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1492), .Y(n_1502) );
AOI221xp5_ASAP7_75t_L g1503 ( .A1(n_1497), .A2(n_1477), .B1(n_1485), .B2(n_1483), .C(n_1479), .Y(n_1503) );
AOI321xp33_ASAP7_75t_L g1504 ( .A1(n_1495), .A2(n_1374), .A3(n_1341), .B1(n_1408), .B2(n_1412), .C(n_1421), .Y(n_1504) );
NOR4xp75_ASAP7_75t_SL g1505 ( .A(n_1498), .B(n_1493), .C(n_1490), .D(n_1402), .Y(n_1505) );
NAND3xp33_ASAP7_75t_L g1506 ( .A(n_1499), .B(n_1419), .C(n_1412), .Y(n_1506) );
AOI22xp5_ASAP7_75t_L g1507 ( .A1(n_1502), .A2(n_1489), .B1(n_1374), .B2(n_1373), .Y(n_1507) );
AOI221xp5_ASAP7_75t_L g1508 ( .A1(n_1503), .A2(n_1419), .B1(n_1413), .B2(n_1421), .C(n_1420), .Y(n_1508) );
BUFx6f_ASAP7_75t_L g1509 ( .A(n_1501), .Y(n_1509) );
OAI221xp5_ASAP7_75t_SL g1510 ( .A1(n_1505), .A2(n_1504), .B1(n_1500), .B2(n_1373), .C(n_1327), .Y(n_1510) );
INVxp33_ASAP7_75t_L g1511 ( .A(n_1509), .Y(n_1511) );
OAI22xp33_ASAP7_75t_L g1512 ( .A1(n_1511), .A2(n_1507), .B1(n_1506), .B2(n_1508), .Y(n_1512) );
INVx4_ASAP7_75t_L g1513 ( .A(n_1512), .Y(n_1513) );
AOI221xp5_ASAP7_75t_L g1514 ( .A1(n_1513), .A2(n_1510), .B1(n_1442), .B2(n_1351), .C(n_1293), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_1514), .A2(n_1322), .B1(n_1286), .B2(n_1400), .Y(n_1515) );
AOI322xp5_ASAP7_75t_L g1516 ( .A1(n_1515), .A2(n_1400), .A3(n_1366), .B1(n_1404), .B2(n_1371), .C1(n_1397), .C2(n_1395), .Y(n_1516) );
AOI21xp5_ASAP7_75t_L g1517 ( .A1(n_1516), .A2(n_1397), .B(n_1398), .Y(n_1517) );
endmodule