module fake_jpeg_15126_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx3_ASAP7_75t_SL g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx5_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

OR2x2_ASAP7_75t_SL g14 ( 
.A(n_7),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_18),
.B1(n_12),
.B2(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_9),
.B(n_5),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_2),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_6),
.C(n_3),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_16),
.A2(n_12),
.B1(n_11),
.B2(n_10),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_22),
.A2(n_23),
.B(n_2),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_14),
.A3(n_19),
.B1(n_18),
.B2(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_21),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.C(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_31),
.B(n_24),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_32),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_5),
.B(n_6),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_3),
.C(n_4),
.Y(n_36)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_4),
.C(n_17),
.Y(n_37)
);


endmodule