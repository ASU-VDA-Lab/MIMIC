module fake_jpeg_11560_n_447 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_9),
.B(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_60),
.B(n_66),
.Y(n_126)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_62),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_70),
.Y(n_164)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_72),
.B(n_73),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_30),
.B(n_15),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_74),
.B(n_83),
.Y(n_143)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_75),
.B(n_82),
.Y(n_134)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

CKINVDCx6p67_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_77),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_78),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_20),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_30),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_35),
.B(n_0),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_84),
.B(n_93),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_42),
.B(n_1),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_87),
.Y(n_155)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_25),
.Y(n_86)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_1),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_89),
.Y(n_179)
);

INVx2_ASAP7_75t_R g90 ( 
.A(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_90),
.B(n_105),
.Y(n_138)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_26),
.Y(n_91)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_92),
.B(n_100),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_14),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_26),
.Y(n_95)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_96),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_99),
.B(n_103),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_28),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_101),
.B(n_102),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_2),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_43),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_104),
.B(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_38),
.B(n_14),
.Y(n_105)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_26),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_38),
.B(n_3),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_108),
.B(n_109),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_113),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g111 ( 
.A(n_26),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_115),
.B1(n_117),
.B2(n_56),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_28),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_114),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

BUFx24_ASAP7_75t_L g115 ( 
.A(n_26),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_118),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_48),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_41),
.B(n_5),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_119),
.B(n_12),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_49),
.B1(n_32),
.B2(n_41),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_120),
.A2(n_137),
.B1(n_157),
.B2(n_163),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_59),
.A2(n_53),
.B1(n_21),
.B2(n_47),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_121),
.A2(n_142),
.B1(n_149),
.B2(n_154),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_122),
.Y(n_245)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_34),
.B(n_37),
.C(n_40),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_130),
.A2(n_181),
.B(n_185),
.C(n_163),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_49),
.B1(n_32),
.B2(n_45),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_115),
.A2(n_29),
.B1(n_49),
.B2(n_32),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_140),
.A2(n_141),
.B1(n_146),
.B2(n_156),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_29),
.B1(n_49),
.B2(n_53),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_63),
.A2(n_53),
.B1(n_44),
.B2(n_45),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_95),
.A2(n_56),
.B1(n_19),
.B2(n_21),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_64),
.A2(n_56),
.B1(n_44),
.B2(n_43),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_80),
.B(n_61),
.C(n_76),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_153),
.B(n_178),
.C(n_181),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_67),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_106),
.A2(n_56),
.B1(n_34),
.B2(n_33),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_70),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_94),
.A2(n_56),
.B1(n_40),
.B2(n_51),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_158),
.A2(n_165),
.B1(n_166),
.B2(n_174),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_78),
.A2(n_19),
.B1(n_51),
.B2(n_47),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_89),
.A2(n_37),
.B1(n_33),
.B2(n_57),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_88),
.A2(n_57),
.B1(n_31),
.B2(n_58),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_79),
.A2(n_57),
.B1(n_31),
.B2(n_7),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_170),
.A2(n_175),
.B1(n_182),
.B2(n_184),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_107),
.A2(n_31),
.B1(n_68),
.B2(n_62),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_81),
.A2(n_58),
.B1(n_28),
.B2(n_8),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_91),
.B(n_58),
.C(n_6),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_62),
.A2(n_58),
.B1(n_6),
.B2(n_8),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_180),
.A2(n_183),
.B1(n_189),
.B2(n_191),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_97),
.A2(n_58),
.B1(n_8),
.B2(n_9),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_99),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_114),
.A2(n_117),
.B1(n_113),
.B2(n_109),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_103),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_187),
.B(n_138),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_114),
.A2(n_12),
.B1(n_13),
.B2(n_117),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_77),
.A2(n_69),
.B1(n_111),
.B2(n_118),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_176),
.Y(n_192)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_192),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g193 ( 
.A(n_143),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_193),
.B(n_201),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_194),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_136),
.B(n_77),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_196),
.Y(n_286)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_130),
.A2(n_111),
.B(n_188),
.C(n_144),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_197),
.A2(n_230),
.B(n_195),
.C(n_198),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_136),
.B(n_186),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_206),
.Y(n_265)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_190),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_200),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_133),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_126),
.Y(n_202)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_202),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_203),
.B(n_205),
.Y(n_296)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_148),
.A2(n_187),
.A3(n_188),
.B1(n_123),
.B2(n_136),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_204),
.B(n_249),
.Y(n_275)
);

OR2x4_ASAP7_75t_L g205 ( 
.A(n_138),
.B(n_168),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_148),
.B(n_123),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_149),
.A2(n_154),
.B1(n_142),
.B2(n_129),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_208),
.A2(n_237),
.B1(n_241),
.B2(n_199),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_171),
.B(n_167),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_209),
.B(n_216),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_210),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_177),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_251),
.C(n_195),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g300 ( 
.A(n_213),
.Y(n_300)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_151),
.Y(n_214)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_155),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_215),
.B(n_219),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_178),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_162),
.Y(n_217)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_173),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_218),
.B(n_227),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_169),
.B(n_147),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_145),
.B(n_173),
.Y(n_221)
);

NAND3xp33_ASAP7_75t_L g258 ( 
.A(n_221),
.B(n_226),
.C(n_235),
.Y(n_258)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

INVx13_ASAP7_75t_L g260 ( 
.A(n_223),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_124),
.Y(n_224)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_224),
.Y(n_277)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_177),
.B(n_150),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_184),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_150),
.B(n_159),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_228),
.B(n_231),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_159),
.B(n_128),
.Y(n_231)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_125),
.Y(n_232)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_132),
.A2(n_161),
.B1(n_152),
.B2(n_172),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_233),
.A2(n_229),
.B1(n_252),
.B2(n_212),
.Y(n_274)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_175),
.A2(n_185),
.B1(n_127),
.B2(n_161),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_234),
.B(n_246),
.Y(n_288)
);

OR2x2_ASAP7_75t_SL g235 ( 
.A(n_147),
.B(n_131),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_242),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_129),
.A2(n_132),
.B1(n_139),
.B2(n_152),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_131),
.B(n_179),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_238),
.B(n_254),
.Y(n_279)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_240),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_125),
.A2(n_139),
.B1(n_152),
.B2(n_164),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_125),
.A2(n_139),
.B1(n_164),
.B2(n_172),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_243),
.A2(n_194),
.B1(n_224),
.B2(n_210),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_164),
.B(n_172),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_160),
.B(n_135),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_247),
.B(n_211),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_248),
.Y(n_287)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_176),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_253),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_136),
.B(n_148),
.C(n_153),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_124),
.Y(n_252)
);

INVx11_ASAP7_75t_L g295 ( 
.A(n_252),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_144),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_155),
.B(n_168),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_255),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_211),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_257),
.B(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_259),
.B(n_299),
.C(n_275),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_270),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_251),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g306 ( 
.A(n_269),
.B(n_197),
.CI(n_222),
.CON(n_306),
.SN(n_306)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_274),
.A2(n_284),
.B1(n_302),
.B2(n_263),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_275),
.B(n_229),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_209),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_227),
.A2(n_199),
.B1(n_206),
.B2(n_216),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_289),
.B(n_305),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_249),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_291),
.B(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_214),
.B(n_230),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_192),
.B(n_196),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_247),
.C(n_245),
.Y(n_299)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

BUFx24_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_235),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_263),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_212),
.B(n_217),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_306),
.B(n_319),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_307),
.B(n_337),
.Y(n_350)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_239),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_308),
.Y(n_365)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_310),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_207),
.B(n_234),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_311),
.A2(n_320),
.B(n_333),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_278),
.B(n_220),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_248),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_271),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_234),
.B(n_240),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_266),
.A2(n_200),
.B(n_225),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_340),
.Y(n_356)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_256),
.Y(n_323)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_267),
.B(n_255),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_324),
.B(n_331),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_280),
.A2(n_232),
.B1(n_233),
.B2(n_288),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_327),
.A2(n_329),
.B1(n_332),
.B2(n_282),
.Y(n_353)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_286),
.Y(n_328)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_291),
.A2(n_284),
.B1(n_267),
.B2(n_265),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_268),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_282),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_296),
.B(n_261),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_265),
.A2(n_304),
.B1(n_259),
.B2(n_289),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_299),
.A2(n_300),
.B(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_334),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_335),
.A2(n_298),
.B1(n_285),
.B2(n_262),
.Y(n_346)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_339),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_257),
.A2(n_269),
.B(n_258),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_338),
.A2(n_307),
.B(n_325),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_268),
.B(n_301),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_294),
.C(n_273),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_296),
.B(n_294),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_341),
.B(n_342),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_300),
.B(n_298),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_346),
.B(n_354),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_295),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_347),
.B(n_333),
.C(n_321),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_308),
.A2(n_277),
.B1(n_262),
.B2(n_264),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_361),
.Y(n_371)
);

AOI32xp33_ASAP7_75t_L g351 ( 
.A1(n_313),
.A2(n_295),
.A3(n_287),
.B1(n_285),
.B2(n_260),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_363),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_353),
.B(n_311),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_327),
.A2(n_277),
.B1(n_264),
.B2(n_290),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_357),
.A2(n_358),
.B1(n_342),
.B2(n_336),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_290),
.B1(n_281),
.B2(n_287),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_308),
.A2(n_281),
.B1(n_287),
.B2(n_260),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_287),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_362),
.B(n_368),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_312),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_320),
.A2(n_303),
.B1(n_313),
.B2(n_324),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_331),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_369),
.B(n_318),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_332),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_373),
.B(n_377),
.C(n_381),
.Y(n_397)
);

OAI21xp33_ASAP7_75t_L g374 ( 
.A1(n_366),
.A2(n_337),
.B(n_333),
.Y(n_374)
);

NOR3xp33_ASAP7_75t_SL g394 ( 
.A(n_374),
.B(n_360),
.C(n_365),
.Y(n_394)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_359),
.Y(n_375)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_375),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_376),
.B(n_387),
.Y(n_400)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_338),
.C(n_340),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_356),
.B(n_309),
.C(n_330),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_350),
.B(n_309),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_350),
.B(n_326),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_317),
.Y(n_385)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_385),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_317),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_355),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_326),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_363),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_389),
.Y(n_395)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_343),
.Y(n_390)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_390),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_391),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g398 ( 
.A1(n_392),
.A2(n_393),
.B1(n_365),
.B2(n_380),
.Y(n_398)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_380),
.A2(n_349),
.B1(n_348),
.B2(n_361),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_373),
.B(n_381),
.C(n_382),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_408),
.C(n_386),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_355),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_380),
.A2(n_349),
.B1(n_346),
.B2(n_344),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_377),
.B(n_353),
.C(n_344),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_362),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_410),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_367),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_378),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_412),
.B(n_414),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_383),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_395),
.Y(n_415)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_384),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_416),
.B(n_339),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_371),
.B1(n_351),
.B2(n_357),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_407),
.B1(n_410),
.B2(n_409),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_388),
.B(n_352),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_L g425 ( 
.A1(n_418),
.A2(n_422),
.B(n_394),
.C(n_402),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_393),
.B1(n_306),
.B2(n_367),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_400),
.B(n_315),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_408),
.A2(n_358),
.B(n_314),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_424),
.B(n_426),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_425),
.B(n_429),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_402),
.C(n_407),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_427),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_405),
.C(n_396),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_416),
.C(n_422),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_430),
.B(n_431),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_423),
.B(n_418),
.C(n_420),
.Y(n_431)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_432),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_421),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_419),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_437),
.B(n_434),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_428),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_440),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_436),
.B(n_433),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_443),
.A2(n_413),
.B(n_403),
.Y(n_444)
);

AOI321xp33_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_442),
.A3(n_399),
.B1(n_364),
.B2(n_345),
.C(n_310),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_445),
.B(n_364),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_316),
.Y(n_447)
);


endmodule