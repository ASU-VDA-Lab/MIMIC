module fake_jpeg_4453_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_20;
wire n_59;
wire n_35;
wire n_71;
wire n_68;
wire n_52;
wire n_48;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_44;
wire n_24;
wire n_28;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx10_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_41),
.Y(n_57)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_24),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_47),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_3),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_4),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_5),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_30),
.A2(n_15),
.B1(n_16),
.B2(n_33),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_36),
.B1(n_37),
.B2(n_22),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_53),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.C(n_59),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_57),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.B(n_49),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_58),
.B(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_55),
.Y(n_66)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_51),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_67),
.B(n_42),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_70),
.B(n_55),
.C(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_23),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_50),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_47),
.A3(n_60),
.B1(n_34),
.B2(n_52),
.C1(n_48),
.C2(n_54),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_43),
.Y(n_74)
);


endmodule