module fake_netlist_6_2290_n_1069 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_229, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1069);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1069;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_278;
wire n_362;
wire n_341;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_988;
wire n_969;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_1057;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_638;
wire n_910;
wire n_486;
wire n_947;
wire n_381;
wire n_911;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_904;
wire n_366;
wire n_870;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_1041;
wire n_252;
wire n_757;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_982;
wire n_964;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_1055;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1063;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_137),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_88),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_188),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_138),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_136),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_53),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_176),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_224),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_23),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_233),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_189),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_106),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_2),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_76),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_223),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_44),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_125),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_56),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_74),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_69),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_134),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_169),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_131),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_107),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_37),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_160),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_112),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_185),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_61),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_144),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_151),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_117),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_8),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_232),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_119),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_41),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_55),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_21),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_236),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g283 ( 
.A(n_179),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_7),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_190),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_164),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_184),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_124),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_229),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_128),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_219),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_110),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_228),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_181),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_198),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_122),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_73),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_142),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_0),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_227),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_58),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_154),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_135),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_120),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_6),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_20),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_70),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_17),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_140),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_220),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_167),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_159),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_153),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_78),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_222),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_130),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_40),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_211),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_52),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_57),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_15),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_79),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_40),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_95),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_182),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_96),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_48),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_59),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_21),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_82),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_168),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_93),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_150),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_19),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_207),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_158),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_253),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_332),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_271),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_322),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_244),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_325),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_293),
.B(n_0),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_273),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_247),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_256),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_256),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_283),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_305),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_307),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_309),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_1),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_292),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_324),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_254),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_276),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_283),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_330),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_242),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_279),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_238),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_325),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_242),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_281),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_241),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_312),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_243),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_334),
.B(n_1),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_287),
.B(n_2),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_245),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_246),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_287),
.B(n_3),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_239),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_240),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_255),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_248),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_259),
.Y(n_384)
);

INVxp67_ASAP7_75t_SL g385 ( 
.A(n_260),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_249),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_266),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_269),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_250),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_313),
.B(n_3),
.Y(n_390)
);

INVxp33_ASAP7_75t_L g391 ( 
.A(n_247),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_252),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_257),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_272),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_346),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_351),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_369),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_343),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_387),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_343),
.Y(n_402)
);

OAI21x1_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_277),
.B(n_274),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_339),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_299),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_R g406 ( 
.A(n_365),
.B(n_261),
.Y(n_406)
);

NAND2xp33_ASAP7_75t_SL g407 ( 
.A(n_353),
.B(n_299),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_377),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_344),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_372),
.B(n_345),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_368),
.B(n_282),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_363),
.B(n_348),
.Y(n_412)
);

OR2x6_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_285),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_349),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_286),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_383),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_358),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_348),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

OR2x6_ASAP7_75t_L g421 ( 
.A(n_369),
.B(n_290),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_382),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_384),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_389),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_355),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_367),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_394),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

OA21x2_ASAP7_75t_L g431 ( 
.A1(n_393),
.A2(n_294),
.B(n_291),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_361),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_371),
.B(n_298),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_371),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_340),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_362),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_373),
.B(n_306),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_341),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_356),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_356),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_350),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_370),
.Y(n_445)
);

OA21x2_ASAP7_75t_L g446 ( 
.A1(n_374),
.A2(n_317),
.B(n_308),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_378),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_360),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_359),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_375),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_347),
.A2(n_321),
.B(n_319),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_364),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_373),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_366),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_342),
.A2(n_318),
.B1(n_284),
.B2(n_251),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_450),
.B(n_379),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_432),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_450),
.B(n_390),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_292),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_450),
.B(n_400),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_399),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_398),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_416),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_396),
.A2(n_386),
.B1(n_376),
.B2(n_392),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_450),
.B(n_268),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_400),
.B(n_292),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_455),
.B(n_318),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_420),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_376),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_401),
.Y(n_475)
);

INVx8_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_418),
.B(n_292),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_364),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_422),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_442),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_398),
.B(n_323),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_418),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_433),
.B(n_386),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_408),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_423),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_399),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_392),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g491 ( 
.A(n_425),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_439),
.B(n_312),
.Y(n_492)
);

INVxp67_ASAP7_75t_SL g493 ( 
.A(n_418),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_404),
.Y(n_494)
);

AND2x6_ASAP7_75t_L g495 ( 
.A(n_411),
.B(n_268),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

INVxp33_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_408),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_399),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_414),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_427),
.B(n_391),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_445),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_445),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_402),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_447),
.Y(n_505)
);

OAI21xp33_ASAP7_75t_L g506 ( 
.A1(n_448),
.A2(n_328),
.B(n_289),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_447),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

INVx6_ASAP7_75t_L g509 ( 
.A(n_427),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_427),
.B(n_258),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_446),
.B(n_292),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_403),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_446),
.B(n_292),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_446),
.B(n_315),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_437),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_434),
.B(n_315),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_434),
.B(n_268),
.Y(n_520)
);

BUFx6f_ASAP7_75t_SL g521 ( 
.A(n_413),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_444),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_417),
.Y(n_524)
);

AND2x6_ASAP7_75t_L g525 ( 
.A(n_444),
.B(n_268),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_419),
.B(n_296),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_431),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_431),
.B(n_315),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_451),
.A2(n_315),
.B1(n_304),
.B2(n_338),
.Y(n_529)
);

NAND2x1p5_ASAP7_75t_L g530 ( 
.A(n_403),
.B(n_262),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_451),
.B(n_315),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_459),
.B(n_413),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_463),
.A2(n_413),
.B(n_421),
.Y(n_533)
);

AO22x1_ASAP7_75t_L g534 ( 
.A1(n_526),
.A2(n_453),
.B1(n_429),
.B2(n_443),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_413),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_472),
.B(n_406),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_472),
.B(n_441),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_475),
.B(n_419),
.Y(n_538)
);

NOR3xp33_ASAP7_75t_L g539 ( 
.A(n_475),
.B(n_412),
.C(n_407),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_456),
.B(n_421),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_474),
.B(n_410),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_456),
.B(n_421),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_458),
.B(n_421),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_462),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_458),
.B(n_263),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_478),
.B(n_405),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_497),
.A2(n_436),
.B1(n_440),
.B2(n_397),
.Y(n_548)
);

O2A1O1Ixp5_ASAP7_75t_L g549 ( 
.A1(n_527),
.A2(n_522),
.B(n_511),
.C(n_517),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_512),
.B(n_315),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_493),
.B(n_264),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_493),
.B(n_265),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_484),
.B(n_463),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_483),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_457),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_513),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_490),
.B(n_417),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_501),
.B(n_424),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_461),
.B(n_270),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_424),
.Y(n_562)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_524),
.B(n_492),
.Y(n_563)
);

OR2x2_ASAP7_75t_SL g564 ( 
.A(n_470),
.B(n_442),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_467),
.B(n_428),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_465),
.B(n_428),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_529),
.A2(n_314),
.B1(n_278),
.B2(n_280),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_466),
.A2(n_452),
.B1(n_449),
.B2(n_320),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_473),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_479),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_L g571 ( 
.A(n_506),
.B(n_487),
.C(n_486),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_480),
.B(n_4),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_483),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_489),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_509),
.B(n_275),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_515),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_502),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_494),
.B(n_288),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_503),
.Y(n_579)
);

O2A1O1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_511),
.A2(n_452),
.B(n_449),
.C(n_440),
.Y(n_580)
);

O2A1O1Ixp5_ASAP7_75t_L g581 ( 
.A1(n_522),
.A2(n_295),
.B(n_297),
.C(n_300),
.Y(n_581)
);

O2A1O1Ixp5_ASAP7_75t_L g582 ( 
.A1(n_516),
.A2(n_301),
.B(n_302),
.C(n_303),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_461),
.B(n_310),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_481),
.B(n_311),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_481),
.B(n_316),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_496),
.B(n_326),
.Y(n_586)
);

NOR2x2_ASAP7_75t_L g587 ( 
.A(n_470),
.B(n_397),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

NAND2x1p5_ASAP7_75t_L g589 ( 
.A(n_512),
.B(n_45),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_500),
.B(n_327),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_507),
.B(n_331),
.Y(n_591)
);

INVx8_ASAP7_75t_L g592 ( 
.A(n_476),
.Y(n_592)
);

AO22x1_ASAP7_75t_L g593 ( 
.A1(n_468),
.A2(n_333),
.B1(n_335),
.B2(n_337),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_518),
.Y(n_594)
);

NAND3xp33_ASAP7_75t_L g595 ( 
.A(n_516),
.B(n_436),
.C(n_4),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_509),
.B(n_5),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_523),
.B(n_46),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_468),
.B(n_47),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_468),
.B(n_49),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_514),
.B(n_5),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_521),
.B(n_485),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_508),
.B(n_50),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_514),
.B(n_6),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_468),
.B(n_51),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_471),
.B(n_54),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_498),
.B(n_7),
.Y(n_607)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_517),
.A2(n_528),
.B(n_531),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_482),
.B(n_60),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_464),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_512),
.B(n_8),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_521),
.B(n_480),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_488),
.B(n_62),
.Y(n_614)
);

NOR2x1p5_ASAP7_75t_L g615 ( 
.A(n_531),
.B(n_9),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_562),
.B(n_530),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_599),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_592),
.Y(n_620)
);

A2O1A1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_542),
.A2(n_528),
.B(n_519),
.C(n_469),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_557),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_553),
.B(n_519),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_542),
.A2(n_530),
.B1(n_499),
.B2(n_495),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_469),
.Y(n_625)
);

AOI21xp33_ASAP7_75t_L g626 ( 
.A1(n_540),
.A2(n_477),
.B(n_464),
.Y(n_626)
);

INVx5_ASAP7_75t_L g627 ( 
.A(n_550),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_569),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_570),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_574),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_538),
.B(n_477),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_543),
.B(n_9),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_559),
.B(n_495),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_587),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_594),
.Y(n_635)
);

AND2x4_ASAP7_75t_SL g636 ( 
.A(n_539),
.B(n_63),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_609),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_564),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_608),
.B(n_495),
.Y(n_639)
);

AOI211xp5_ASAP7_75t_L g640 ( 
.A1(n_534),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_577),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_579),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_588),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_548),
.B(n_547),
.Y(n_645)
);

CKINVDCx8_ASAP7_75t_R g646 ( 
.A(n_592),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_576),
.Y(n_647)
);

AOI22x1_ASAP7_75t_L g648 ( 
.A1(n_541),
.A2(n_495),
.B1(n_520),
.B2(n_525),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_555),
.B(n_64),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_546),
.B(n_520),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_563),
.B(n_65),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_576),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_572),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_616),
.B(n_10),
.Y(n_655)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_550),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_568),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_545),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_544),
.B(n_12),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_558),
.B(n_520),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_SL g661 ( 
.A(n_595),
.B(n_580),
.C(n_604),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_554),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_612),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_537),
.B(n_13),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

NOR2x1_ASAP7_75t_L g666 ( 
.A(n_536),
.B(n_66),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_607),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_611),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_532),
.B(n_520),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_603),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_550),
.Y(n_671)
);

OR2x6_ASAP7_75t_L g672 ( 
.A(n_533),
.B(n_13),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_601),
.B(n_14),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_613),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_578),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_L g676 ( 
.A(n_550),
.B(n_525),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_R g677 ( 
.A(n_612),
.B(n_67),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_573),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_R g679 ( 
.A(n_535),
.B(n_68),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_578),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_571),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_571),
.Y(n_682)
);

NOR2x1_ASAP7_75t_L g683 ( 
.A(n_665),
.B(n_566),
.Y(n_683)
);

OAI21x1_ASAP7_75t_L g684 ( 
.A1(n_625),
.A2(n_549),
.B(n_606),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_617),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_623),
.B(n_561),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_663),
.A2(n_589),
.B1(n_596),
.B2(n_615),
.Y(n_687)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_663),
.A2(n_589),
.B1(n_596),
.B2(n_533),
.Y(n_688)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_646),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_L g690 ( 
.A1(n_621),
.A2(n_549),
.B(n_582),
.Y(n_690)
);

HB1xp67_ASAP7_75t_L g691 ( 
.A(n_654),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_664),
.A2(n_560),
.B(n_580),
.C(n_565),
.Y(n_692)
);

OAI21xp5_ASAP7_75t_L g693 ( 
.A1(n_625),
.A2(n_582),
.B(n_581),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_639),
.A2(n_614),
.B(n_610),
.Y(n_694)
);

OR2x2_ASAP7_75t_L g695 ( 
.A(n_634),
.B(n_584),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_L g696 ( 
.A(n_670),
.B(n_539),
.Y(n_696)
);

AOI21x1_ASAP7_75t_L g697 ( 
.A1(n_639),
.A2(n_583),
.B(n_552),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_631),
.B(n_551),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_654),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_622),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_620),
.B(n_575),
.Y(n_701)
);

OAI21x1_ASAP7_75t_SL g702 ( 
.A1(n_665),
.A2(n_666),
.B(n_681),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_670),
.Y(n_703)
);

AOI21x1_ASAP7_75t_SL g704 ( 
.A1(n_652),
.A2(n_600),
.B(n_598),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_623),
.B(n_550),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_682),
.B(n_575),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_651),
.A2(n_597),
.B(n_581),
.Y(n_707)
);

AO31x2_ASAP7_75t_L g708 ( 
.A1(n_632),
.A2(n_567),
.A3(n_605),
.B(n_591),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_627),
.A2(n_585),
.B(n_586),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_632),
.B(n_590),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_659),
.B(n_590),
.Y(n_711)
);

NAND2x1_ASAP7_75t_L g712 ( 
.A(n_670),
.B(n_525),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_651),
.A2(n_593),
.B(n_123),
.Y(n_713)
);

OAI21x1_ASAP7_75t_L g714 ( 
.A1(n_669),
.A2(n_668),
.B(n_637),
.Y(n_714)
);

OAI21x1_ASAP7_75t_SL g715 ( 
.A1(n_626),
.A2(n_121),
.B(n_237),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_659),
.B(n_618),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_628),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_619),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_664),
.B(n_525),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_14),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_667),
.B(n_15),
.Y(n_722)
);

BUFx2_ASAP7_75t_L g723 ( 
.A(n_638),
.Y(n_723)
);

INVx3_ASAP7_75t_SL g724 ( 
.A(n_655),
.Y(n_724)
);

OAI21xp5_ASAP7_75t_L g725 ( 
.A1(n_626),
.A2(n_624),
.B(n_660),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_627),
.B(n_71),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_630),
.B(n_72),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_637),
.A2(n_127),
.B(n_231),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_627),
.Y(n_729)
);

AO31x2_ASAP7_75t_L g730 ( 
.A1(n_635),
.A2(n_16),
.A3(n_17),
.B(n_18),
.Y(n_730)
);

AO31x2_ASAP7_75t_L g731 ( 
.A1(n_662),
.A2(n_16),
.A3(n_18),
.B(n_19),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_649),
.Y(n_732)
);

BUFx4f_ASAP7_75t_SL g733 ( 
.A(n_620),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_680),
.B(n_20),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_673),
.B(n_22),
.Y(n_735)
);

OAI21x1_ASAP7_75t_L g736 ( 
.A1(n_668),
.A2(n_132),
.B(n_230),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_641),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_648),
.A2(n_678),
.B(n_658),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_675),
.B(n_75),
.Y(n_739)
);

AOI21x1_ASAP7_75t_L g740 ( 
.A1(n_653),
.A2(n_133),
.B(n_226),
.Y(n_740)
);

OAI21xp5_ASAP7_75t_L g741 ( 
.A1(n_661),
.A2(n_129),
.B(n_225),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_661),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_742)
);

AO21x2_ASAP7_75t_L g743 ( 
.A1(n_693),
.A2(n_677),
.B(n_679),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_705),
.A2(n_642),
.B(n_644),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

OAI21x1_ASAP7_75t_L g746 ( 
.A1(n_738),
.A2(n_647),
.B(n_633),
.Y(n_746)
);

OAI21x1_ASAP7_75t_L g747 ( 
.A1(n_714),
.A2(n_627),
.B(n_656),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_700),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_742),
.A2(n_672),
.B1(n_657),
.B2(n_655),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_718),
.Y(n_750)
);

OAI21x1_ASAP7_75t_L g751 ( 
.A1(n_704),
.A2(n_656),
.B(n_671),
.Y(n_751)
);

AOI22xp5_ASAP7_75t_L g752 ( 
.A1(n_696),
.A2(n_645),
.B1(n_636),
.B2(n_652),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_716),
.A2(n_656),
.B1(n_671),
.B2(n_672),
.Y(n_753)
);

OAI21x1_ASAP7_75t_L g754 ( 
.A1(n_684),
.A2(n_671),
.B(n_656),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_737),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_732),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_719),
.Y(n_757)
);

OAI22xp33_ASAP7_75t_L g758 ( 
.A1(n_742),
.A2(n_672),
.B1(n_655),
.B2(n_671),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_697),
.A2(n_676),
.B(n_679),
.Y(n_759)
);

NOR2xp67_ASAP7_75t_L g760 ( 
.A(n_695),
.B(n_643),
.Y(n_760)
);

OAI21xp5_ASAP7_75t_L g761 ( 
.A1(n_705),
.A2(n_650),
.B(n_640),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_698),
.A2(n_650),
.B(n_677),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_729),
.B(n_643),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_703),
.B(n_643),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_721),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_741),
.A2(n_674),
.B1(n_649),
.B2(n_26),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_SL g767 ( 
.A1(n_741),
.A2(n_674),
.B(n_25),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_710),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_691),
.Y(n_769)
);

INVx1_ASAP7_75t_SL g770 ( 
.A(n_723),
.Y(n_770)
);

OA21x2_ASAP7_75t_L g771 ( 
.A1(n_693),
.A2(n_27),
.B(n_28),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_699),
.Y(n_772)
);

AO31x2_ASAP7_75t_L g773 ( 
.A1(n_688),
.A2(n_27),
.A3(n_28),
.B(n_29),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_727),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_706),
.A2(n_143),
.B(n_221),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_694),
.A2(n_141),
.B(n_218),
.Y(n_776)
);

AO21x2_ASAP7_75t_L g777 ( 
.A1(n_690),
.A2(n_139),
.B(n_217),
.Y(n_777)
);

OAI21x1_ASAP7_75t_L g778 ( 
.A1(n_713),
.A2(n_126),
.B(n_216),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_703),
.B(n_77),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_686),
.B(n_29),
.Y(n_780)
);

AO31x2_ASAP7_75t_L g781 ( 
.A1(n_688),
.A2(n_30),
.A3(n_31),
.B(n_32),
.Y(n_781)
);

NAND2x1p5_ASAP7_75t_L g782 ( 
.A(n_729),
.B(n_80),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_686),
.B(n_30),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_727),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_716),
.A2(n_146),
.B(n_215),
.Y(n_785)
);

CKINVDCx6p67_ASAP7_75t_R g786 ( 
.A(n_724),
.Y(n_786)
);

OAI21x1_ASAP7_75t_L g787 ( 
.A1(n_707),
.A2(n_145),
.B(n_214),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_729),
.Y(n_788)
);

OAI21x1_ASAP7_75t_L g789 ( 
.A1(n_728),
.A2(n_118),
.B(n_213),
.Y(n_789)
);

CKINVDCx11_ASAP7_75t_R g790 ( 
.A(n_689),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_711),
.B(n_735),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_729),
.Y(n_792)
);

AO31x2_ASAP7_75t_L g793 ( 
.A1(n_687),
.A2(n_31),
.A3(n_32),
.B(n_33),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_717),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_722),
.B(n_33),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_687),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_R g797 ( 
.A(n_756),
.B(n_701),
.Y(n_797)
);

AND2x4_ASAP7_75t_L g798 ( 
.A(n_764),
.B(n_739),
.Y(n_798)
);

INVx3_ASAP7_75t_L g799 ( 
.A(n_763),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_752),
.A2(n_683),
.B1(n_739),
.B2(n_734),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_745),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_774),
.B(n_692),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_770),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_745),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_756),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_769),
.Y(n_806)
);

A2O1A1Ixp33_ASAP7_75t_L g807 ( 
.A1(n_767),
.A2(n_766),
.B(n_762),
.C(n_765),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_766),
.A2(n_715),
.B1(n_702),
.B2(n_725),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_790),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_763),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_749),
.A2(n_720),
.B(n_725),
.C(n_726),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_755),
.Y(n_812)
);

OR2x6_ASAP7_75t_L g813 ( 
.A(n_782),
.B(n_736),
.Y(n_813)
);

AO32x2_ASAP7_75t_L g814 ( 
.A1(n_796),
.A2(n_731),
.A3(n_730),
.B1(n_690),
.B2(n_708),
.Y(n_814)
);

AND2x4_ASAP7_75t_L g815 ( 
.A(n_764),
.B(n_717),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_743),
.A2(n_709),
.B(n_712),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_794),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_749),
.A2(n_758),
.B1(n_761),
.B2(n_785),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_758),
.A2(n_717),
.B1(n_733),
.B2(n_708),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_791),
.A2(n_708),
.B1(n_731),
.B2(n_740),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_743),
.A2(n_730),
.B(n_149),
.Y(n_821)
);

BUFx2_ASAP7_75t_L g822 ( 
.A(n_794),
.Y(n_822)
);

BUFx4f_ASAP7_75t_SL g823 ( 
.A(n_786),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_755),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_746),
.A2(n_730),
.B(n_731),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_784),
.B(n_780),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_744),
.A2(n_783),
.B(n_775),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_760),
.B(n_34),
.Y(n_828)
);

CKINVDCx6p67_ASAP7_75t_R g829 ( 
.A(n_790),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_764),
.B(n_81),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_748),
.Y(n_831)
);

CKINVDCx20_ASAP7_75t_R g832 ( 
.A(n_795),
.Y(n_832)
);

AO31x2_ASAP7_75t_L g833 ( 
.A1(n_753),
.A2(n_35),
.A3(n_36),
.B(n_37),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_750),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_757),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_773),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_772),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_773),
.Y(n_838)
);

NOR2x1_ASAP7_75t_SL g839 ( 
.A(n_777),
.B(n_83),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_792),
.Y(n_840)
);

OAI21x1_ASAP7_75t_L g841 ( 
.A1(n_754),
.A2(n_155),
.B(n_212),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_768),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_792),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_773),
.B(n_38),
.Y(n_844)
);

OAI221xp5_ASAP7_75t_L g845 ( 
.A1(n_771),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.C(n_84),
.Y(n_845)
);

OR2x6_ASAP7_75t_L g846 ( 
.A(n_782),
.B(n_157),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_779),
.B(n_161),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_773),
.B(n_42),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_788),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_751),
.B(n_162),
.Y(n_850)
);

INVx6_ASAP7_75t_L g851 ( 
.A(n_779),
.Y(n_851)
);

AOI221xp5_ASAP7_75t_L g852 ( 
.A1(n_777),
.A2(n_43),
.B1(n_85),
.B2(n_86),
.C(n_87),
.Y(n_852)
);

OAI22xp33_ASAP7_75t_L g853 ( 
.A1(n_771),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_781),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_781),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_779),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_842),
.A2(n_771),
.B1(n_793),
.B2(n_789),
.Y(n_857)
);

BUFx6f_ASAP7_75t_L g858 ( 
.A(n_815),
.Y(n_858)
);

NOR2x1_ASAP7_75t_SL g859 ( 
.A(n_850),
.B(n_781),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_826),
.B(n_793),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_840),
.B(n_793),
.Y(n_861)
);

AOI222xp33_ASAP7_75t_L g862 ( 
.A1(n_818),
.A2(n_793),
.B1(n_781),
.B2(n_788),
.C1(n_789),
.C2(n_787),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_827),
.A2(n_776),
.B1(n_759),
.B2(n_778),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_804),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_834),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_800),
.A2(n_778),
.B1(n_747),
.B2(n_97),
.Y(n_866)
);

OAI21x1_ASAP7_75t_L g867 ( 
.A1(n_816),
.A2(n_92),
.B(n_94),
.Y(n_867)
);

BUFx2_ASAP7_75t_L g868 ( 
.A(n_803),
.Y(n_868)
);

OAI211xp5_ASAP7_75t_L g869 ( 
.A1(n_845),
.A2(n_98),
.B(n_99),
.C(n_100),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_SL g870 ( 
.A1(n_845),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_826),
.B(n_104),
.Y(n_871)
);

AOI21xp33_ASAP7_75t_L g872 ( 
.A1(n_827),
.A2(n_105),
.B(n_108),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_852),
.A2(n_109),
.B1(n_111),
.B2(n_113),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_SL g874 ( 
.A1(n_839),
.A2(n_846),
.B1(n_851),
.B2(n_847),
.Y(n_874)
);

OAI21x1_ASAP7_75t_SL g875 ( 
.A1(n_811),
.A2(n_114),
.B(n_115),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_846),
.A2(n_116),
.B1(n_147),
.B2(n_148),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_SL g877 ( 
.A1(n_846),
.A2(n_152),
.B1(n_156),
.B2(n_165),
.Y(n_877)
);

OAI22xp33_ASAP7_75t_L g878 ( 
.A1(n_852),
.A2(n_166),
.B1(n_170),
.B2(n_171),
.Y(n_878)
);

OAI221xp5_ASAP7_75t_L g879 ( 
.A1(n_807),
.A2(n_808),
.B1(n_819),
.B2(n_828),
.C(n_802),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_856),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_843),
.B(n_824),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_812),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_801),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_831),
.Y(n_884)
);

AND2x2_ASAP7_75t_L g885 ( 
.A(n_856),
.B(n_798),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_851),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_832),
.A2(n_235),
.B1(n_178),
.B2(n_180),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_798),
.B(n_177),
.Y(n_888)
);

INVxp67_ASAP7_75t_R g889 ( 
.A(n_806),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_849),
.Y(n_890)
);

AO21x2_ASAP7_75t_L g891 ( 
.A1(n_821),
.A2(n_183),
.B(n_186),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_835),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_825),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_815),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_802),
.A2(n_208),
.B1(n_191),
.B2(n_192),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_797),
.A2(n_187),
.B1(n_193),
.B2(n_194),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_847),
.B(n_195),
.Y(n_897)
);

OAI22xp33_ASAP7_75t_L g898 ( 
.A1(n_844),
.A2(n_196),
.B1(n_197),
.B2(n_201),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_841),
.A2(n_202),
.B(n_203),
.Y(n_899)
);

OAI211xp5_ASAP7_75t_L g900 ( 
.A1(n_844),
.A2(n_848),
.B(n_820),
.C(n_836),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_817),
.B(n_204),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_848),
.Y(n_902)
);

AOI21xp33_ASAP7_75t_L g903 ( 
.A1(n_853),
.A2(n_205),
.B(n_206),
.Y(n_903)
);

OAI221xp5_ASAP7_75t_L g904 ( 
.A1(n_837),
.A2(n_805),
.B1(n_809),
.B2(n_813),
.C(n_850),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_SL g905 ( 
.A1(n_830),
.A2(n_823),
.B1(n_850),
.B2(n_813),
.Y(n_905)
);

AO31x2_ASAP7_75t_L g906 ( 
.A1(n_838),
.A2(n_855),
.A3(n_854),
.B(n_814),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_906),
.B(n_814),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_906),
.Y(n_908)
);

HB1xp67_ASAP7_75t_L g909 ( 
.A(n_906),
.Y(n_909)
);

AND2x2_ASAP7_75t_L g910 ( 
.A(n_906),
.B(n_814),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_893),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_902),
.Y(n_912)
);

INVx4_ASAP7_75t_L g913 ( 
.A(n_891),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_860),
.B(n_833),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_861),
.B(n_833),
.Y(n_915)
);

AND2x4_ASAP7_75t_L g916 ( 
.A(n_893),
.B(n_813),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_865),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_864),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_882),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_859),
.B(n_833),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_883),
.B(n_849),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_892),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_868),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_883),
.Y(n_925)
);

OAI31xp33_ASAP7_75t_L g926 ( 
.A1(n_878),
.A2(n_869),
.A3(n_898),
.B(n_879),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_884),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_881),
.Y(n_928)
);

OR2x2_ASAP7_75t_L g929 ( 
.A(n_900),
.B(n_822),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_867),
.Y(n_930)
);

INVxp67_ASAP7_75t_R g931 ( 
.A(n_867),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_862),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_890),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_899),
.Y(n_934)
);

OAI21x1_ASAP7_75t_L g935 ( 
.A1(n_863),
.A2(n_799),
.B(n_810),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_890),
.Y(n_936)
);

BUFx3_ASAP7_75t_L g937 ( 
.A(n_904),
.Y(n_937)
);

NOR2xp67_ASAP7_75t_SL g938 ( 
.A(n_878),
.B(n_799),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_899),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_898),
.B(n_810),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_891),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_871),
.B(n_829),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_924),
.B(n_885),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_914),
.B(n_857),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_924),
.Y(n_945)
);

NAND2x1p5_ASAP7_75t_L g946 ( 
.A(n_929),
.B(n_886),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

OAI22xp5_ASAP7_75t_L g948 ( 
.A1(n_937),
.A2(n_873),
.B1(n_870),
.B2(n_905),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_917),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_924),
.B(n_889),
.Y(n_950)
);

NOR4xp25_ASAP7_75t_SL g951 ( 
.A(n_932),
.B(n_872),
.C(n_903),
.D(n_873),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_923),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_938),
.A2(n_874),
.B1(n_887),
.B2(n_896),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_926),
.A2(n_887),
.B1(n_895),
.B2(n_877),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_935),
.B(n_921),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_914),
.B(n_857),
.Y(n_956)
);

AO21x2_ASAP7_75t_L g957 ( 
.A1(n_939),
.A2(n_930),
.B(n_932),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_937),
.B(n_894),
.Y(n_958)
);

AOI22xp33_ASAP7_75t_SL g959 ( 
.A1(n_937),
.A2(n_866),
.B1(n_875),
.B2(n_880),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_936),
.B(n_894),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_908),
.Y(n_961)
);

AOI22xp33_ASAP7_75t_SL g962 ( 
.A1(n_940),
.A2(n_897),
.B1(n_830),
.B2(n_888),
.Y(n_962)
);

OAI211xp5_ASAP7_75t_L g963 ( 
.A1(n_926),
.A2(n_895),
.B(n_876),
.C(n_863),
.Y(n_963)
);

OAI221xp5_ASAP7_75t_L g964 ( 
.A1(n_942),
.A2(n_858),
.B1(n_886),
.B2(n_901),
.C(n_940),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_936),
.Y(n_965)
);

OAI33xp33_ASAP7_75t_L g966 ( 
.A1(n_912),
.A2(n_858),
.A3(n_927),
.B1(n_929),
.B2(n_923),
.B3(n_933),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_936),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_965),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_955),
.B(n_921),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_947),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_949),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_957),
.B(n_915),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_957),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_952),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_955),
.B(n_945),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_967),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_961),
.Y(n_977)
);

OR2x2_ASAP7_75t_L g978 ( 
.A(n_944),
.B(n_915),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_955),
.B(n_921),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_961),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_946),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_960),
.B(n_916),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_946),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_970),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_971),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_974),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_973),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_978),
.A2(n_954),
.B1(n_953),
.B2(n_948),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_980),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_980),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_977),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_968),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_982),
.B(n_975),
.Y(n_993)
);

AO21x1_ASAP7_75t_L g994 ( 
.A1(n_988),
.A2(n_972),
.B(n_913),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_989),
.B(n_978),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_984),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_987),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_993),
.B(n_975),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_990),
.B(n_985),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_987),
.Y(n_1000)
);

AND2x2_ASAP7_75t_L g1001 ( 
.A(n_991),
.B(n_982),
.Y(n_1001)
);

AOI22x1_ASAP7_75t_L g1002 ( 
.A1(n_986),
.A2(n_983),
.B1(n_972),
.B2(n_981),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_1002),
.A2(n_988),
.B1(n_954),
.B2(n_964),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_996),
.B(n_992),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_999),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_999),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_997),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_1007),
.Y(n_1008)
);

INVxp67_ASAP7_75t_SL g1009 ( 
.A(n_1006),
.Y(n_1009)
);

NOR2x1_ASAP7_75t_L g1010 ( 
.A(n_1003),
.B(n_997),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_SL g1011 ( 
.A1(n_1009),
.A2(n_1005),
.B(n_1004),
.C(n_1000),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_1010),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_1008),
.B(n_1001),
.Y(n_1013)
);

AOI211xp5_ASAP7_75t_L g1014 ( 
.A1(n_1009),
.A2(n_994),
.B(n_963),
.C(n_942),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_1012),
.B(n_951),
.C(n_959),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_1014),
.B(n_998),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1013),
.A2(n_995),
.B1(n_969),
.B2(n_979),
.Y(n_1017)
);

AOI211xp5_ASAP7_75t_L g1018 ( 
.A1(n_1011),
.A2(n_938),
.B(n_958),
.C(n_995),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_1012),
.A2(n_959),
.B(n_958),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_1012),
.B(n_979),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_1012),
.B(n_969),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_1012),
.B(n_983),
.Y(n_1022)
);

OAI221xp5_ASAP7_75t_SL g1023 ( 
.A1(n_1018),
.A2(n_956),
.B1(n_950),
.B2(n_929),
.C(n_962),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1020),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_1016),
.B(n_976),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_SL g1026 ( 
.A(n_1015),
.B(n_1022),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_SL g1027 ( 
.A1(n_1019),
.A2(n_913),
.B1(n_941),
.B2(n_915),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_1021),
.B(n_966),
.Y(n_1028)
);

AOI22xp33_ASAP7_75t_L g1029 ( 
.A1(n_1017),
.A2(n_913),
.B1(n_938),
.B2(n_941),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1024),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_1025),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1028),
.Y(n_1032)
);

OAI21xp33_ASAP7_75t_L g1033 ( 
.A1(n_1026),
.A2(n_962),
.B(n_943),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1023),
.A2(n_976),
.B1(n_968),
.B2(n_982),
.Y(n_1034)
);

AO22x2_ASAP7_75t_L g1035 ( 
.A1(n_1027),
.A2(n_913),
.B1(n_941),
.B2(n_933),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_1029),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_1032),
.B(n_966),
.C(n_913),
.Y(n_1037)
);

NAND4xp75_ASAP7_75t_L g1038 ( 
.A(n_1030),
.B(n_927),
.C(n_912),
.D(n_939),
.Y(n_1038)
);

AND3x4_ASAP7_75t_L g1039 ( 
.A(n_1036),
.B(n_960),
.C(n_916),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_1033),
.A2(n_941),
.B1(n_858),
.B2(n_931),
.Y(n_1040)
);

OAI21xp33_ASAP7_75t_L g1041 ( 
.A1(n_1031),
.A2(n_928),
.B(n_941),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1034),
.B(n_928),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1035),
.B(n_858),
.Y(n_1043)
);

NOR2xp67_ASAP7_75t_L g1044 ( 
.A(n_1040),
.B(n_1035),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1039),
.Y(n_1045)
);

NAND3xp33_ASAP7_75t_L g1046 ( 
.A(n_1042),
.B(n_930),
.C(n_934),
.Y(n_1046)
);

NOR4xp25_ASAP7_75t_L g1047 ( 
.A(n_1041),
.B(n_934),
.C(n_930),
.D(n_920),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_922),
.Y(n_1048)
);

XNOR2x1_ASAP7_75t_L g1049 ( 
.A(n_1038),
.B(n_935),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1045),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_1044),
.B(n_1037),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1048),
.B(n_920),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1046),
.Y(n_1053)
);

NAND3x1_ASAP7_75t_L g1054 ( 
.A(n_1051),
.B(n_1049),
.C(n_1047),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_1050),
.B(n_934),
.Y(n_1055)
);

AOI31xp33_ASAP7_75t_L g1056 ( 
.A1(n_1053),
.A2(n_920),
.A3(n_922),
.B(n_909),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_1052),
.Y(n_1057)
);

AOI21xp33_ASAP7_75t_L g1058 ( 
.A1(n_1057),
.A2(n_934),
.B(n_916),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_1054),
.A2(n_908),
.B1(n_909),
.B2(n_934),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1059),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_1058),
.B(n_1055),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_SL g1062 ( 
.A1(n_1060),
.A2(n_1056),
.B1(n_922),
.B2(n_916),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1061),
.A2(n_931),
.B(n_922),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1062),
.A2(n_1063),
.B(n_931),
.Y(n_1064)
);

AOI222xp33_ASAP7_75t_L g1065 ( 
.A1(n_1062),
.A2(n_916),
.B1(n_922),
.B2(n_907),
.C1(n_910),
.C2(n_918),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1065),
.B1(n_925),
.B2(n_919),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_SL g1067 ( 
.A1(n_1064),
.A2(n_925),
.B1(n_935),
.B2(n_918),
.Y(n_1067)
);

OAI221xp5_ASAP7_75t_R g1068 ( 
.A1(n_1067),
.A2(n_925),
.B1(n_910),
.B2(n_907),
.C(n_918),
.Y(n_1068)
);

AOI211xp5_ASAP7_75t_L g1069 ( 
.A1(n_1068),
.A2(n_1066),
.B(n_919),
.C(n_911),
.Y(n_1069)
);


endmodule