module fake_jpeg_16554_n_292 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_292);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_292;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_38),
.Y(n_52)
);

BUFx2_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_43),
.Y(n_62)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_44),
.B1(n_35),
.B2(n_28),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_38),
.B1(n_41),
.B2(n_40),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_21),
.B1(n_28),
.B2(n_29),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_51),
.B(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_29),
.B1(n_43),
.B2(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_24),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_40),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_18),
.B1(n_19),
.B2(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_85)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_23),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_36),
.Y(n_65)
);

NAND2x1_ASAP7_75t_SL g67 ( 
.A(n_47),
.B(n_34),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_67),
.A2(n_94),
.B(n_5),
.C(n_7),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_36),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_69),
.B(n_80),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_70),
.A2(n_91),
.B1(n_100),
.B2(n_57),
.Y(n_106)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

O2A1O1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_38),
.B(n_32),
.C(n_17),
.Y(n_74)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_41),
.B(n_61),
.C(n_58),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_75),
.B(n_79),
.Y(n_127)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_77),
.B(n_81),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_92),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_50),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_60),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_82),
.B(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_22),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_83),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_56),
.B(n_22),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_34),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_53),
.B(n_24),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_47),
.A2(n_39),
.B(n_1),
.C(n_2),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_49),
.A2(n_38),
.B1(n_31),
.B2(n_30),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_95),
.A2(n_102),
.B1(n_58),
.B2(n_9),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_61),
.Y(n_108)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_53),
.B(n_0),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_41),
.B1(n_31),
.B2(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_103),
.Y(n_129)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_39),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_39),
.C(n_41),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_128),
.C(n_130),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_118),
.B1(n_70),
.B2(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_108),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_109),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_1),
.B(n_4),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_114),
.B(n_115),
.Y(n_138)
);

AND2x6_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_4),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_65),
.B(n_5),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_72),
.B(n_16),
.C(n_9),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_66),
.C(n_84),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_124),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_133),
.B(n_142),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_104),
.B(n_78),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_134),
.A2(n_136),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_123),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_156),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_78),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_137),
.B(n_139),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_81),
.Y(n_140)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_141),
.A2(n_100),
.B1(n_128),
.B2(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_80),
.Y(n_144)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_144),
.Y(n_174)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_120),
.A2(n_85),
.B(n_94),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_154),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_85),
.B1(n_66),
.B2(n_91),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_114),
.B1(n_117),
.B2(n_106),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_97),
.B1(n_68),
.B2(n_73),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_152),
.A2(n_73),
.B1(n_102),
.B2(n_88),
.Y(n_189)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_74),
.B(n_67),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_115),
.B(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_68),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_135),
.B(n_125),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_161),
.B(n_189),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_163),
.A2(n_167),
.B(n_133),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_153),
.B(n_111),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_170),
.C(n_172),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_107),
.B(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_107),
.C(n_131),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_107),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_158),
.A2(n_122),
.B1(n_117),
.B2(n_113),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_180),
.B1(n_187),
.B2(n_188),
.Y(n_196)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

INVxp67_ASAP7_75t_SL g198 ( 
.A(n_176),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_90),
.C(n_132),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_182),
.C(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_126),
.Y(n_179)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_179),
.Y(n_213)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_149),
.A2(n_110),
.B1(n_122),
.B2(n_117),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_184),
.B1(n_146),
.B2(n_154),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_134),
.B(n_136),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_143),
.B(n_126),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_145),
.A2(n_67),
.B1(n_76),
.B2(n_116),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_136),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_173),
.B(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_197),
.C(n_172),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_194),
.A2(n_204),
.B(n_167),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_206),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g200 ( 
.A(n_173),
.B(n_138),
.C(n_155),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_200),
.B(n_182),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_147),
.Y(n_201)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_138),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_202),
.Y(n_214)
);

OAI22x1_ASAP7_75t_SL g205 ( 
.A1(n_180),
.A2(n_155),
.B1(n_137),
.B2(n_139),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_171),
.B1(n_178),
.B2(n_164),
.Y(n_215)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_183),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_210),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_176),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_98),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_211),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_186),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_212),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_227),
.B1(n_203),
.B2(n_206),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_231),
.B(n_8),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g219 ( 
.A(n_205),
.B(n_185),
.C(n_175),
.Y(n_219)
);

NAND3xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_196),
.C(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_197),
.C(n_195),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_77),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_171),
.B1(n_177),
.B2(n_170),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_163),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_230),
.B(n_196),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_202),
.A2(n_181),
.B(n_188),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_189),
.B1(n_165),
.B2(n_77),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_222),
.C(n_225),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

OAI322xp33_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_190),
.A3(n_192),
.B1(n_213),
.B2(n_193),
.C1(n_203),
.C2(n_211),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_243),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_218),
.A2(n_194),
.B(n_213),
.Y(n_236)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

BUFx12_ASAP7_75t_L g237 ( 
.A(n_226),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_241),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_240),
.Y(n_261)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_249),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_191),
.A3(n_195),
.B1(n_198),
.B2(n_210),
.C(n_96),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_244),
.A2(n_247),
.B1(n_248),
.B2(n_223),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_232),
.C(n_229),
.Y(n_252)
);

OA21x2_ASAP7_75t_SL g248 ( 
.A1(n_219),
.A2(n_9),
.B(n_10),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_16),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_251),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_215),
.C(n_227),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_247),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_214),
.C(n_221),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_260),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_214),
.C(n_223),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_263),
.B(n_268),
.Y(n_276)
);

AOI211xp5_ASAP7_75t_SL g266 ( 
.A1(n_258),
.A2(n_236),
.B(n_259),
.C(n_254),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_245),
.C(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_237),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_270),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_245),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_229),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_269),
.B(n_249),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_237),
.Y(n_270)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_257),
.Y(n_272)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_272),
.A2(n_274),
.B(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_217),
.Y(n_281)
);

NOR2x1_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_228),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_217),
.B1(n_261),
.B2(n_240),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_268),
.C(n_263),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_14),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_278),
.A2(n_271),
.B(n_240),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_11),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_283),
.B(n_15),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_10),
.C(n_11),
.Y(n_283)
);

AOI322xp5_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_273),
.A3(n_276),
.B1(n_12),
.B2(n_13),
.C1(n_10),
.C2(n_15),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_286),
.B(n_287),
.Y(n_289)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_289),
.B(n_14),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_14),
.Y(n_292)
);


endmodule