module real_jpeg_4274_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_0),
.B(n_124),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_0),
.B(n_177),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_0),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_0),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_0),
.B(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_0),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_0),
.B(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_1),
.Y(n_97)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_1),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_1),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_1),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_1),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_1),
.Y(n_313)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_2),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_2),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_2),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_3),
.B(n_179),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_3),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_3),
.B(n_293),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_3),
.B(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_3),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_3),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_3),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_4),
.B(n_32),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_4),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_4),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_4),
.B(n_221),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_4),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_4),
.B(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_5),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_5),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_47),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_5),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_5),
.B(n_296),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_5),
.B(n_400),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_6),
.Y(n_94)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_6),
.Y(n_116)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_6),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g385 ( 
.A(n_6),
.Y(n_385)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_7),
.Y(n_483)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_10),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_10),
.Y(n_214)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_12),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_12),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_12),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_12),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_13),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_13),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_13),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_13),
.B(n_81),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_14),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_14),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_14),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_14),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_14),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_14),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_14),
.B(n_358),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_14),
.B(n_221),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_15),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_16),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_16),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_16),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_16),
.B(n_274),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_16),
.B(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_16),
.B(n_369),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_16),
.B(n_385),
.Y(n_384)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_18),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_18),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_18),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_18),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_18),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_18),
.B(n_270),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_18),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_19),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_19),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_19),
.B(n_84),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_19),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g215 ( 
.A(n_19),
.B(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_481),
.B(n_484),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_182),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_181),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_143),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_25),
.B(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_104),
.B2(n_142),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_73),
.C(n_88),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_28),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_45),
.C(n_59),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_29),
.A2(n_30),
.B1(n_45),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_31),
.B(n_36),
.C(n_41),
.Y(n_118)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_40),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_40),
.Y(n_373)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_40),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_44),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_44),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g395 ( 
.A(n_44),
.Y(n_395)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_45),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.C(n_54),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_46),
.B(n_54),
.Y(n_163)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_50),
.B(n_163),
.Y(n_162)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_58),
.Y(n_173)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_58),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_58),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_59),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_66),
.C(n_69),
.Y(n_117)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_63),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_69),
.B2(n_72),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_66),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_108),
.C(n_112),
.Y(n_129)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_68),
.Y(n_271)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_68),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_91),
.C(n_95),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_69),
.A2(n_72),
.B1(n_95),
.B2(n_96),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g257 ( 
.A(n_71),
.Y(n_257)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_71),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_73),
.A2(n_88),
.B1(n_89),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_79),
.C(n_87),
.Y(n_127)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_83),
.B2(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_82),
.Y(n_342)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_86),
.Y(n_280)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_86),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_86),
.Y(n_383)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_101),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_90),
.B(n_165),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_91),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_95),
.A2(n_96),
.B1(n_158),
.B2(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_154),
.C(n_158),
.Y(n_153)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_97),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_102),
.Y(n_165)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_101),
.A2(n_102),
.B1(n_175),
.B2(n_176),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_102),
.B(n_167),
.C(n_175),
.Y(n_166)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_103),
.Y(n_250)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_119),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_117),
.C(n_118),
.Y(n_105)
);

FAx1_ASAP7_75t_SL g148 ( 
.A(n_106),
.B(n_117),
.CI(n_118),
.CON(n_148),
.SN(n_148)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_109),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_114),
.Y(n_254)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_128),
.B2(n_141),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_127),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_139),
.B2(n_140),
.Y(n_128)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_129),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_138),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_148),
.C(n_149),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_144),
.A2(n_145),
.B1(n_148),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_148),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_148),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_149),
.B(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.C(n_166),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_150),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_162),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_151),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_153),
.B(n_162),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_158),
.Y(n_204)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx8_ASAP7_75t_L g358 ( 
.A(n_160),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_161),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_164),
.B(n_166),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.C(n_174),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_174),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_189),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AO21x1_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_473),
.B(n_479),
.Y(n_182)
);

OAI21x1_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_281),
.B(n_472),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_232),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_185),
.B(n_232),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_226),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_186),
.B(n_227),
.C(n_230),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_205),
.C(n_207),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_187),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_202),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_188),
.B(n_458),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_190),
.A2(n_191),
.B1(n_202),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.C(n_198),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_192),
.B(n_198),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_193),
.B(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_200),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_202),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_205),
.B(n_207),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_220),
.C(n_222),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_208),
.B(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.C(n_215),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_209),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_215),
.Y(n_244)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_220),
.B(n_222),
.Y(n_262)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_239),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_234),
.B(n_237),
.Y(n_468)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_239),
.B(n_468),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_260),
.C(n_263),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_241),
.B(n_461),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_242),
.A2(n_243),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_245),
.A2(n_246),
.B(n_248),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_245),
.B(n_251),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_258),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_416)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_258),
.B(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_259),
.B(n_271),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_260),
.A2(n_261),
.B1(n_263),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_263),
.Y(n_462)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_276),
.C(n_277),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_265),
.B(n_450),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_269),
.C(n_272),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_266),
.B(n_428),
.Y(n_427)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_269),
.A2(n_272),
.B1(n_273),
.B2(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g429 ( 
.A(n_269),
.Y(n_429)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_276),
.B(n_277),
.Y(n_450)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI21x1_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_466),
.B(n_471),
.Y(n_281)
);

OAI21x1_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_453),
.B(n_465),
.Y(n_282)
);

AOI21x1_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_435),
.B(n_452),
.Y(n_283)
);

OAI21x1_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_409),
.B(n_434),
.Y(n_284)
);

AOI21x1_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_377),
.B(n_408),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_346),
.B(n_376),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_324),
.B(n_345),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_303),
.B(n_323),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_299),
.B(n_302),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_297),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_297),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_295),
.Y(n_304)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g404 ( 
.A(n_301),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_305),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_314),
.B2(n_315),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_306),
.B(n_317),
.C(n_321),
.Y(n_344)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_312),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_312),
.Y(n_335)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_321),
.B2(n_322),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_344),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_344),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_336),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_335),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_327),
.B(n_335),
.C(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_332),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_332),
.Y(n_351)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_337),
.B(n_362),
.C(n_363),
.Y(n_361)
);

INVx5_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_341),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_343),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_349),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_360),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_350),
.B(n_361),
.C(n_364),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_351),
.B(n_353),
.C(n_354),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_359),
.Y(n_354)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_355),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_359),
.Y(n_386)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_367),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g406 ( 
.A(n_365),
.B(n_371),
.C(n_374),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_371),
.B1(n_374),
.B2(n_375),
.Y(n_367)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_371),
.Y(n_375)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_378),
.B(n_407),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_407),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_388),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_387),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_380),
.B(n_387),
.C(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_386),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_384),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_423),
.C(n_424),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_388),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_396),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_389),
.B(n_398),
.C(n_405),
.Y(n_412)
);

BUFx24_ASAP7_75t_SL g488 ( 
.A(n_389),
.Y(n_488)
);

FAx1_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_392),
.CI(n_393),
.CON(n_389),
.SN(n_389)
);

MAJx2_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_392),
.C(n_393),
.Y(n_420)
);

INVx3_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_405),
.B2(n_406),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_399),
.B(n_402),
.Y(n_419)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx3_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_432),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_432),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_421),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_412),
.B(n_413),
.C(n_421),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_417),
.B2(n_418),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_444),
.C(n_445),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_419),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_420),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g421 ( 
.A(n_422),
.B(n_425),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_422),
.B(n_426),
.C(n_431),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_427),
.B1(n_430),
.B2(n_431),
.Y(n_425)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_426),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_427),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_436),
.B(n_451),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_436),
.B(n_451),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_437),
.B(n_442),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_441),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_441),
.C(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_439),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_442),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_443),
.B(n_446),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_443),
.B(n_447),
.C(n_449),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_449),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_463),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_454),
.B(n_463),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_455),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_460),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_457),
.B(n_460),
.C(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_469),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_467),
.B(n_469),
.Y(n_471)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_475),
.B(n_478),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_478),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx4f_ASAP7_75t_SL g481 ( 
.A(n_482),
.Y(n_481)
);

INVx13_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx8_ASAP7_75t_L g485 ( 
.A(n_483),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);


endmodule