module fake_jpeg_12349_n_634 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_634);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_634;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_SL g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_3),
.B(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_64),
.B(n_68),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_65),
.Y(n_189)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_26),
.A2(n_33),
.B1(n_29),
.B2(n_44),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_67),
.A2(n_127),
.B1(n_56),
.B2(n_29),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_17),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_69),
.B(n_82),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_70),
.Y(n_206)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_74),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_79),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_80),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_17),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_85),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_21),
.B(n_30),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_16),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_90),
.B(n_91),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_31),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_92),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_95),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_19),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_98),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_20),
.B(n_1),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_99),
.B(n_104),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_103),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_37),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_106),
.Y(n_160)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_110),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_111),
.Y(n_176)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_113),
.B(n_119),
.Y(n_212)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_22),
.Y(n_115)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_116),
.Y(n_211)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_22),
.Y(n_117)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_118),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_37),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_25),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_125),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_21),
.B(n_30),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_54),
.B(n_16),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_126),
.B(n_15),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_26),
.A2(n_33),
.B1(n_29),
.B2(n_23),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_32),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_134),
.B(n_144),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_68),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_135),
.B(n_154),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_99),
.B(n_54),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_32),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_153),
.B(n_155),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_84),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_42),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_74),
.B(n_42),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_161),
.B(n_164),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_66),
.B(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_169),
.B(n_174),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_45),
.Y(n_174)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_65),
.B(n_45),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_182),
.B(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_185),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_84),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_123),
.B1(n_120),
.B2(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_89),
.Y(n_192)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_192),
.Y(n_239)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_114),
.B(n_38),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_172),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_71),
.A2(n_26),
.B1(n_33),
.B2(n_29),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_198),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_97),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_76),
.Y(n_237)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_60),
.Y(n_202)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_202),
.Y(n_248)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_61),
.Y(n_203)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_203),
.Y(n_290)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_62),
.Y(n_204)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_204),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_83),
.A2(n_23),
.B1(n_46),
.B2(n_56),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_205),
.A2(n_108),
.B1(n_101),
.B2(n_105),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_217),
.A2(n_227),
.B1(n_163),
.B2(n_195),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_38),
.C(n_36),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_218),
.B(n_260),
.C(n_275),
.Y(n_295)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_220),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_221),
.A2(n_268),
.B1(n_151),
.B2(n_130),
.Y(n_348)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_213),
.A2(n_46),
.B1(n_23),
.B2(n_210),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_223),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_96),
.Y(n_224)
);

OAI21xp33_ASAP7_75t_L g334 ( 
.A1(n_224),
.A2(n_236),
.B(n_238),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_133),
.A2(n_98),
.B1(n_85),
.B2(n_80),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_228),
.Y(n_335)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_230),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_206),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_231),
.B(n_247),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_131),
.A2(n_46),
.B1(n_96),
.B2(n_34),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_232),
.Y(n_349)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_235),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_141),
.B(n_50),
.Y(n_236)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_SL g238 ( 
.A(n_188),
.B(n_49),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_142),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_241),
.Y(n_291)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_139),
.Y(n_242)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_242),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_159),
.B(n_49),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_244),
.B(n_269),
.Y(n_326)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_178),
.Y(n_245)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_141),
.B(n_159),
.Y(n_247)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_148),
.Y(n_250)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_250),
.Y(n_300)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_156),
.Y(n_251)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_251),
.Y(n_309)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_158),
.Y(n_252)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_129),
.Y(n_253)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_253),
.Y(n_340)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_166),
.Y(n_255)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_255),
.Y(n_319)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_160),
.Y(n_256)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_256),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_258),
.B(n_266),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_212),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_271),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_157),
.B(n_47),
.C(n_34),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_205),
.A2(n_75),
.B1(n_50),
.B2(n_55),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_261),
.A2(n_262),
.B1(n_270),
.B2(n_278),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_190),
.A2(n_55),
.B1(n_53),
.B2(n_47),
.Y(n_262)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_263),
.Y(n_346)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_145),
.Y(n_264)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_264),
.Y(n_307)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_145),
.Y(n_265)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_167),
.B(n_53),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_267),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_137),
.A2(n_36),
.B1(n_59),
.B2(n_4),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_183),
.B(n_15),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_152),
.A2(n_59),
.B1(n_15),
.B2(n_37),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g273 ( 
.A(n_215),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_273),
.B(n_285),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_138),
.Y(n_274)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_274),
.Y(n_344)
);

XNOR2x1_ASAP7_75t_L g275 ( 
.A(n_183),
.B(n_2),
.Y(n_275)
);

INVx11_ASAP7_75t_L g276 ( 
.A(n_211),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_129),
.Y(n_279)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_280),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_212),
.B(n_4),
.C(n_5),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_281),
.B(n_283),
.C(n_8),
.Y(n_316)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_194),
.Y(n_282)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_152),
.B(n_5),
.C(n_7),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_184),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_284),
.B(n_245),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_214),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_214),
.B(n_5),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_286),
.B(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_149),
.B(n_7),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_130),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_288),
.B(n_136),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_165),
.B(n_175),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_289),
.B(n_168),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_293),
.A2(n_151),
.B1(n_253),
.B2(n_228),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_276),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_297),
.B(n_314),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_261),
.A2(n_140),
.B1(n_147),
.B2(n_146),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_304),
.A2(n_342),
.B1(n_288),
.B2(n_279),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_217),
.A2(n_146),
.B1(n_179),
.B2(n_140),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g375 ( 
.A1(n_306),
.A2(n_304),
.B1(n_342),
.B2(n_298),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_246),
.B(n_170),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_308),
.B(n_318),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_221),
.A2(n_147),
.B1(n_195),
.B2(n_186),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_313),
.A2(n_327),
.B1(n_336),
.B2(n_339),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_266),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_316),
.B(n_320),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_171),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_272),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_226),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_225),
.Y(n_365)
);

NAND3xp33_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_325),
.C(n_10),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_216),
.B(n_162),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_258),
.A2(n_227),
.B1(n_219),
.B2(n_223),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_224),
.B(n_143),
.C(n_186),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_328),
.B(n_231),
.C(n_232),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_218),
.A2(n_136),
.B1(n_181),
.B2(n_150),
.Y(n_336)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_247),
.A2(n_208),
.B(n_143),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_233),
.B(n_132),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_341),
.B(n_347),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_262),
.A2(n_179),
.B1(n_181),
.B2(n_150),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_345),
.B(n_267),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_234),
.B(n_163),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_271),
.B1(n_230),
.B2(n_242),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g351 ( 
.A(n_339),
.B(n_236),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_SL g409 ( 
.A(n_351),
.B(n_393),
.C(n_330),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_376),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_281),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_301),
.B(n_277),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_354),
.B(n_355),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_315),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_356),
.B(n_369),
.C(n_395),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_290),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_294),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_366),
.Y(n_404)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_361),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_229),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_362),
.B(n_365),
.Y(n_405)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_295),
.B(n_249),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_367),
.A2(n_382),
.B1(n_349),
.B2(n_327),
.Y(n_402)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_368),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_295),
.B(n_275),
.C(n_239),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_307),
.Y(n_371)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_371),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_254),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_374),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_305),
.B(n_274),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g396 ( 
.A1(n_375),
.A2(n_384),
.B1(n_293),
.B2(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_377),
.Y(n_399)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_335),
.Y(n_378)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_378),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_317),
.B(n_240),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_386),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_345),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_381),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_298),
.A2(n_268),
.B1(n_264),
.B2(n_265),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_255),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_383),
.A2(n_344),
.B(n_329),
.Y(n_403)
);

INVx13_ASAP7_75t_L g385 ( 
.A(n_291),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_300),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_339),
.B(n_263),
.Y(n_387)
);

NOR2x1_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_394),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_300),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_344),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g389 ( 
.A1(n_312),
.A2(n_257),
.B1(n_271),
.B2(n_235),
.Y(n_389)
);

OAI22xp33_ASAP7_75t_SL g411 ( 
.A1(n_389),
.A2(n_390),
.B1(n_292),
.B2(n_343),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_299),
.B(n_284),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_391),
.Y(n_410)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_392),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_334),
.B(n_208),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_316),
.B(n_336),
.C(n_323),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_396),
.A2(n_402),
.B1(n_414),
.B2(n_417),
.Y(n_442)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_370),
.A2(n_349),
.B(n_312),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_418),
.Y(n_443)
);

NAND2xp33_ASAP7_75t_SL g462 ( 
.A(n_403),
.B(n_352),
.Y(n_462)
);

AO21x1_ASAP7_75t_L g455 ( 
.A1(n_409),
.A2(n_364),
.B(n_351),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_356),
.B1(n_383),
.B2(n_376),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_393),
.B(n_343),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_370),
.Y(n_457)
);

AND2x2_ASAP7_75t_SL g413 ( 
.A(n_360),
.B(n_296),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_432),
.B(n_380),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_382),
.A2(n_329),
.B1(n_296),
.B2(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_415),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_367),
.A2(n_340),
.B1(n_333),
.B2(n_319),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_350),
.B(n_319),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g419 ( 
.A(n_357),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_419),
.B(n_430),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_330),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_423),
.B(n_425),
.C(n_433),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_350),
.B(n_355),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_395),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_353),
.B(n_309),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_354),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_387),
.A2(n_303),
.B(n_302),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_309),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_435),
.Y(n_469)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_437),
.Y(n_474)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_426),
.Y(n_438)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

INVx4_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_439),
.A2(n_450),
.B1(n_454),
.B2(n_458),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_440),
.Y(n_472)
);

BUFx12f_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_441),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_449),
.Y(n_473)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_421),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_459),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_446),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_358),
.Y(n_448)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_448),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_358),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_426),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_451),
.A2(n_455),
.B1(n_457),
.B2(n_373),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_415),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_452),
.B(n_465),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_401),
.B(n_362),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_453),
.B(n_410),
.Y(n_480)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_397),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_407),
.B(n_359),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_456),
.Y(n_484)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_407),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_404),
.B(n_383),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_460),
.B(n_467),
.C(n_427),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_398),
.B(n_381),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_461),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_462),
.A2(n_468),
.B(n_432),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_398),
.B(n_363),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_463),
.Y(n_490)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_403),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_464),
.B(n_466),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_405),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_420),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_427),
.B(n_379),
.C(n_371),
.Y(n_467)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_397),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_470),
.B(n_479),
.C(n_488),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_476),
.B(n_466),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_440),
.A2(n_413),
.B(n_404),
.Y(n_478)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_478),
.A2(n_499),
.B(n_399),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_433),
.C(n_423),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_480),
.B(n_496),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_425),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_481),
.B(n_483),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_436),
.B(n_413),
.Y(n_483)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_486),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_454),
.A2(n_402),
.B1(n_414),
.B2(n_417),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_487),
.A2(n_491),
.B1(n_375),
.B2(n_378),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_408),
.Y(n_488)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_408),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_489),
.B(n_385),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_443),
.A2(n_390),
.B1(n_412),
.B2(n_409),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_492),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_459),
.B(n_373),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_464),
.B(n_461),
.C(n_455),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_501),
.C(n_388),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_443),
.A2(n_400),
.B(n_431),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_447),
.B(n_422),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_500),
.B(n_431),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_448),
.B(n_352),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_493),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_503),
.B(n_509),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_482),
.A2(n_458),
.B1(n_451),
.B2(n_434),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_504),
.A2(n_505),
.B1(n_506),
.B2(n_507),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_490),
.A2(n_434),
.B1(n_463),
.B2(n_449),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_490),
.A2(n_456),
.B1(n_457),
.B2(n_442),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_498),
.A2(n_450),
.B1(n_435),
.B2(n_400),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_446),
.Y(n_508)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_471),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_477),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_511),
.A2(n_524),
.B1(n_526),
.B2(n_527),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_497),
.B(n_441),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_512),
.B(n_515),
.Y(n_539)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_469),
.Y(n_513)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_469),
.Y(n_514)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_514),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_516),
.B(n_519),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_485),
.A2(n_375),
.B1(n_441),
.B2(n_439),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_517),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_361),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_518),
.B(n_529),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_473),
.B(n_441),
.Y(n_521)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_521),
.Y(n_546)
);

CKINVDCx14_ASAP7_75t_R g524 ( 
.A(n_473),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_474),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_SL g528 ( 
.A1(n_491),
.A2(n_399),
.B1(n_445),
.B2(n_420),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_528),
.A2(n_476),
.B(n_499),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_487),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_488),
.B(n_386),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_531),
.B(n_501),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_522),
.B(n_470),
.C(n_479),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_532),
.B(n_535),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_534),
.A2(n_494),
.B(n_514),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_483),
.C(n_472),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_536),
.B(n_555),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_525),
.B(n_472),
.C(n_489),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_541),
.B(n_548),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g548 ( 
.A1(n_503),
.A2(n_528),
.B(n_529),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_518),
.B(n_478),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_549),
.B(n_532),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_525),
.B(n_520),
.C(n_516),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_552),
.C(n_502),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_523),
.B(n_498),
.C(n_484),
.Y(n_552)
);

INVxp33_ASAP7_75t_SL g553 ( 
.A(n_508),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_553),
.A2(n_511),
.B1(n_494),
.B2(n_509),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_554),
.B(n_517),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_519),
.B(n_475),
.Y(n_555)
);

XOR2xp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_530),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_556),
.B(n_560),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_546),
.Y(n_557)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_557),
.Y(n_581)
);

FAx1_ASAP7_75t_SL g558 ( 
.A(n_535),
.B(n_484),
.CI(n_510),
.CON(n_558),
.SN(n_558)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_558),
.B(n_539),
.Y(n_576)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_533),
.Y(n_559)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_559),
.Y(n_585)
);

BUFx12_ASAP7_75t_L g561 ( 
.A(n_545),
.Y(n_561)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_561),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_562),
.B(n_563),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_550),
.B(n_551),
.C(n_541),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_SL g588 ( 
.A(n_564),
.B(n_385),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_547),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_565),
.B(n_567),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_542),
.B(n_502),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_566),
.B(n_574),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_SL g590 ( 
.A1(n_568),
.A2(n_377),
.B(n_368),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_540),
.A2(n_513),
.B1(n_527),
.B2(n_475),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_570),
.A2(n_544),
.B1(n_552),
.B2(n_542),
.Y(n_580)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_571),
.B(n_572),
.Y(n_586)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_543),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_540),
.A2(n_495),
.B1(n_375),
.B2(n_392),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_576),
.A2(n_587),
.B(n_569),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_SL g577 ( 
.A1(n_558),
.A2(n_544),
.B(n_537),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_577),
.A2(n_566),
.B1(n_568),
.B2(n_556),
.Y(n_597)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_580),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_575),
.B(n_554),
.C(n_555),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_584),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_560),
.B(n_495),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g587 ( 
.A1(n_573),
.A2(n_292),
.B(n_346),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_588),
.B(n_592),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_SL g598 ( 
.A1(n_590),
.A2(n_567),
.B(n_561),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_SL g592 ( 
.A(n_564),
.B(n_377),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_569),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_598),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_578),
.B(n_557),
.Y(n_596)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_596),
.Y(n_614)
);

XOR2x1_ASAP7_75t_SL g610 ( 
.A(n_597),
.B(n_588),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_585),
.B(n_565),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_599),
.B(n_600),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_583),
.B(n_563),
.C(n_574),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_601),
.B(n_602),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_586),
.B(n_561),
.Y(n_602)
);

OAI22xp5_ASAP7_75t_SL g603 ( 
.A1(n_591),
.A2(n_303),
.B1(n_302),
.B2(n_337),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_603),
.A2(n_590),
.B1(n_592),
.B2(n_273),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_582),
.B(n_310),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g608 ( 
.A(n_604),
.B(n_581),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_579),
.B(n_337),
.C(n_346),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g616 ( 
.A(n_605),
.B(n_332),
.C(n_310),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_613),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_610),
.B(n_615),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_612),
.B(n_616),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_595),
.B(n_577),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_601),
.B(n_579),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_614),
.A2(n_593),
.B1(n_594),
.B2(n_605),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_618),
.B(n_619),
.Y(n_625)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_609),
.A2(n_598),
.B(n_597),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_607),
.A2(n_611),
.B(n_615),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_621),
.B(n_610),
.C(n_606),
.Y(n_624)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_611),
.Y(n_622)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_622),
.A2(n_606),
.B(n_332),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_SL g628 ( 
.A1(n_624),
.A2(n_626),
.B(n_627),
.Y(n_628)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_620),
.B(n_248),
.C(n_368),
.Y(n_627)
);

AOI322xp5_ASAP7_75t_L g629 ( 
.A1(n_625),
.A2(n_623),
.A3(n_617),
.B1(n_273),
.B2(n_220),
.C1(n_222),
.C2(n_13),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_10),
.C(n_11),
.Y(n_630)
);

MAJx2_ASAP7_75t_L g631 ( 
.A(n_630),
.B(n_628),
.C(n_12),
.Y(n_631)
);

XOR2xp5_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_11),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_632),
.A2(n_13),
.B1(n_14),
.B2(n_220),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_633),
.B(n_13),
.Y(n_634)
);


endmodule