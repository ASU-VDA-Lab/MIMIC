module fake_ariane_1744_n_1773 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1773);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1773;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_26),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_72),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_134),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_33),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_101),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_58),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_86),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_68),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_13),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_115),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_64),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_71),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_121),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_3),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_11),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_28),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_1),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_54),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_67),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_89),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_14),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_30),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_57),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_153),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_107),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_6),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_141),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_27),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_23),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_109),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_23),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_88),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_45),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_65),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_136),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_92),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_16),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_123),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_112),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_22),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_146),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_80),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_26),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_44),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_3),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_73),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_162),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_104),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_34),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_122),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_110),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_124),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_44),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_17),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_74),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_50),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_6),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_75),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_33),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_127),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_32),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_52),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_129),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_93),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_42),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_120),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_135),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_21),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_119),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_51),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_105),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_13),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_142),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_11),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_103),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_55),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g260 ( 
.A(n_21),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_138),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_56),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_132),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_79),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_91),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_18),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_14),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_12),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_38),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_133),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_95),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_1),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_39),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_149),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_49),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_22),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_30),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_83),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_4),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_61),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_98),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_5),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_19),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_57),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_43),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_108),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_46),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_156),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_53),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_53),
.Y(n_296)
);

INVx4_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_139),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_85),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_145),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_155),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_78),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_41),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_147),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_47),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_19),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_116),
.Y(n_308)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_58),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_161),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_38),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_25),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_160),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_35),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_42),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_7),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_49),
.Y(n_317)
);

INVxp33_ASAP7_75t_SL g318 ( 
.A(n_25),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_62),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_15),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_29),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_10),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_51),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_20),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_223),
.Y(n_326)
);

NOR2xp67_ASAP7_75t_L g327 ( 
.A(n_280),
.B(n_2),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_223),
.Y(n_328)
);

CKINVDCx14_ASAP7_75t_R g329 ( 
.A(n_253),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_239),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_239),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_223),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_223),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_218),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_221),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_223),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_223),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_236),
.Y(n_338)
);

INVxp33_ASAP7_75t_SL g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_223),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_237),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_302),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_318),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_164),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_167),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_L g346 ( 
.A(n_280),
.B(n_219),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_169),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_223),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_171),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_174),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_223),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_271),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_227),
.B(n_2),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_260),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_190),
.Y(n_356)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_199),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_215),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_227),
.B(n_4),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_168),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_168),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_181),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_182),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_176),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_178),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_183),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_178),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_187),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_224),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_275),
.Y(n_371)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_184),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_187),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_189),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_283),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_198),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_189),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_252),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_180),
.Y(n_379)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_180),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_199),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_195),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_200),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_203),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_209),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_195),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_252),
.B(n_7),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_197),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_271),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_191),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_197),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_199),
.Y(n_392)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_202),
.B(n_8),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_208),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_202),
.B(n_9),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_210),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_217),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_212),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_205),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_217),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_205),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_211),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_309),
.B(n_211),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_271),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_326),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_360),
.B(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_385),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_333),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_328),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_336),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_333),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_361),
.B(n_244),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_403),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_357),
.B(n_225),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_337),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_340),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_364),
.B(n_244),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_387),
.B(n_207),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_340),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_348),
.Y(n_431)
);

AND3x2_ASAP7_75t_L g432 ( 
.A(n_355),
.B(n_300),
.C(n_288),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_357),
.B(n_220),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_357),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_263),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_352),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_365),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_365),
.B(n_263),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_366),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_366),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_368),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_330),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_368),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_369),
.B(n_288),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_373),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_374),
.B(n_303),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_374),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_331),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_334),
.Y(n_457)
);

AND3x2_ASAP7_75t_L g458 ( 
.A(n_354),
.B(n_304),
.C(n_303),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_377),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_359),
.B(n_327),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_377),
.B(n_304),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_344),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

OA21x2_ASAP7_75t_L g465 ( 
.A1(n_386),
.A2(n_226),
.B(n_220),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_388),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_391),
.B(n_317),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

AND2x4_ASAP7_75t_L g472 ( 
.A(n_399),
.B(n_317),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_353),
.B(n_226),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_401),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_217),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_402),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_345),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_423),
.B(n_389),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_423),
.B(n_329),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_459),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_426),
.Y(n_481)
);

INVxp33_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_460),
.A2(n_339),
.B1(n_378),
.B2(n_327),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_459),
.B(n_462),
.Y(n_484)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_473),
.B(n_350),
.C(n_347),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_402),
.Y(n_486)
);

HB1xp67_ASAP7_75t_SL g487 ( 
.A(n_463),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_429),
.B(n_372),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_406),
.B(n_379),
.Y(n_489)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_456),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

BUFx8_ASAP7_75t_SL g492 ( 
.A(n_463),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_459),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_459),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_426),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_444),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_459),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_406),
.B(n_380),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_429),
.B(n_460),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_463),
.Y(n_501)
);

BUFx6f_ASAP7_75t_SL g502 ( 
.A(n_475),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_R g504 ( 
.A(n_457),
.B(n_335),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_424),
.B(n_351),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_457),
.B(n_338),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_424),
.B(n_362),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_454),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_439),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g513 ( 
.A(n_477),
.B(n_393),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_449),
.B(n_363),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_449),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_426),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_431),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_441),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_R g519 ( 
.A(n_432),
.B(n_356),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_434),
.Y(n_520)
);

BUFx10_ASAP7_75t_L g521 ( 
.A(n_477),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_431),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_441),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_451),
.B(n_367),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_465),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_434),
.B(n_376),
.Y(n_527)
);

AO22x1_ASAP7_75t_L g528 ( 
.A1(n_473),
.A2(n_343),
.B1(n_398),
.B2(n_396),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_440),
.B(n_393),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

AND2x6_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_246),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_431),
.Y(n_532)
);

INVxp33_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_465),
.A2(n_400),
.B1(n_397),
.B2(n_392),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_441),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_440),
.B(n_395),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_451),
.B(n_383),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_459),
.B(n_384),
.Y(n_538)
);

INVx5_ASAP7_75t_L g539 ( 
.A(n_459),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_442),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_462),
.Y(n_541)
);

INVx2_ASAP7_75t_SL g542 ( 
.A(n_406),
.Y(n_542)
);

INVx8_ASAP7_75t_L g543 ( 
.A(n_475),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_442),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_442),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_434),
.B(n_394),
.Y(n_547)
);

INVx4_ASAP7_75t_L g548 ( 
.A(n_451),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_462),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_455),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_451),
.B(n_390),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_434),
.B(n_341),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_443),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_443),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_453),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

AND2x2_ASAP7_75t_SL g558 ( 
.A(n_465),
.B(n_194),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_451),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_462),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_455),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_462),
.B(n_468),
.Y(n_565)
);

BUFx3_ASAP7_75t_L g566 ( 
.A(n_420),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_476),
.B(n_346),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_476),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_462),
.B(n_468),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_445),
.B(n_342),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_346),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_475),
.A2(n_251),
.B1(n_325),
.B2(n_323),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_462),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_438),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_476),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_448),
.B(n_395),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_440),
.B(n_422),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_462),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_421),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_422),
.B(n_191),
.Y(n_580)
);

BUFx6f_ASAP7_75t_SL g581 ( 
.A(n_475),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_258),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_450),
.B(n_466),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_421),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_465),
.Y(n_586)
);

HAxp5_ASAP7_75t_SL g587 ( 
.A(n_432),
.B(n_358),
.CON(n_587),
.SN(n_587)
);

INVx8_ASAP7_75t_L g588 ( 
.A(n_475),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_450),
.B(n_246),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_468),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

OR2x6_ASAP7_75t_L g592 ( 
.A(n_422),
.B(n_193),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_404),
.B(n_254),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_468),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_421),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_466),
.B(n_254),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_469),
.B(n_264),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_421),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_469),
.B(n_258),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_474),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_471),
.B(n_264),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_412),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_468),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_412),
.Y(n_604)
);

AND3x2_ASAP7_75t_L g605 ( 
.A(n_404),
.B(n_196),
.C(n_193),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_404),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_412),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_474),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_446),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_446),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_446),
.Y(n_611)
);

OR2x6_ASAP7_75t_L g612 ( 
.A(n_422),
.B(n_196),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_405),
.B(n_273),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_412),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_422),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_405),
.B(n_273),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_446),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_407),
.B(n_409),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_468),
.B(n_292),
.Y(n_619)
);

NOR2x1p5_ASAP7_75t_L g620 ( 
.A(n_404),
.B(n_234),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_L g621 ( 
.A1(n_465),
.A2(n_312),
.B1(n_248),
.B2(n_245),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_407),
.B(n_292),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_435),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_412),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_435),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_464),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_409),
.B(n_305),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_464),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_505),
.B(n_435),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_509),
.B(n_435),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_579),
.Y(n_631)
);

A2O1A1Ixp33_ASAP7_75t_L g632 ( 
.A1(n_500),
.A2(n_464),
.B(n_467),
.C(n_470),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_490),
.B(n_435),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_504),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_478),
.B(n_437),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_L g636 ( 
.A1(n_558),
.A2(n_465),
.B1(n_470),
.B2(n_447),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_488),
.B(n_437),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_564),
.B(n_404),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_420),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_606),
.B(n_437),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_527),
.B(n_437),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_606),
.B(n_437),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_521),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_586),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_547),
.B(n_404),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_570),
.A2(n_593),
.B1(n_531),
.B2(n_581),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_486),
.B(n_433),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_566),
.Y(n_648)
);

BUFx8_ASAP7_75t_L g649 ( 
.A(n_564),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_521),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_542),
.B(n_433),
.Y(n_651)
);

NOR2xp67_ASAP7_75t_L g652 ( 
.A(n_485),
.B(n_479),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_542),
.B(n_414),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_579),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_551),
.B(n_414),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_585),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_585),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_583),
.B(n_416),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_503),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_521),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_520),
.Y(n_661)
);

NAND2x1_ASAP7_75t_L g662 ( 
.A(n_623),
.B(n_464),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_558),
.A2(n_621),
.B1(n_526),
.B2(n_593),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_508),
.Y(n_664)
);

OR2x2_ASAP7_75t_L g665 ( 
.A(n_497),
.B(n_422),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_600),
.B(n_416),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_595),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_552),
.B(n_418),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_514),
.B(n_418),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_595),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_499),
.B(n_608),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_499),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_512),
.Y(n_673)
);

INVx8_ASAP7_75t_L g674 ( 
.A(n_543),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_598),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_550),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_526),
.B(n_420),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_580),
.A2(n_612),
.B1(n_592),
.B2(n_482),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_598),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_525),
.B(n_419),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_526),
.B(n_623),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_481),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_481),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_524),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_593),
.A2(n_472),
.B1(n_470),
.B2(n_428),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_543),
.Y(n_687)
);

INVx2_ASAP7_75t_SL g688 ( 
.A(n_550),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_535),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_540),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_537),
.B(n_615),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_577),
.B(n_428),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_571),
.B(n_419),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_623),
.B(n_425),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_593),
.A2(n_472),
.B1(n_470),
.B2(n_428),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_544),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_580),
.A2(n_467),
.B1(n_234),
.B2(n_235),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_510),
.B(n_428),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_489),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_496),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_545),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_625),
.B(n_425),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_513),
.B(n_427),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_496),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_511),
.Y(n_705)
);

INVxp67_ASAP7_75t_L g706 ( 
.A(n_487),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_593),
.A2(n_472),
.B1(n_470),
.B2(n_428),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_546),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_553),
.Y(n_709)
);

AND2x4_ASAP7_75t_SL g710 ( 
.A(n_513),
.B(n_370),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_593),
.A2(n_472),
.B1(n_470),
.B2(n_428),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_520),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_489),
.B(n_427),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_554),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_482),
.B(n_533),
.Y(n_715)
);

NAND2x1p5_ASAP7_75t_L g716 ( 
.A(n_577),
.B(n_436),
.Y(n_716)
);

INVxp67_ASAP7_75t_L g717 ( 
.A(n_507),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_489),
.B(n_430),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_620),
.B(n_458),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_586),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_576),
.B(n_430),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_467),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_543),
.Y(n_723)
);

AOI221xp5_ASAP7_75t_L g724 ( 
.A1(n_483),
.A2(n_248),
.B1(n_261),
.B2(n_268),
.C(n_269),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_511),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_516),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_528),
.B(n_467),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_516),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_555),
.B(n_436),
.Y(n_729)
);

NOR2x1p5_ASAP7_75t_L g730 ( 
.A(n_492),
.B(n_216),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_559),
.B(n_472),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_625),
.B(n_436),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_R g733 ( 
.A(n_501),
.B(n_371),
.Y(n_733)
);

INVxp33_ASAP7_75t_SL g734 ( 
.A(n_572),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_517),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_560),
.B(n_436),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_568),
.B(n_436),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_575),
.B(n_436),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_582),
.B(n_472),
.Y(n_739)
);

OR2x2_ASAP7_75t_SL g740 ( 
.A(n_587),
.B(n_375),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_531),
.A2(n_461),
.B1(n_452),
.B2(n_447),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_543),
.A2(n_270),
.B1(n_287),
.B2(n_259),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_513),
.B(n_458),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_609),
.Y(n_744)
);

AO221x1_ASAP7_75t_L g745 ( 
.A1(n_587),
.A2(n_312),
.B1(n_296),
.B2(n_235),
.C(n_241),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_517),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_594),
.B(n_447),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_588),
.A2(n_618),
.B1(n_580),
.B2(n_612),
.Y(n_748)
);

NOR3xp33_ASAP7_75t_L g749 ( 
.A(n_538),
.B(n_245),
.C(n_241),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_594),
.B(n_603),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_492),
.B(n_207),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_599),
.B(n_461),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_627),
.B(n_461),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_513),
.B(n_447),
.Y(n_754)
);

HB1xp67_ASAP7_75t_L g755 ( 
.A(n_501),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_523),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_531),
.B(n_461),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_531),
.B(n_461),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_529),
.B(n_447),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_588),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_531),
.B(n_461),
.Y(n_761)
);

NAND3xp33_ASAP7_75t_L g762 ( 
.A(n_533),
.B(n_229),
.C(n_222),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_610),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_531),
.B(n_447),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_534),
.A2(n_269),
.B1(n_289),
.B2(n_279),
.C(n_296),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_602),
.B(n_452),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_502),
.A2(n_452),
.B1(n_314),
.B2(n_307),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_602),
.B(n_452),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_594),
.B(n_603),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_523),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_530),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_611),
.Y(n_772)
);

XNOR2xp5_ASAP7_75t_L g773 ( 
.A(n_605),
.B(n_452),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_529),
.B(n_452),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_305),
.Y(n_775)
);

O2A1O1Ixp5_ASAP7_75t_L g776 ( 
.A1(n_538),
.A2(n_417),
.B(n_415),
.C(n_411),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_617),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_589),
.B(n_279),
.C(n_268),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_626),
.A2(n_289),
.B(n_306),
.C(n_307),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_529),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_604),
.B(n_306),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_530),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_628),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_607),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_594),
.B(n_194),
.Y(n_785)
);

INVx4_ASAP7_75t_L g786 ( 
.A(n_588),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_607),
.B(n_314),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_603),
.B(n_232),
.Y(n_788)
);

OAI221xp5_ASAP7_75t_L g789 ( 
.A1(n_536),
.A2(n_257),
.B1(n_238),
.B2(n_322),
.C(n_321),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_536),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_502),
.A2(n_207),
.B1(n_230),
.B2(n_308),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_532),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_532),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_556),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_614),
.B(n_624),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_614),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_536),
.B(n_588),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_624),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_659),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_734),
.B(n_536),
.Y(n_800)
);

CKINVDCx6p67_ASAP7_75t_R g801 ( 
.A(n_755),
.Y(n_801)
);

O2A1O1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_637),
.A2(n_622),
.B(n_613),
.C(n_616),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_641),
.A2(n_495),
.B(n_491),
.Y(n_803)
);

AND2x2_ASAP7_75t_L g804 ( 
.A(n_676),
.B(n_580),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_631),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_699),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_672),
.B(n_592),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_637),
.B(n_592),
.Y(n_808)
);

AND2x2_ASAP7_75t_SL g809 ( 
.A(n_663),
.B(n_232),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_713),
.B(n_592),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_671),
.A2(n_596),
.B(n_601),
.C(n_597),
.Y(n_811)
);

INVxp67_ASAP7_75t_SL g812 ( 
.A(n_687),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_668),
.A2(n_548),
.B1(n_491),
.B2(n_495),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_691),
.A2(n_556),
.B(n_557),
.C(n_563),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_677),
.A2(n_495),
.B(n_491),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_678),
.B(n_612),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_677),
.A2(n_522),
.B(n_515),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_649),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_664),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_631),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_681),
.A2(n_522),
.B(n_515),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_776),
.A2(n_565),
.B(n_484),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_654),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_674),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_718),
.B(n_612),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_691),
.B(n_515),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_669),
.A2(n_563),
.B(n_574),
.C(n_557),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_688),
.B(n_574),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_649),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_681),
.A2(n_548),
.B(n_522),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_797),
.A2(n_581),
.B1(n_502),
.B2(n_484),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_629),
.A2(n_630),
.B(n_644),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_760),
.Y(n_834)
);

OAI21xp5_ASAP7_75t_L g835 ( 
.A1(n_669),
.A2(n_569),
.B(n_565),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_663),
.B(n_791),
.Y(n_836)
);

BUFx4f_ASAP7_75t_L g837 ( 
.A(n_674),
.Y(n_837)
);

OAI21xp5_ASAP7_75t_L g838 ( 
.A1(n_680),
.A2(n_642),
.B(n_640),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_647),
.B(n_548),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_760),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_654),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_720),
.A2(n_569),
.B(n_561),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_760),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_651),
.A2(n_619),
.B(n_561),
.C(n_498),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_750),
.A2(n_498),
.B(n_480),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_680),
.A2(n_642),
.B(n_640),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_635),
.B(n_480),
.Y(n_847)
);

AND2x2_ASAP7_75t_SL g848 ( 
.A(n_791),
.B(n_265),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_750),
.A2(n_619),
.B(n_410),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_715),
.B(n_243),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_769),
.A2(n_498),
.B(n_480),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_635),
.B(n_562),
.Y(n_852)
);

INVx2_ASAP7_75t_SL g853 ( 
.A(n_733),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_692),
.B(n_562),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_769),
.A2(n_573),
.B(n_562),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_692),
.B(n_573),
.Y(n_856)
);

INVx4_ASAP7_75t_L g857 ( 
.A(n_674),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_692),
.B(n_573),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_760),
.B(n_603),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_780),
.B(n_581),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_703),
.B(n_578),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_703),
.B(n_578),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_694),
.A2(n_584),
.B(n_578),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_658),
.B(n_584),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_645),
.A2(n_584),
.B(n_603),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_634),
.B(n_255),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_666),
.B(n_493),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_795),
.A2(n_591),
.B(n_493),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_753),
.B(n_493),
.Y(n_869)
);

OAI22xp5_ASAP7_75t_L g870 ( 
.A1(n_786),
.A2(n_646),
.B1(n_653),
.B2(n_636),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_656),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_759),
.B(n_494),
.Y(n_872)
);

OAI21xp33_ASAP7_75t_L g873 ( 
.A1(n_739),
.A2(n_295),
.B(n_267),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_673),
.Y(n_874)
);

NAND2x1p5_ASAP7_75t_L g875 ( 
.A(n_786),
.B(n_723),
.Y(n_875)
);

CKINVDCx10_ASAP7_75t_R g876 ( 
.A(n_733),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_684),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_685),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_732),
.A2(n_265),
.B(n_308),
.C(n_417),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_723),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_655),
.A2(n_591),
.B(n_494),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_759),
.B(n_494),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_748),
.B(n_652),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_716),
.Y(n_884)
);

OAI21xp5_ASAP7_75t_L g885 ( 
.A1(n_694),
.A2(n_632),
.B(n_702),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_689),
.B(n_494),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_797),
.B(n_506),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_732),
.A2(n_308),
.B(n_415),
.C(n_411),
.Y(n_888)
);

AO21x1_ASAP7_75t_L g889 ( 
.A1(n_727),
.A2(n_410),
.B(n_411),
.Y(n_889)
);

BUFx4f_ASAP7_75t_L g890 ( 
.A(n_643),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_702),
.A2(n_417),
.B(n_410),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_638),
.B(n_506),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_633),
.A2(n_591),
.B(n_506),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_656),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_721),
.A2(n_693),
.B(n_662),
.Y(n_895)
);

OAI21xp5_ASAP7_75t_L g896 ( 
.A1(n_632),
.A2(n_539),
.B(n_590),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_657),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_690),
.B(n_506),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_650),
.B(n_549),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_706),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_717),
.B(n_274),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_661),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_724),
.A2(n_591),
.B(n_549),
.C(n_277),
.Y(n_903)
);

OAI321xp33_ASAP7_75t_L g904 ( 
.A1(n_697),
.A2(n_228),
.A3(n_209),
.B1(n_417),
.B2(n_408),
.C(n_415),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_636),
.A2(n_549),
.B1(n_315),
.B2(n_311),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_665),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_696),
.A2(n_549),
.B(n_278),
.C(n_281),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_752),
.A2(n_731),
.B(n_736),
.C(n_729),
.Y(n_908)
);

INVx2_ASAP7_75t_SL g909 ( 
.A(n_710),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_766),
.A2(n_768),
.B(n_747),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_701),
.A2(n_290),
.B(n_293),
.C(n_316),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_745),
.A2(n_207),
.B1(n_230),
.B2(n_320),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_737),
.A2(n_408),
.B(n_410),
.C(n_411),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_722),
.A2(n_590),
.B(n_541),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_740),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_784),
.A2(n_590),
.B(n_541),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_747),
.A2(n_590),
.B(n_541),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_796),
.A2(n_590),
.B(n_541),
.Y(n_918)
);

NAND2x1p5_ASAP7_75t_L g919 ( 
.A(n_661),
.B(n_539),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_708),
.B(n_539),
.Y(n_920)
);

OAI22xp5_ASAP7_75t_L g921 ( 
.A1(n_648),
.A2(n_541),
.B1(n_539),
.B2(n_165),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_712),
.Y(n_922)
);

INVx1_ASAP7_75t_SL g923 ( 
.A(n_710),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_709),
.B(n_539),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_754),
.B(n_9),
.Y(n_925)
);

O2A1O1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_738),
.A2(n_408),
.B(n_415),
.C(n_16),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_798),
.A2(n_408),
.B(n_242),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_714),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_682),
.A2(n_240),
.B(n_247),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_754),
.B(n_166),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_682),
.A2(n_231),
.B(n_233),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_686),
.B(n_413),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_765),
.B(n_170),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_683),
.A2(n_262),
.B(n_177),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_698),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_774),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_767),
.B(n_172),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_767),
.B(n_173),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_657),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_695),
.B(n_175),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_789),
.A2(n_763),
.B(n_744),
.C(n_772),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_660),
.B(n_519),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_707),
.B(n_179),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_790),
.B(n_10),
.Y(n_944)
);

OAI21xp5_ASAP7_75t_L g945 ( 
.A1(n_683),
.A2(n_276),
.B(n_188),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_712),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_700),
.A2(n_214),
.B(n_185),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_700),
.A2(n_213),
.B(n_186),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_757),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_777),
.A2(n_15),
.B(n_18),
.C(n_20),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_719),
.B(n_751),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_719),
.B(n_24),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_711),
.B(n_192),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_741),
.A2(n_228),
.A3(n_209),
.B1(n_519),
.B2(n_230),
.C(n_413),
.Y(n_954)
);

BUFx2_ASAP7_75t_L g955 ( 
.A(n_773),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_743),
.A2(n_284),
.B1(n_324),
.B2(n_319),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_704),
.A2(n_282),
.B(n_313),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_758),
.B(n_201),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_704),
.A2(n_272),
.B(n_310),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_749),
.B(n_204),
.Y(n_960)
);

BUFx4f_ASAP7_75t_L g961 ( 
.A(n_783),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_705),
.A2(n_285),
.B(n_301),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_778),
.B(n_206),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_705),
.A2(n_794),
.B(n_793),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_761),
.A2(n_266),
.B(n_299),
.C(n_298),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_743),
.B(n_764),
.Y(n_967)
);

AO21x2_ASAP7_75t_L g968 ( 
.A1(n_785),
.A2(n_297),
.B(n_230),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_762),
.B(n_24),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_725),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_725),
.B(n_249),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_794),
.B(n_250),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_726),
.B(n_413),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_726),
.A2(n_286),
.B(n_256),
.Y(n_974)
);

CKINVDCx6p67_ASAP7_75t_R g975 ( 
.A(n_787),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_728),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_735),
.A2(n_294),
.B(n_413),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_730),
.B(n_228),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_735),
.A2(n_413),
.B(n_228),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_793),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_742),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_667),
.Y(n_982)
);

AOI22xp5_ASAP7_75t_L g983 ( 
.A1(n_746),
.A2(n_228),
.B1(n_209),
.B2(n_413),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_746),
.A2(n_228),
.B(n_209),
.C(n_413),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_756),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_756),
.B(n_413),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_770),
.B(n_792),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_770),
.A2(n_297),
.B(n_209),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_836),
.A2(n_792),
.B1(n_771),
.B2(n_782),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_827),
.A2(n_639),
.B(n_771),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_827),
.A2(n_782),
.B(n_670),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_839),
.A2(n_679),
.B(n_670),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_833),
.A2(n_679),
.B(n_675),
.Y(n_993)
);

NOR3xp33_ASAP7_75t_SL g994 ( 
.A(n_911),
.B(n_779),
.C(n_775),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_813),
.A2(n_675),
.B(n_667),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_825),
.Y(n_996)
);

OR2x6_ASAP7_75t_SL g997 ( 
.A(n_876),
.B(n_779),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_816),
.A2(n_788),
.B1(n_785),
.B2(n_32),
.Y(n_998)
);

OAI21xp33_ASAP7_75t_L g999 ( 
.A1(n_925),
.A2(n_788),
.B(n_31),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_838),
.A2(n_29),
.B(n_35),
.C(n_36),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_803),
.A2(n_82),
.B(n_154),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_799),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_846),
.A2(n_36),
.B(n_37),
.C(n_39),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_967),
.B(n_37),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_819),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_808),
.A2(n_40),
.B(n_41),
.C(n_43),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_825),
.B(n_40),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_817),
.B(n_45),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_816),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_800),
.B(n_50),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_837),
.B(n_52),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_867),
.A2(n_106),
.B(n_150),
.Y(n_1012)
);

OR2x2_ASAP7_75t_L g1013 ( 
.A(n_906),
.B(n_54),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_800),
.B(n_55),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_837),
.B(n_961),
.Y(n_1015)
);

OR2x6_ASAP7_75t_L g1016 ( 
.A(n_909),
.B(n_853),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_883),
.A2(n_59),
.B(n_60),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_925),
.A2(n_63),
.B(n_69),
.C(n_77),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_836),
.A2(n_81),
.B1(n_90),
.B2(n_94),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_847),
.A2(n_852),
.B(n_869),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_805),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_R g1022 ( 
.A(n_830),
.B(n_96),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_900),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_906),
.B(n_99),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_883),
.A2(n_100),
.B(n_113),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_935),
.B(n_114),
.Y(n_1026)
);

CKINVDCx20_ASAP7_75t_R g1027 ( 
.A(n_801),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_935),
.B(n_117),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_961),
.B(n_126),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_951),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_807),
.B(n_128),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_850),
.B(n_131),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_864),
.A2(n_137),
.B(n_140),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_821),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_820),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_981),
.A2(n_807),
.B1(n_848),
.B2(n_804),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_834),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_969),
.A2(n_143),
.B(n_148),
.C(n_163),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_923),
.Y(n_1039)
);

OAI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_809),
.A2(n_848),
.B1(n_826),
.B2(n_810),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_890),
.B(n_857),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_949),
.B(n_936),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_895),
.A2(n_908),
.B(n_831),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_936),
.B(n_817),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_857),
.Y(n_1045)
);

NOR3xp33_ASAP7_75t_L g1046 ( 
.A(n_969),
.B(n_866),
.C(n_950),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_809),
.A2(n_878),
.B1(n_877),
.B2(n_874),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_941),
.A2(n_907),
.B(n_811),
.C(n_873),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_824),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_822),
.A2(n_802),
.B(n_865),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_815),
.A2(n_818),
.B(n_914),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_978),
.B(n_884),
.Y(n_1052)
);

O2A1O1Ixp5_ASAP7_75t_L g1053 ( 
.A1(n_859),
.A2(n_958),
.B(n_889),
.C(n_885),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_884),
.B(n_812),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_964),
.A2(n_858),
.B(n_854),
.C(n_856),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_834),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_SL g1057 ( 
.A1(n_859),
.A2(n_966),
.B(n_924),
.C(n_920),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_SL g1058 ( 
.A1(n_915),
.A2(n_955),
.B1(n_942),
.B2(n_952),
.Y(n_1058)
);

A2O1A1Ixp33_ASAP7_75t_L g1059 ( 
.A1(n_835),
.A2(n_903),
.B(n_944),
.C(n_962),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_928),
.A2(n_870),
.B1(n_812),
.B2(n_892),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_949),
.B(n_910),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_868),
.A2(n_881),
.B(n_893),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_944),
.A2(n_892),
.B(n_844),
.C(n_862),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_806),
.B(n_952),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_890),
.B(n_834),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_976),
.B(n_985),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_863),
.A2(n_855),
.B(n_851),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_872),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_814),
.A2(n_828),
.B(n_861),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_829),
.B(n_975),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_901),
.B(n_930),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_845),
.A2(n_842),
.B(n_823),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_886),
.A2(n_898),
.B1(n_882),
.B2(n_912),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_896),
.A2(n_916),
.B(n_918),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_912),
.B(n_948),
.C(n_945),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_841),
.B(n_894),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_973),
.A2(n_986),
.B(n_988),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_978),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_956),
.B(n_860),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_871),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_973),
.A2(n_986),
.B(n_917),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_840),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_937),
.A2(n_938),
.B1(n_933),
.B2(n_905),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_860),
.B(n_902),
.Y(n_1084)
);

NOR2x1p5_ASAP7_75t_L g1085 ( 
.A(n_843),
.B(n_960),
.Y(n_1085)
);

O2A1O1Ixp5_ASAP7_75t_L g1086 ( 
.A1(n_899),
.A2(n_957),
.B(n_927),
.C(n_932),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_926),
.A2(n_932),
.B(n_953),
.C(n_940),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_943),
.A2(n_913),
.B(n_902),
.C(n_978),
.Y(n_1088)
);

HB1xp67_ASAP7_75t_L g1089 ( 
.A(n_970),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_965),
.A2(n_987),
.B(n_904),
.Y(n_1090)
);

INVxp67_ASAP7_75t_L g1091 ( 
.A(n_971),
.Y(n_1091)
);

OR2x6_ASAP7_75t_L g1092 ( 
.A(n_875),
.B(n_887),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_875),
.A2(n_922),
.B1(n_946),
.B2(n_832),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_880),
.B(n_954),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_897),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_987),
.A2(n_921),
.B(n_946),
.Y(n_1096)
);

BUFx12f_ASAP7_75t_L g1097 ( 
.A(n_880),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_922),
.A2(n_843),
.B1(n_919),
.B2(n_972),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_970),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_939),
.B(n_982),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_977),
.A2(n_959),
.B(n_974),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_970),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_929),
.A2(n_947),
.B(n_934),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_980),
.B(n_931),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_980),
.B(n_919),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_963),
.B(n_879),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_888),
.B(n_983),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_849),
.B(n_979),
.Y(n_1108)
);

INVx6_ASAP7_75t_L g1109 ( 
.A(n_891),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_984),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_968),
.A2(n_827),
.B(n_839),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_838),
.B(n_846),
.Y(n_1112)
);

INVx3_ASAP7_75t_L g1113 ( 
.A(n_857),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_800),
.B(n_734),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_883),
.A2(n_870),
.B(n_846),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_876),
.B(n_634),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_816),
.A2(n_800),
.B1(n_743),
.B2(n_688),
.Y(n_1117)
);

OR2x2_ASAP7_75t_L g1118 ( 
.A(n_906),
.B(n_564),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_827),
.A2(n_839),
.B(n_641),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_805),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_838),
.A2(n_846),
.B(n_925),
.C(n_637),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_838),
.A2(n_423),
.B(n_488),
.C(n_505),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_853),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_800),
.B(n_564),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_891),
.A2(n_849),
.B(n_965),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_853),
.Y(n_1126)
);

OAI21x1_ASAP7_75t_L g1127 ( 
.A1(n_891),
.A2(n_849),
.B(n_965),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_817),
.B(n_884),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_808),
.A2(n_836),
.B1(n_925),
.B2(n_809),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_816),
.A2(n_734),
.B1(n_501),
.B2(n_688),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_800),
.B(n_734),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_827),
.A2(n_839),
.B(n_641),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_R g1133 ( 
.A(n_876),
.B(n_634),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_838),
.B(n_846),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_825),
.B(n_676),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_800),
.B(n_505),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_827),
.A2(n_839),
.B(n_641),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1129),
.A2(n_1046),
.B1(n_1114),
.B2(n_1131),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1136),
.B(n_1130),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1071),
.C(n_1075),
.Y(n_1140)
);

OAI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1129),
.A2(n_1134),
.B(n_1112),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1119),
.A2(n_1137),
.B(n_1132),
.Y(n_1142)
);

AO21x1_ASAP7_75t_L g1143 ( 
.A1(n_1047),
.A2(n_1019),
.B(n_1048),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_1116),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1064),
.B(n_1118),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1023),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1079),
.B(n_1010),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1112),
.B(n_1134),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_999),
.A2(n_1087),
.B(n_1059),
.C(n_1055),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1061),
.B(n_1040),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1051),
.A2(n_1043),
.B(n_1062),
.Y(n_1152)
);

OAI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1053),
.A2(n_1020),
.B(n_1069),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1111),
.A2(n_1074),
.B(n_990),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1002),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1050),
.A2(n_991),
.B(n_1115),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1035),
.Y(n_1157)
);

O2A1O1Ixp33_ASAP7_75t_SL g1158 ( 
.A1(n_1063),
.A2(n_1003),
.B(n_1029),
.C(n_1004),
.Y(n_1158)
);

AOI31xp67_ASAP7_75t_L g1159 ( 
.A1(n_1108),
.A2(n_1106),
.A3(n_1110),
.B(n_1107),
.Y(n_1159)
);

INVxp67_ASAP7_75t_L g1160 ( 
.A(n_1044),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1095),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1014),
.B(n_1091),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1110),
.A2(n_1047),
.A3(n_1090),
.B(n_1077),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1067),
.A2(n_1057),
.B(n_995),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1042),
.B(n_1128),
.Y(n_1165)
);

O2A1O1Ixp5_ASAP7_75t_SL g1166 ( 
.A1(n_1019),
.A2(n_1098),
.B(n_1073),
.C(n_1060),
.Y(n_1166)
);

AND2x4_ASAP7_75t_L g1167 ( 
.A(n_1128),
.B(n_996),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1034),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1054),
.B(n_1084),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_993),
.A2(n_1081),
.B(n_992),
.Y(n_1170)
);

HB1xp67_ASAP7_75t_L g1171 ( 
.A(n_1054),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1096),
.A2(n_1101),
.B(n_1001),
.Y(n_1172)
);

BUFx6f_ASAP7_75t_L g1173 ( 
.A(n_996),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1049),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1061),
.B(n_1040),
.Y(n_1175)
);

O2A1O1Ixp5_ASAP7_75t_L g1176 ( 
.A1(n_1103),
.A2(n_1086),
.B(n_1098),
.C(n_1060),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1017),
.A2(n_1025),
.B(n_1093),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1080),
.Y(n_1178)
);

NAND3xp33_ASAP7_75t_L g1179 ( 
.A(n_1000),
.B(n_1009),
.C(n_1083),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1093),
.A2(n_1088),
.B(n_1031),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1004),
.A2(n_1094),
.B(n_1033),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1073),
.A2(n_1104),
.A3(n_1066),
.B(n_1117),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1039),
.B(n_1030),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_996),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_994),
.A2(n_989),
.B(n_998),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1012),
.A2(n_1068),
.B(n_1018),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_SL g1187 ( 
.A(n_1036),
.B(n_1070),
.Y(n_1187)
);

NAND3xp33_ASAP7_75t_L g1188 ( 
.A(n_1006),
.B(n_1038),
.C(n_1032),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1024),
.A2(n_1026),
.B(n_1028),
.C(n_1085),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1008),
.B(n_1058),
.Y(n_1190)
);

BUFx2_ASAP7_75t_R g1191 ( 
.A(n_1015),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1008),
.A2(n_1105),
.B(n_1065),
.C(n_1007),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1123),
.B(n_1126),
.Y(n_1193)
);

BUFx2_ASAP7_75t_L g1194 ( 
.A(n_1027),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1133),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1076),
.A2(n_1100),
.B(n_1056),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1089),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1013),
.A2(n_1011),
.B(n_1120),
.Y(n_1198)
);

BUFx10_ASAP7_75t_L g1199 ( 
.A(n_1016),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1082),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1016),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1041),
.A2(n_1135),
.B(n_1113),
.C(n_1045),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1005),
.Y(n_1203)
);

NOR2x1_ASAP7_75t_SL g1204 ( 
.A(n_1092),
.B(n_1099),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1078),
.B(n_1052),
.Y(n_1205)
);

INVx5_ASAP7_75t_L g1206 ( 
.A(n_1097),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1016),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1102),
.B(n_1092),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_1022),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_997),
.B(n_1052),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1045),
.A2(n_1109),
.B(n_1037),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1109),
.A2(n_1127),
.B(n_1125),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1002),
.Y(n_1213)
);

BUFx3_ASAP7_75t_L g1214 ( 
.A(n_1023),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_1099),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1002),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1129),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1071),
.C(n_1136),
.Y(n_1220)
);

CKINVDCx6p67_ASAP7_75t_R g1221 ( 
.A(n_1027),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1222)
);

AND2x6_ASAP7_75t_L g1223 ( 
.A(n_1008),
.B(n_816),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1136),
.B(n_423),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1136),
.B(n_734),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1021),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1071),
.C(n_1136),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_SL g1229 ( 
.A1(n_1121),
.A2(n_1122),
.B1(n_1000),
.B2(n_1003),
.C(n_1112),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1118),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_996),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1129),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1237)
);

BUFx3_ASAP7_75t_L g1238 ( 
.A(n_1023),
.Y(n_1238)
);

AO32x2_ASAP7_75t_L g1239 ( 
.A1(n_1129),
.A2(n_1047),
.A3(n_1060),
.B1(n_1040),
.B2(n_1073),
.Y(n_1239)
);

NAND2x2_ASAP7_75t_L g1240 ( 
.A(n_1023),
.B(n_676),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1136),
.B(n_423),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1092),
.B(n_1093),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1128),
.B(n_817),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1118),
.B(n_1130),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1002),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1002),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1046),
.A2(n_836),
.B1(n_765),
.B2(n_734),
.Y(n_1251)
);

O2A1O1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1136),
.C(n_423),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1002),
.Y(n_1253)
);

AO31x2_ASAP7_75t_L g1254 ( 
.A1(n_1115),
.A2(n_889),
.A3(n_1110),
.B(n_1111),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_996),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1023),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1136),
.B(n_423),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1023),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1115),
.A2(n_889),
.A3(n_1110),
.B(n_1111),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1002),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1136),
.B(n_423),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1115),
.A2(n_1048),
.B(n_1055),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1267)
);

O2A1O1Ixp33_ASAP7_75t_L g1268 ( 
.A1(n_1122),
.A2(n_1121),
.B(n_1136),
.C(n_423),
.Y(n_1268)
);

BUFx3_ASAP7_75t_L g1269 ( 
.A(n_1023),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1112),
.B(n_1134),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1129),
.A2(n_836),
.B1(n_734),
.B2(n_925),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1112),
.B(n_1134),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1108),
.A2(n_1111),
.B(n_1074),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1124),
.B(n_1131),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1121),
.A2(n_1132),
.B(n_1119),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_996),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1134),
.C(n_1112),
.Y(n_1279)
);

INVxp67_ASAP7_75t_SL g1280 ( 
.A(n_1054),
.Y(n_1280)
);

OAI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1130),
.A2(n_1009),
.B1(n_1079),
.B2(n_1008),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1125),
.A2(n_1127),
.B(n_1072),
.Y(n_1282)
);

AO31x2_ASAP7_75t_L g1283 ( 
.A1(n_1115),
.A2(n_889),
.A3(n_1110),
.B(n_1111),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1155),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1157),
.Y(n_1285)
);

OAI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1147),
.A2(n_1140),
.B(n_1138),
.Y(n_1286)
);

CKINVDCx8_ASAP7_75t_R g1287 ( 
.A(n_1209),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1223),
.A2(n_1179),
.B1(n_1190),
.B2(n_1185),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1251),
.A2(n_1271),
.B1(n_1143),
.B2(n_1281),
.Y(n_1289)
);

INVxp67_ASAP7_75t_L g1290 ( 
.A(n_1183),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1138),
.A2(n_1271),
.B1(n_1227),
.B2(n_1220),
.Y(n_1291)
);

BUFx12f_ASAP7_75t_L g1292 ( 
.A(n_1144),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1196),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1179),
.A2(n_1223),
.B1(n_1185),
.B2(n_1139),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1225),
.A2(n_1236),
.B1(n_1218),
.B2(n_1188),
.Y(n_1295)
);

BUFx12f_ASAP7_75t_L g1296 ( 
.A(n_1195),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1223),
.A2(n_1218),
.B1(n_1236),
.B2(n_1188),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1213),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1223),
.B1(n_1235),
.B2(n_1244),
.Y(n_1299)
);

INVx6_ASAP7_75t_L g1300 ( 
.A(n_1206),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1247),
.A2(n_1187),
.B1(n_1262),
.B2(n_1267),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1159),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1221),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_SL g1304 ( 
.A1(n_1210),
.A2(n_1245),
.B1(n_1265),
.B2(n_1151),
.Y(n_1304)
);

AOI21xp33_ASAP7_75t_L g1305 ( 
.A1(n_1229),
.A2(n_1150),
.B(n_1189),
.Y(n_1305)
);

CKINVDCx6p67_ASAP7_75t_R g1306 ( 
.A(n_1203),
.Y(n_1306)
);

CKINVDCx11_ASAP7_75t_R g1307 ( 
.A(n_1240),
.Y(n_1307)
);

BUFx4f_ASAP7_75t_SL g1308 ( 
.A(n_1146),
.Y(n_1308)
);

BUFx2_ASAP7_75t_SL g1309 ( 
.A(n_1214),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1243),
.A2(n_1276),
.B1(n_1233),
.B2(n_1141),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1224),
.B(n_1241),
.Y(n_1311)
);

HB1xp67_ASAP7_75t_L g1312 ( 
.A(n_1233),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1257),
.B(n_1264),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1256),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1217),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1145),
.B(n_1160),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1141),
.A2(n_1151),
.B1(n_1175),
.B2(n_1250),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1175),
.A2(n_1249),
.B1(n_1253),
.B2(n_1263),
.Y(n_1318)
);

INVx3_ASAP7_75t_L g1319 ( 
.A(n_1173),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1238),
.Y(n_1320)
);

CKINVDCx11_ASAP7_75t_R g1321 ( 
.A(n_1194),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1161),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_L g1323 ( 
.A(n_1246),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1258),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1252),
.A2(n_1268),
.B1(n_1280),
.B2(n_1169),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1165),
.B(n_1246),
.Y(n_1326)
);

BUFx2_ASAP7_75t_SL g1327 ( 
.A(n_1269),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1168),
.A2(n_1174),
.B1(n_1178),
.B2(n_1198),
.Y(n_1328)
);

OAI22x1_ASAP7_75t_L g1329 ( 
.A1(n_1207),
.A2(n_1201),
.B1(n_1171),
.B2(n_1200),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1193),
.A2(n_1148),
.B1(n_1270),
.B2(n_1272),
.Y(n_1330)
);

CKINVDCx11_ASAP7_75t_R g1331 ( 
.A(n_1184),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1226),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1198),
.A2(n_1153),
.B1(n_1180),
.B2(n_1148),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1153),
.A2(n_1204),
.B1(n_1239),
.B2(n_1186),
.Y(n_1334)
);

BUFx2_ASAP7_75t_SL g1335 ( 
.A(n_1167),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1184),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1184),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1270),
.A2(n_1272),
.B1(n_1192),
.B2(n_1232),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1181),
.A2(n_1248),
.B1(n_1242),
.B2(n_1277),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1197),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1197),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1239),
.A2(n_1205),
.B1(n_1199),
.B2(n_1208),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1219),
.A2(n_1259),
.B1(n_1237),
.B2(n_1273),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_1234),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1216),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1208),
.Y(n_1346)
);

BUFx2_ASAP7_75t_SL g1347 ( 
.A(n_1234),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1216),
.A2(n_1255),
.B1(n_1234),
.B2(n_1278),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1182),
.Y(n_1349)
);

BUFx10_ASAP7_75t_L g1350 ( 
.A(n_1255),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1182),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1278),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1182),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1230),
.A2(n_1266),
.B1(n_1261),
.B2(n_1239),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1191),
.A2(n_1142),
.B1(n_1164),
.B2(n_1156),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1279),
.B(n_1229),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1202),
.B(n_1158),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_1212),
.Y(n_1358)
);

CKINVDCx6p67_ASAP7_75t_R g1359 ( 
.A(n_1211),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1211),
.A2(n_1166),
.B1(n_1177),
.B2(n_1154),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1274),
.A2(n_1176),
.B1(n_1163),
.B2(n_1172),
.Y(n_1361)
);

BUFx8_ASAP7_75t_SL g1362 ( 
.A(n_1254),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1163),
.Y(n_1363)
);

CKINVDCx6p67_ASAP7_75t_R g1364 ( 
.A(n_1254),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1254),
.Y(n_1365)
);

AOI22xp5_ASAP7_75t_L g1366 ( 
.A1(n_1170),
.A2(n_1149),
.B1(n_1282),
.B2(n_1215),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1152),
.A2(n_1222),
.B1(n_1228),
.B2(n_1231),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1275),
.A2(n_1260),
.B(n_1283),
.Y(n_1368)
);

CKINVDCx11_ASAP7_75t_R g1369 ( 
.A(n_1260),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1283),
.A2(n_1147),
.B1(n_836),
.B2(n_745),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1147),
.A2(n_1138),
.B1(n_1271),
.B2(n_1121),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1256),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1146),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1221),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1155),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1173),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_1144),
.Y(n_1377)
);

OAI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1271),
.A2(n_1138),
.B1(n_1147),
.B2(n_1129),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_1280),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1251),
.A2(n_836),
.B1(n_1147),
.B2(n_1271),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_SL g1381 ( 
.A1(n_1147),
.A2(n_501),
.B1(n_1225),
.B2(n_1138),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1155),
.Y(n_1382)
);

BUFx2_ASAP7_75t_R g1383 ( 
.A(n_1209),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1173),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1256),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1155),
.Y(n_1386)
);

INVx3_ASAP7_75t_SL g1387 ( 
.A(n_1209),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1251),
.A2(n_836),
.B1(n_1147),
.B2(n_1271),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1147),
.A2(n_734),
.B1(n_1271),
.B2(n_1251),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1251),
.A2(n_836),
.B1(n_1147),
.B2(n_1271),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1155),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1251),
.A2(n_836),
.B1(n_1147),
.B2(n_1271),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1183),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1147),
.A2(n_1138),
.B1(n_1271),
.B2(n_1121),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1251),
.A2(n_836),
.B1(n_1147),
.B2(n_1271),
.Y(n_1395)
);

BUFx8_ASAP7_75t_SL g1396 ( 
.A(n_1203),
.Y(n_1396)
);

BUFx8_ASAP7_75t_L g1397 ( 
.A(n_1144),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1271),
.A2(n_1138),
.B1(n_1147),
.B2(n_1129),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1349),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1351),
.Y(n_1400)
);

INVx4_ASAP7_75t_L g1401 ( 
.A(n_1359),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1308),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1353),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1317),
.B(n_1363),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1341),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1330),
.B(n_1316),
.Y(n_1406)
);

AOI21xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1286),
.A2(n_1295),
.B(n_1371),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1312),
.Y(n_1409)
);

AO21x2_ASAP7_75t_L g1410 ( 
.A1(n_1368),
.A2(n_1302),
.B(n_1361),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1358),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1365),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1298),
.B(n_1315),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1364),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1340),
.Y(n_1415)
);

INVx4_ASAP7_75t_L g1416 ( 
.A(n_1300),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1375),
.Y(n_1417)
);

OAI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1389),
.A2(n_1381),
.B1(n_1294),
.B2(n_1289),
.C(n_1392),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1382),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1379),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1300),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1339),
.A2(n_1343),
.B(n_1367),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1339),
.A2(n_1343),
.B(n_1367),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1386),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1357),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1293),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1391),
.Y(n_1427)
);

BUFx2_ASAP7_75t_L g1428 ( 
.A(n_1362),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1322),
.Y(n_1429)
);

HB1xp67_ASAP7_75t_L g1430 ( 
.A(n_1346),
.Y(n_1430)
);

INVx4_ASAP7_75t_SL g1431 ( 
.A(n_1300),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1354),
.A2(n_1360),
.B(n_1366),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1318),
.B(n_1310),
.Y(n_1433)
);

AND2x6_ASAP7_75t_SL g1434 ( 
.A(n_1311),
.B(n_1313),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1318),
.B(n_1310),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1338),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1332),
.Y(n_1437)
);

BUFx6f_ASAP7_75t_L g1438 ( 
.A(n_1369),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1356),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1369),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1288),
.A2(n_1388),
.B1(n_1380),
.B2(n_1390),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1333),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1290),
.B(n_1393),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1354),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1329),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1334),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1360),
.A2(n_1355),
.B(n_1291),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1328),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1326),
.Y(n_1449)
);

INVx8_ASAP7_75t_L g1450 ( 
.A(n_1336),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1328),
.Y(n_1451)
);

INVxp67_ASAP7_75t_L g1452 ( 
.A(n_1314),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1297),
.A2(n_1394),
.B(n_1294),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1297),
.B(n_1301),
.Y(n_1454)
);

OAI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1325),
.A2(n_1289),
.B(n_1319),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1378),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1378),
.A2(n_1398),
.B(n_1305),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1398),
.B(n_1301),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1299),
.B(n_1380),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1342),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1323),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1304),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1308),
.B(n_1320),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1370),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1395),
.B(n_1385),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1345),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1348),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1337),
.A2(n_1344),
.B1(n_1352),
.B2(n_1296),
.Y(n_1469)
);

BUFx2_ASAP7_75t_L g1470 ( 
.A(n_1467),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1409),
.B(n_1373),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1430),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1458),
.B(n_1327),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1415),
.B(n_1309),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1436),
.B(n_1324),
.Y(n_1475)
);

OAI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1407),
.A2(n_1384),
.B(n_1376),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1420),
.B(n_1324),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1401),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1418),
.A2(n_1335),
.B1(n_1331),
.B2(n_1307),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1466),
.B(n_1321),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1466),
.B(n_1321),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_SL g1482 ( 
.A1(n_1406),
.A2(n_1307),
.B(n_1396),
.Y(n_1482)
);

NAND4xp25_ASAP7_75t_L g1483 ( 
.A(n_1439),
.B(n_1452),
.C(n_1436),
.D(n_1441),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1438),
.B(n_1374),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1405),
.B(n_1306),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1442),
.A2(n_1303),
.B1(n_1387),
.B2(n_1347),
.C(n_1383),
.Y(n_1486)
);

A2O1A1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1453),
.A2(n_1292),
.B(n_1296),
.C(n_1377),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1408),
.B(n_1387),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1438),
.B(n_1397),
.Y(n_1489)
);

OR2x2_ASAP7_75t_L g1490 ( 
.A(n_1417),
.B(n_1396),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1408),
.B(n_1413),
.Y(n_1491)
);

AND2x4_ASAP7_75t_L g1492 ( 
.A(n_1438),
.B(n_1397),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1457),
.A2(n_1350),
.B(n_1377),
.Y(n_1493)
);

AOI221xp5_ASAP7_75t_L g1494 ( 
.A1(n_1442),
.A2(n_1287),
.B1(n_1292),
.B2(n_1350),
.C(n_1456),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1413),
.B(n_1404),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1465),
.A2(n_1454),
.B1(n_1463),
.B2(n_1457),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1439),
.B(n_1456),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1404),
.B(n_1444),
.Y(n_1498)
);

NOR2xp67_ASAP7_75t_L g1499 ( 
.A(n_1401),
.B(n_1469),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1438),
.B(n_1414),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1417),
.B(n_1419),
.Y(n_1501)
);

OA21x2_ASAP7_75t_L g1502 ( 
.A1(n_1447),
.A2(n_1422),
.B(n_1423),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1440),
.B(n_1428),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1457),
.A2(n_1447),
.B(n_1422),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1459),
.A2(n_1465),
.B(n_1460),
.C(n_1454),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1444),
.B(n_1425),
.Y(n_1506)
);

AO32x2_ASAP7_75t_L g1507 ( 
.A1(n_1401),
.A2(n_1421),
.A3(n_1416),
.B1(n_1434),
.B2(n_1433),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1402),
.B(n_1464),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1419),
.B(n_1424),
.Y(n_1509)
);

O2A1O1Ixp5_ASAP7_75t_L g1510 ( 
.A1(n_1446),
.A2(n_1459),
.B(n_1463),
.C(n_1412),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1460),
.A2(n_1446),
.B(n_1455),
.C(n_1433),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1425),
.B(n_1427),
.Y(n_1512)
);

A2O1A1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1455),
.A2(n_1435),
.B(n_1461),
.C(n_1448),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1425),
.B(n_1429),
.Y(n_1514)
);

OAI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1448),
.A2(n_1451),
.B(n_1435),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1491),
.B(n_1432),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1495),
.B(n_1502),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1502),
.B(n_1410),
.Y(n_1518)
);

CKINVDCx5p33_ASAP7_75t_R g1519 ( 
.A(n_1470),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1498),
.B(n_1432),
.Y(n_1520)
);

NAND3xp33_ASAP7_75t_L g1521 ( 
.A(n_1504),
.B(n_1432),
.C(n_1443),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1512),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1500),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1496),
.A2(n_1468),
.B1(n_1445),
.B2(n_1449),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_SL g1525 ( 
.A(n_1476),
.B(n_1462),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1498),
.B(n_1412),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1512),
.B(n_1426),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1497),
.B(n_1472),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1501),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1514),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1507),
.Y(n_1531)
);

INVxp67_ASAP7_75t_R g1532 ( 
.A(n_1476),
.Y(n_1532)
);

AOI222xp33_ASAP7_75t_L g1533 ( 
.A1(n_1505),
.A2(n_1450),
.B1(n_1431),
.B2(n_1399),
.C1(n_1403),
.C2(n_1400),
.Y(n_1533)
);

HB1xp67_ASAP7_75t_L g1534 ( 
.A(n_1506),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1509),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1506),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1483),
.A2(n_1450),
.B1(n_1437),
.B2(n_1399),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1507),
.B(n_1411),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1507),
.B(n_1411),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1522),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1490),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1517),
.B(n_1507),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1522),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1530),
.Y(n_1544)
);

OAI22xp5_ASAP7_75t_SL g1545 ( 
.A1(n_1531),
.A2(n_1489),
.B1(n_1492),
.B2(n_1484),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1523),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1547)
);

AOI33xp33_ASAP7_75t_L g1548 ( 
.A1(n_1537),
.A2(n_1481),
.A3(n_1486),
.B1(n_1479),
.B2(n_1471),
.B3(n_1473),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1488),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1516),
.B(n_1475),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1538),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1531),
.B(n_1520),
.Y(n_1553)
);

OAI21xp33_ASAP7_75t_L g1554 ( 
.A1(n_1521),
.A2(n_1511),
.B(n_1513),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1518),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1519),
.B(n_1474),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1518),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1538),
.B(n_1503),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1530),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1518),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1531),
.B(n_1477),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1534),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1534),
.Y(n_1563)
);

NAND2x1_ASAP7_75t_L g1564 ( 
.A(n_1539),
.B(n_1492),
.Y(n_1564)
);

OAI21xp33_ASAP7_75t_L g1565 ( 
.A1(n_1521),
.A2(n_1524),
.B(n_1537),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1540),
.B(n_1536),
.Y(n_1566)
);

BUFx2_ASAP7_75t_L g1567 ( 
.A(n_1552),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1540),
.B(n_1536),
.Y(n_1568)
);

BUFx3_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1542),
.B(n_1539),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1539),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1543),
.B(n_1536),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1552),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1543),
.B(n_1529),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1552),
.B(n_1532),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1541),
.B(n_1528),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1532),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1544),
.B(n_1529),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1544),
.B(n_1559),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1547),
.B(n_1532),
.Y(n_1580)
);

OR2x2_ASAP7_75t_L g1581 ( 
.A(n_1553),
.B(n_1526),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1549),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1529),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1546),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1553),
.B(n_1526),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1547),
.B(n_1527),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1564),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1562),
.B(n_1535),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1546),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1562),
.B(n_1535),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

OR2x6_ASAP7_75t_SL g1593 ( 
.A(n_1579),
.B(n_1485),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1569),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1574),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1569),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1573),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1588),
.B(n_1561),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1574),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1578),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1569),
.Y(n_1603)
);

A2O1A1Ixp33_ASAP7_75t_L g1604 ( 
.A1(n_1576),
.A2(n_1565),
.B(n_1554),
.C(n_1548),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1588),
.B(n_1561),
.Y(n_1606)
);

NAND2x1_ASAP7_75t_SL g1607 ( 
.A(n_1575),
.B(n_1563),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1578),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1583),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1583),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1576),
.B(n_1551),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1589),
.Y(n_1612)
);

AOI32xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1579),
.A2(n_1541),
.A3(n_1556),
.B1(n_1508),
.B2(n_1551),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1561),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1589),
.Y(n_1615)
);

NAND2x1p5_ASAP7_75t_L g1616 ( 
.A(n_1569),
.B(n_1525),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1591),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1573),
.Y(n_1619)
);

INVx2_ASAP7_75t_SL g1620 ( 
.A(n_1587),
.Y(n_1620)
);

AOI211xp5_ASAP7_75t_L g1621 ( 
.A1(n_1584),
.A2(n_1565),
.B(n_1554),
.C(n_1499),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1591),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1570),
.A2(n_1524),
.B1(n_1515),
.B2(n_1533),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1566),
.Y(n_1624)
);

AOI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1570),
.A2(n_1524),
.B1(n_1533),
.B2(n_1520),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1581),
.B(n_1563),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1582),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1587),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1584),
.B(n_1548),
.Y(n_1629)
);

AND2x4_ASAP7_75t_L g1630 ( 
.A(n_1587),
.B(n_1590),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1566),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1570),
.B(n_1558),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1581),
.B(n_1528),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1581),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1575),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1590),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1556),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1634),
.B(n_1585),
.Y(n_1638)
);

NAND3x1_ASAP7_75t_L g1639 ( 
.A(n_1629),
.B(n_1486),
.C(n_1575),
.Y(n_1639)
);

INVx2_ASAP7_75t_L g1640 ( 
.A(n_1597),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1598),
.B(n_1571),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1585),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1597),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1626),
.B(n_1585),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1601),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1626),
.B(n_1568),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1605),
.B(n_1571),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1599),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1622),
.Y(n_1649)
);

OR2x2_ASAP7_75t_L g1650 ( 
.A(n_1633),
.B(n_1568),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1605),
.B(n_1571),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1618),
.B(n_1632),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1624),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1633),
.B(n_1572),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1631),
.B(n_1611),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1602),
.B(n_1572),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1599),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1587),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1632),
.B(n_1577),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1621),
.A2(n_1487),
.B(n_1577),
.C(n_1545),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1602),
.B(n_1592),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1593),
.B(n_1577),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1601),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1593),
.B(n_1586),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1619),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1596),
.B(n_1564),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1623),
.A2(n_1510),
.B(n_1493),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1606),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1606),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1608),
.B(n_1582),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1625),
.B(n_1545),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1637),
.B(n_1594),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1637),
.B(n_1648),
.Y(n_1673)
);

AOI221xp5_ASAP7_75t_L g1674 ( 
.A1(n_1671),
.A2(n_1609),
.B1(n_1610),
.B2(n_1612),
.C(n_1608),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1648),
.Y(n_1675)
);

A2O1A1Ixp33_ASAP7_75t_L g1676 ( 
.A1(n_1667),
.A2(n_1607),
.B(n_1613),
.C(n_1614),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1657),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1667),
.A2(n_1610),
.B1(n_1612),
.B2(n_1609),
.C(n_1615),
.Y(n_1678)
);

INVxp67_ASAP7_75t_L g1679 ( 
.A(n_1657),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1668),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1664),
.B(n_1596),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1655),
.A2(n_1614),
.A3(n_1613),
.B1(n_1616),
.B2(n_1635),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1662),
.A2(n_1607),
.B(n_1603),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1668),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1669),
.Y(n_1685)
);

OAI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1662),
.A2(n_1600),
.B(n_1595),
.Y(n_1686)
);

OAI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1639),
.A2(n_1616),
.B1(n_1560),
.B2(n_1549),
.C(n_1555),
.Y(n_1687)
);

AOI21xp33_ASAP7_75t_SL g1688 ( 
.A1(n_1655),
.A2(n_1616),
.B(n_1620),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1669),
.B(n_1617),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1664),
.B(n_1630),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1649),
.B(n_1615),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1649),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1652),
.B(n_1630),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1636),
.B(n_1619),
.Y(n_1695)
);

OAI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1639),
.A2(n_1520),
.B1(n_1549),
.B2(n_1555),
.Y(n_1696)
);

OAI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1653),
.A2(n_1628),
.B(n_1620),
.C(n_1567),
.Y(n_1697)
);

NAND3x2_ASAP7_75t_L g1698 ( 
.A(n_1690),
.B(n_1644),
.C(n_1653),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1675),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1672),
.B(n_1673),
.Y(n_1700)
);

INVxp33_ASAP7_75t_L g1701 ( 
.A(n_1690),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1692),
.B(n_1636),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1692),
.B(n_1641),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1676),
.A2(n_1639),
.B(n_1660),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

OR2x2_ASAP7_75t_L g1706 ( 
.A(n_1695),
.B(n_1644),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1694),
.B(n_1641),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1680),
.Y(n_1708)
);

O2A1O1Ixp5_ASAP7_75t_L g1709 ( 
.A1(n_1682),
.A2(n_1640),
.B(n_1643),
.C(n_1665),
.Y(n_1709)
);

AOI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1678),
.A2(n_1656),
.B1(n_1640),
.B2(n_1643),
.C(n_1665),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1696),
.A2(n_1660),
.B1(n_1643),
.B2(n_1665),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1694),
.B(n_1646),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1695),
.B(n_1638),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1681),
.B(n_1647),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1684),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1685),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1687),
.A2(n_1674),
.B1(n_1676),
.B2(n_1683),
.Y(n_1717)
);

INVxp33_ASAP7_75t_L g1718 ( 
.A(n_1712),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1707),
.B(n_1679),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1682),
.Y(n_1720)
);

XOR2x2_ASAP7_75t_L g1721 ( 
.A(n_1704),
.B(n_1691),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1706),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1713),
.Y(n_1723)
);

NOR2xp67_ASAP7_75t_L g1724 ( 
.A(n_1702),
.B(n_1697),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1714),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1704),
.A2(n_1681),
.B1(n_1686),
.B2(n_1645),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1698),
.B(n_1638),
.Y(n_1727)
);

XNOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1717),
.B(n_1693),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1718),
.B(n_1703),
.Y(n_1729)
);

OAI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1720),
.A2(n_1709),
.B(n_1700),
.Y(n_1730)
);

NAND4xp25_ASAP7_75t_L g1731 ( 
.A(n_1724),
.B(n_1709),
.C(n_1699),
.D(n_1707),
.Y(n_1731)
);

NOR4xp75_ASAP7_75t_SL g1732 ( 
.A(n_1726),
.B(n_1689),
.C(n_1656),
.D(n_1661),
.Y(n_1732)
);

OAI21xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1728),
.A2(n_1727),
.B(n_1722),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_SL g1734 ( 
.A(n_1721),
.B(n_1710),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1723),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1719),
.B(n_1710),
.C(n_1711),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1725),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1719),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1731),
.A2(n_1730),
.B(n_1732),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1729),
.B(n_1647),
.Y(n_1740)
);

NAND2x1_ASAP7_75t_L g1741 ( 
.A(n_1738),
.B(n_1735),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1734),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1734),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1737),
.Y(n_1745)
);

AOI22xp5_ASAP7_75t_L g1746 ( 
.A1(n_1742),
.A2(n_1736),
.B1(n_1716),
.B2(n_1715),
.Y(n_1746)
);

OAI311xp33_ASAP7_75t_L g1747 ( 
.A1(n_1739),
.A2(n_1708),
.A3(n_1642),
.B1(n_1646),
.C1(n_1650),
.Y(n_1747)
);

A2O1A1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1742),
.A2(n_1688),
.B(n_1645),
.C(n_1663),
.Y(n_1748)
);

OAI211xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1744),
.A2(n_1640),
.B(n_1663),
.C(n_1645),
.Y(n_1749)
);

AOI222xp33_ASAP7_75t_L g1750 ( 
.A1(n_1743),
.A2(n_1663),
.B1(n_1670),
.B2(n_1661),
.C1(n_1627),
.C2(n_1651),
.Y(n_1750)
);

NOR3xp33_ASAP7_75t_L g1751 ( 
.A(n_1741),
.B(n_1670),
.C(n_1642),
.Y(n_1751)
);

AOI222xp33_ASAP7_75t_L g1752 ( 
.A1(n_1745),
.A2(n_1627),
.B1(n_1651),
.B2(n_1560),
.C1(n_1557),
.C2(n_1555),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1746),
.A2(n_1740),
.B1(n_1666),
.B2(n_1658),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1749),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1751),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1748),
.B(n_1658),
.Y(n_1756)
);

NOR2xp67_ASAP7_75t_L g1757 ( 
.A(n_1747),
.B(n_1628),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1754),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1757),
.B(n_1750),
.Y(n_1759)
);

NOR2x1p5_ASAP7_75t_L g1760 ( 
.A(n_1755),
.B(n_1650),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1760),
.Y(n_1761)
);

OAI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1761),
.A2(n_1759),
.B1(n_1753),
.B2(n_1756),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1762),
.Y(n_1763)
);

XNOR2x1_ASAP7_75t_L g1764 ( 
.A(n_1762),
.B(n_1758),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1763),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1764),
.A2(n_1752),
.B(n_1666),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1765),
.A2(n_1766),
.B1(n_1659),
.B2(n_1484),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1765),
.Y(n_1768)
);

AOI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1768),
.A2(n_1654),
.B(n_1659),
.Y(n_1769)
);

OAI21xp33_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1767),
.B(n_1654),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1770),
.Y(n_1771)
);

OAI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1771),
.A2(n_1567),
.B1(n_1482),
.B2(n_1478),
.C(n_1582),
.Y(n_1772)
);

AOI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1493),
.B(n_1494),
.C(n_1592),
.Y(n_1773)
);


endmodule