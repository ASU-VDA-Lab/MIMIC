module fake_jpeg_3600_n_471 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_471);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_471;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_56),
.Y(n_156)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_21),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_59),
.B(n_104),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_60),
.Y(n_183)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_61),
.Y(n_120)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_64),
.Y(n_151)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_68),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_21),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_77),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_71),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_SL g72 ( 
.A1(n_33),
.A2(n_17),
.B(n_16),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g165 ( 
.A1(n_72),
.A2(n_36),
.B(n_5),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_48),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_113),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_75),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_54),
.A2(n_55),
.B1(n_29),
.B2(n_38),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_76),
.A2(n_23),
.B1(n_43),
.B2(n_41),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_31),
.B(n_52),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_18),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_79),
.A2(n_40),
.B1(n_25),
.B2(n_53),
.Y(n_140)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_81),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_31),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_82),
.B(n_108),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_83),
.Y(n_174)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_86),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_89),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_92),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_99),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_102),
.B(n_103),
.Y(n_149)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_106),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_35),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_1),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_26),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_114),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_111),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_27),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_82),
.B(n_53),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_124),
.B(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_131),
.A2(n_135),
.B1(n_124),
.B2(n_151),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_78),
.A2(n_24),
.B1(n_43),
.B2(n_41),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_76),
.A2(n_40),
.B1(n_25),
.B2(n_24),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_137),
.A2(n_140),
.B1(n_163),
.B2(n_175),
.Y(n_201)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_70),
.A2(n_27),
.B(n_22),
.C(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_143),
.B(n_164),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_114),
.A2(n_37),
.B1(n_30),
.B2(n_20),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_150),
.A2(n_153),
.B1(n_119),
.B2(n_171),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_77),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_152),
.B(n_157),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_99),
.A2(n_37),
.B1(n_30),
.B2(n_20),
.Y(n_153)
);

CKINVDCx12_ASAP7_75t_R g154 ( 
.A(n_96),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_154),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_2),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_3),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_112),
.B(n_3),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_37),
.B1(n_36),
.B2(n_22),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_73),
.A2(n_22),
.B(n_36),
.C(n_6),
.Y(n_164)
);

NOR2x1_ASAP7_75t_R g244 ( 
.A(n_165),
.B(n_177),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_101),
.B(n_10),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_166),
.B(n_179),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_56),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_85),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_178),
.A2(n_188),
.B1(n_153),
.B2(n_150),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_104),
.B(n_7),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_7),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_114),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_9),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_184),
.B(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_60),
.B(n_67),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_87),
.B(n_68),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_69),
.A2(n_71),
.B1(n_89),
.B2(n_90),
.Y(n_188)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_93),
.B1(n_100),
.B2(n_102),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_192),
.A2(n_215),
.B1(n_226),
.B2(n_228),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_126),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_197),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_199),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_117),
.B(n_111),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_234),
.Y(n_267)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_202),
.Y(n_270)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_203),
.Y(n_291)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_189),
.B(n_113),
.CI(n_143),
.CON(n_205),
.SN(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_206),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_207),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_131),
.A2(n_135),
.B1(n_164),
.B2(n_180),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_209),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_180),
.A2(n_181),
.B1(n_161),
.B2(n_172),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_211),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_136),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_212),
.B(n_230),
.C(n_244),
.Y(n_290)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_132),
.Y(n_213)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_214),
.A2(n_219),
.B1(n_220),
.B2(n_225),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_171),
.B1(n_170),
.B2(n_119),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_122),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_218),
.Y(n_284)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_186),
.A2(n_125),
.B1(n_139),
.B2(n_138),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_221),
.B(n_224),
.Y(n_259)
);

AO22x1_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_237),
.B1(n_201),
.B2(n_235),
.Y(n_255)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_149),
.A2(n_159),
.B1(n_162),
.B2(n_151),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_159),
.A2(n_149),
.B1(n_162),
.B2(n_183),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_128),
.A2(n_190),
.B1(n_118),
.B2(n_123),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_227),
.A2(n_235),
.B1(n_237),
.B2(n_241),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_142),
.A2(n_146),
.B1(n_127),
.B2(n_149),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_129),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_229),
.B(n_245),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_133),
.B(n_141),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_147),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.Y(n_262)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_123),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_155),
.B(n_185),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_155),
.A2(n_185),
.B1(n_168),
.B2(n_183),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_147),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_236),
.B(n_238),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_168),
.A2(n_141),
.B1(n_144),
.B2(n_174),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_144),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_174),
.A2(n_130),
.B1(n_148),
.B2(n_132),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_130),
.A2(n_148),
.B1(n_167),
.B2(n_120),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_130),
.A2(n_148),
.B1(n_167),
.B2(n_120),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_167),
.B(n_147),
.Y(n_242)
);

OR2x6_ASAP7_75t_SL g257 ( 
.A(n_242),
.B(n_244),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_173),
.A2(n_145),
.B1(n_117),
.B2(n_137),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_243),
.A2(n_252),
.B1(n_195),
.B2(n_207),
.Y(n_298)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_173),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_177),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_125),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_248),
.B(n_217),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_131),
.A2(n_163),
.B1(n_37),
.B2(n_135),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_251),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_145),
.A2(n_117),
.B1(n_137),
.B2(n_189),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_200),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_254),
.B(n_267),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_255),
.A2(n_274),
.B1(n_281),
.B2(n_260),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_256),
.A2(n_247),
.B1(n_224),
.B2(n_236),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_257),
.Y(n_320)
);

O2A1O1Ixp33_ASAP7_75t_SL g261 ( 
.A1(n_216),
.A2(n_205),
.B(n_223),
.C(n_219),
.Y(n_261)
);

A2O1A1O1Ixp25_ASAP7_75t_L g300 ( 
.A1(n_261),
.A2(n_257),
.B(n_272),
.C(n_258),
.D(n_267),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_242),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_282),
.Y(n_306)
);

OAI32xp33_ASAP7_75t_L g273 ( 
.A1(n_194),
.A2(n_205),
.A3(n_208),
.B1(n_249),
.B2(n_193),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_277),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_222),
.A2(n_234),
.B1(n_226),
.B2(n_197),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_223),
.A2(n_218),
.B(n_229),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_296),
.B(n_271),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_202),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_199),
.B(n_206),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_287),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_223),
.A2(n_239),
.B1(n_233),
.B2(n_204),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_213),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_225),
.B(n_196),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_191),
.B(n_238),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_231),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_298),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_203),
.B(n_245),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_246),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_282),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_299),
.A2(n_300),
.B(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_301),
.Y(n_335)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_305),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_307),
.B(n_286),
.Y(n_352)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_278),
.B(n_258),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_310),
.B(n_312),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_254),
.B(n_274),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_275),
.B(n_293),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_314),
.B(n_315),
.Y(n_357)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_266),
.B1(n_298),
.B2(n_276),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_326),
.B1(n_291),
.B2(n_253),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_275),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_284),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_322),
.Y(n_355)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_257),
.B(n_261),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_321),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_284),
.Y(n_322)
);

BUFx8_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

INVx11_ASAP7_75t_L g363 ( 
.A(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_284),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_324),
.B(n_327),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_325),
.Y(n_344)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_280),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_328),
.B(n_329),
.Y(n_360)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_280),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_255),
.A2(n_266),
.B1(n_281),
.B2(n_260),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_330),
.A2(n_334),
.B1(n_294),
.B2(n_264),
.Y(n_340)
);

OR2x4_ASAP7_75t_L g331 ( 
.A(n_261),
.B(n_290),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_331),
.B(n_332),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_263),
.B(n_262),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_289),
.B(n_269),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_333),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_255),
.A2(n_283),
.B1(n_294),
.B2(n_256),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_323),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_361),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_264),
.B(n_296),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_337),
.A2(n_351),
.B(n_308),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_307),
.B(n_285),
.C(n_259),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_346),
.C(n_347),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_340),
.A2(n_311),
.B1(n_305),
.B2(n_304),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_343),
.A2(n_334),
.B1(n_330),
.B2(n_326),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_320),
.B(n_285),
.C(n_268),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_268),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_323),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_349),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_320),
.A2(n_291),
.B(n_288),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_352),
.B(n_347),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_303),
.B(n_288),
.C(n_286),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_356),
.B(n_362),
.C(n_324),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_323),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_303),
.B(n_292),
.C(n_253),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_318),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_381),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_357),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_370),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_367),
.A2(n_371),
.B(n_375),
.Y(n_388)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_360),
.Y(n_368)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_369),
.B(n_353),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_349),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_331),
.B(n_317),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_373),
.A2(n_376),
.B1(n_378),
.B2(n_386),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_354),
.B(n_301),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_379),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_341),
.A2(n_321),
.B(n_313),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_351),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_354),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_340),
.A2(n_311),
.B1(n_302),
.B2(n_316),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_357),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_357),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_385),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_358),
.B(n_316),
.Y(n_383)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_383),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_339),
.B(n_321),
.C(n_306),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_346),
.C(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_349),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_343),
.A2(n_302),
.B1(n_306),
.B2(n_332),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_372),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_387),
.B(n_393),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_389),
.B(n_391),
.C(n_404),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_338),
.C(n_362),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_373),
.A2(n_337),
.B1(n_335),
.B2(n_359),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_376),
.B1(n_365),
.B2(n_382),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_367),
.A2(n_359),
.B(n_350),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_394),
.A2(n_355),
.B(n_358),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_406),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_344),
.Y(n_396)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_396),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_353),
.Y(n_397)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_397),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_374),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_368),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_380),
.B(n_338),
.C(n_359),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_321),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_398),
.B(n_381),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_395),
.Y(n_430)
);

FAx1_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_375),
.CI(n_371),
.CON(n_412),
.SN(n_412)
);

O2A1O1Ixp33_ASAP7_75t_L g434 ( 
.A1(n_412),
.A2(n_394),
.B(n_400),
.C(n_401),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_369),
.C(n_379),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_413),
.B(n_422),
.C(n_406),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_414),
.A2(n_415),
.B1(n_418),
.B2(n_419),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_387),
.A2(n_378),
.B1(n_383),
.B2(n_350),
.Y(n_415)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_416),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_390),
.A2(n_335),
.B1(n_342),
.B2(n_345),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_402),
.A2(n_355),
.B1(n_342),
.B2(n_345),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_336),
.C(n_361),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_430),
.Y(n_440)
);

BUFx24_ASAP7_75t_SL g425 ( 
.A(n_423),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_425),
.B(n_435),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_409),
.B(n_389),
.C(n_404),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_426),
.B(n_431),
.C(n_424),
.Y(n_438)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_419),
.Y(n_428)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_428),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_418),
.A2(n_390),
.B1(n_392),
.B2(n_400),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_429),
.A2(n_405),
.B1(n_407),
.B2(n_399),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_388),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g436 ( 
.A1(n_434),
.A2(n_412),
.B(n_415),
.C(n_410),
.D(n_401),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_421),
.Y(n_435)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_436),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_437),
.A2(n_442),
.B1(n_405),
.B2(n_429),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_438),
.A2(n_430),
.B(n_413),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_427),
.B(n_410),
.Y(n_441)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_441),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_434),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_409),
.C(n_411),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_443),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_432),
.A2(n_412),
.B(n_399),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_445),
.A2(n_432),
.B(n_433),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_447),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_441),
.B(n_408),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_448),
.B(n_450),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_445),
.A2(n_422),
.B(n_431),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_451),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_452),
.B(n_439),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_438),
.Y(n_460)
);

AOI322xp5_ASAP7_75t_L g456 ( 
.A1(n_448),
.A2(n_453),
.A3(n_449),
.B1(n_407),
.B2(n_436),
.C1(n_444),
.C2(n_348),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_456),
.B(n_458),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_443),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_462),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_455),
.B(n_440),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_457),
.B(n_440),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_463),
.B(n_461),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_460),
.B(n_459),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_466),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_465),
.A2(n_457),
.B(n_417),
.Y(n_467)
);

AOI322xp5_ASAP7_75t_L g469 ( 
.A1(n_467),
.A2(n_385),
.A3(n_333),
.B1(n_360),
.B2(n_363),
.C1(n_348),
.C2(n_370),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_469),
.B(n_366),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_470),
.B(n_468),
.Y(n_471)
);


endmodule