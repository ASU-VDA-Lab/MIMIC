module fake_jpeg_19389_n_168 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_168);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_11),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_4),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_7),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_4),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_33),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_6),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_69),
.Y(n_81)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_81),
.Y(n_88)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_83),
.Y(n_87)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_67),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_68),
.B1(n_76),
.B2(n_75),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_93),
.A2(n_57),
.B1(n_63),
.B2(n_77),
.Y(n_107)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_106),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_66),
.B1(n_80),
.B2(n_71),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_100),
.B1(n_62),
.B2(n_67),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_62),
.B1(n_49),
.B2(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_103),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_84),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_79),
.B1(n_49),
.B2(n_57),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_108),
.B1(n_90),
.B2(n_91),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_0),
.C(n_1),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_94),
.B1(n_96),
.B2(n_55),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_73),
.C(n_70),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_120),
.B(n_125),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_65),
.B1(n_60),
.B2(n_58),
.Y(n_128)
);

AO21x2_ASAP7_75t_L g112 ( 
.A1(n_104),
.A2(n_100),
.B(n_94),
.Y(n_112)
);

AO21x2_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_72),
.B(n_25),
.Y(n_132)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_127),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_54),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_123),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_74),
.B1(n_59),
.B2(n_64),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_118),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_99),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_123),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_54),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

NAND2x1_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_0),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_76),
.C(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_134),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_112),
.B1(n_26),
.B2(n_32),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_136),
.B(n_140),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_20),
.B(n_44),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_15),
.C(n_43),
.Y(n_146)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_142),
.B(n_145),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_149),
.B1(n_150),
.B2(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_148),
.Y(n_152)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_47),
.Y(n_148)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_135),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_12),
.C(n_39),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_143),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_156),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_148),
.Y(n_156)
);

OAI322xp33_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_152),
.A3(n_154),
.B1(n_151),
.B2(n_132),
.C1(n_149),
.C2(n_133),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_132),
.Y(n_160)
);

OAI21x1_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_133),
.B(n_128),
.Y(n_161)
);

OAI21x1_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_138),
.B(n_2),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_42),
.C(n_38),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_36),
.B(n_35),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_164),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_34),
.B1(n_16),
.B2(n_3),
.Y(n_166)
);

AO221x1_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.C(n_7),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_167),
.B(n_8),
.Y(n_168)
);


endmodule