module real_jpeg_25288_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_213;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_202;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx3_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_1),
.A2(n_69),
.B1(n_71),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_1),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_84),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_84),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_29),
.B1(n_41),
.B2(n_42),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_5),
.A2(n_69),
.B1(n_71),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_5),
.A2(n_41),
.B1(n_42),
.B2(n_133),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_133),
.Y(n_255)
);

INVx8_ASAP7_75t_SL g78 ( 
.A(n_6),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_7),
.A2(n_63),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_63),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_63),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_8),
.A2(n_33),
.B1(n_41),
.B2(n_42),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_11),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_12),
.B(n_71),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_12),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_12),
.B(n_80),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_12),
.B(n_42),
.C(n_55),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_12),
.A2(n_58),
.B1(n_59),
.B2(n_181),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_12),
.B(n_152),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_12),
.A2(n_41),
.B1(n_42),
.B2(n_181),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_12),
.B(n_28),
.C(n_46),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_12),
.A2(n_30),
.B(n_243),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_43),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_15),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_15),
.A2(n_41),
.B1(n_42),
.B2(n_68),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_68),
.Y(n_242)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_16),
.Y(n_191)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_16),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_114),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_20),
.B(n_114),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_113),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.C(n_65),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_25),
.A2(n_37),
.B1(n_38),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_25),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_26),
.A2(n_30),
.B1(n_100),
.B2(n_122),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_27),
.B(n_267),
.Y(n_266)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_31),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_30),
.A2(n_32),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_30),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_30),
.A2(n_157),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_30),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_30),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_35),
.A2(n_123),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_35),
.B(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_40),
.A2(n_48),
.B1(n_91),
.B2(n_125),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_42),
.B1(n_55),
.B2(n_56),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_42),
.B(n_250),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_44),
.A2(n_49),
.B1(n_51),
.B2(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_44),
.B(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_44),
.A2(n_51),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_48),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_48),
.A2(n_125),
.B(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_48),
.A2(n_174),
.B(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_48),
.B(n_181),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_51),
.B(n_175),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_52),
.B(n_65),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_64),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_54),
.B1(n_64),
.B2(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_53),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_53),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_53),
.A2(n_151),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_62),
.B(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_54),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_54),
.A2(n_128),
.B(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_59),
.B1(n_76),
.B2(n_77),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_69),
.A3(n_77),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g160 ( 
.A(n_59),
.B(n_76),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_59),
.B(n_206),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_73),
.B(n_81),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_74),
.B1(n_80),
.B2(n_132),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_70),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_70),
.Y(n_180)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_74),
.A2(n_82),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_108),
.B(n_111),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_79),
.A2(n_111),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_96),
.B2(n_97),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B(n_95),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_90),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_91),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_91),
.A2(n_231),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_105),
.B1(n_106),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_99),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_99),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_100),
.B(n_181),
.Y(n_267)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.C(n_119),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_118),
.Y(n_162)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_126),
.C(n_131),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_121),
.B(n_124),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_127),
.B1(n_131),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_150),
.B1(n_152),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_132),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_163),
.B(n_291),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_161),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_138),
.B(n_161),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.C(n_145),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_143),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_145),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.C(n_153),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_148),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_153),
.B(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_158),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_154),
.B(n_158),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_155),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

O2A1O1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_198),
.B(n_285),
.C(n_290),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_192),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_192),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_183),
.C(n_184),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_166),
.A2(n_167),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_176),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_172),
.C(n_176),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B(n_182),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_183),
.B(n_184),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.C(n_189),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_225),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_193),
.B(n_196),
.C(n_197),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_279),
.B(n_284),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_232),
.B(n_278),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_221),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_203),
.B(n_221),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_214),
.C(n_218),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_204),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_207),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_207),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B(n_212),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_211),
.A2(n_255),
.B(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_214),
.A2(n_218),
.B1(n_219),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_214),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_222),
.B(n_228),
.C(n_229),
.Y(n_283)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_272),
.B(n_277),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_251),
.B(n_271),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_245),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_245),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_242),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_249),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_247),
.B1(n_249),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_249),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_260),
.B(n_270),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_258),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_258),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_265),
.B(n_269),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_263),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_268),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_276),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_287),
.Y(n_290)
);


endmodule