module fake_aes_2144_n_1118 (n_117, n_219, n_44, n_133, n_149, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_16, n_13, n_198, n_169, n_193, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_270, n_246, n_153, n_61, n_259, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_1118);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
output n_1118;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1092;
wire n_1077;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_1059;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_1093;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_1056;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_1095;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_1074;
wire n_436;
wire n_588;
wire n_275;
wire n_1048;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_1087;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_476;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_1012;
wire n_1098;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_345;
wire n_360;
wire n_1090;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_286;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1024;
wire n_1016;
wire n_1078;
wire n_572;
wire n_1017;
wire n_324;
wire n_1097;
wire n_773;
wire n_847;
wire n_1094;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_279;
wire n_303;
wire n_1042;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_1081;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_880;
wire n_1101;
wire n_630;
wire n_511;
wire n_277;
wire n_1002;
wire n_467;
wire n_1072;
wire n_692;
wire n_865;
wire n_1064;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_274;
wire n_1018;
wire n_738;
wire n_979;
wire n_282;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_1063;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_1062;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_1091;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_950;
wire n_910;
wire n_460;
wire n_1046;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_928;
wire n_938;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_1076;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_805;
wire n_729;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_1061;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_1106;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_1113;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_302;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_1041;
wire n_542;
wire n_1080;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_1099;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_1065;
wire n_549;
wire n_622;
wire n_875;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_1047;
wire n_320;
wire n_768;
wire n_1107;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_1089;
wire n_1058;
wire n_370;
wire n_1050;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_1049;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_970;
wire n_822;
wire n_984;
wire n_390;
wire n_682;
wire n_1082;
wire n_1052;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_1066;
wire n_539;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_1116;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_1114;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_1071;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_1079;
wire n_409;
wire n_315;
wire n_363;
wire n_733;
wire n_861;
wire n_899;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_1057;
wire n_681;
wire n_435;
wire n_577;
wire n_1068;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_1051;
wire n_615;
wire n_1029;
wire n_472;
wire n_1100;
wire n_1088;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_1060;
wire n_429;
wire n_488;
wire n_1037;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_1110;
wire n_325;
wire n_1102;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_1069;
wire n_811;
wire n_1039;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_1054;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_1044;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_947;
wire n_620;
wire n_1043;
wire n_924;
wire n_841;
wire n_912;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_1096;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_1117;
wire n_1040;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_1053;
wire n_774;
wire n_867;
wire n_1070;
wire n_377;
wire n_510;
wire n_343;
wire n_1075;
wire n_1112;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_1084;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_1083;
wire n_356;
wire n_281;
wire n_1038;
wire n_341;
wire n_470;
wire n_600;
wire n_1103;
wire n_1085;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_1073;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_1111;
wire n_1045;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1115;
wire n_521;
wire n_695;
wire n_625;
wire n_650;
wire n_469;
wire n_1104;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_1067;
wire n_736;
wire n_1108;
wire n_287;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_1105;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_1086;
wire n_385;
wire n_992;
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_62), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_263), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g274 ( .A(n_256), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_43), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_261), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_140), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_120), .Y(n_278) );
CKINVDCx5p33_ASAP7_75t_R g279 ( .A(n_225), .Y(n_279) );
CKINVDCx5p33_ASAP7_75t_R g280 ( .A(n_190), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_161), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_145), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_126), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_259), .Y(n_285) );
BUFx2_ASAP7_75t_SL g286 ( .A(n_223), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_49), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_176), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_141), .B(n_146), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_211), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_69), .Y(n_292) );
CKINVDCx5p33_ASAP7_75t_R g293 ( .A(n_14), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_240), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_124), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_43), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_253), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_64), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_269), .Y(n_299) );
CKINVDCx5p33_ASAP7_75t_R g300 ( .A(n_266), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_191), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_137), .Y(n_303) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_46), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_0), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_251), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_154), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_94), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g310 ( .A(n_212), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_252), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_237), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_38), .Y(n_313) );
INVxp67_ASAP7_75t_L g314 ( .A(n_164), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_245), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_116), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_167), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_175), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_52), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_136), .Y(n_320) );
INVxp33_ASAP7_75t_SL g321 ( .A(n_108), .Y(n_321) );
INVx3_ASAP7_75t_L g322 ( .A(n_9), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_242), .Y(n_323) );
BUFx6f_ASAP7_75t_L g324 ( .A(n_118), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_200), .Y(n_325) );
BUFx5_ASAP7_75t_L g326 ( .A(n_94), .Y(n_326) );
XNOR2x1_ASAP7_75t_L g327 ( .A(n_55), .B(n_119), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_149), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_192), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_155), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_160), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_180), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_15), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_219), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_93), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_134), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_71), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_271), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_177), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_68), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_202), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_131), .Y(n_343) );
CKINVDCx14_ASAP7_75t_R g344 ( .A(n_125), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_203), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_8), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_23), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_217), .Y(n_348) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_125), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_40), .Y(n_350) );
INVxp33_ASAP7_75t_SL g351 ( .A(n_61), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_89), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_132), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_67), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_59), .Y(n_355) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_255), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_186), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_63), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_166), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_229), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_57), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_6), .Y(n_362) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_81), .Y(n_363) );
BUFx6f_ASAP7_75t_L g364 ( .A(n_3), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_230), .Y(n_365) );
BUFx3_ASAP7_75t_L g366 ( .A(n_29), .Y(n_366) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_2), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_218), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_174), .Y(n_369) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_195), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_221), .B(n_130), .Y(n_371) );
INVx1_ASAP7_75t_SL g372 ( .A(n_183), .Y(n_372) );
CKINVDCx16_ASAP7_75t_R g373 ( .A(n_224), .Y(n_373) );
CKINVDCx5p33_ASAP7_75t_R g374 ( .A(n_246), .Y(n_374) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_171), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_194), .Y(n_376) );
BUFx10_ASAP7_75t_L g377 ( .A(n_241), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_188), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_179), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_185), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_198), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_234), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_222), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_81), .Y(n_384) );
CKINVDCx5p33_ASAP7_75t_R g385 ( .A(n_126), .Y(n_385) );
NOR2xp67_ASAP7_75t_L g386 ( .A(n_143), .B(n_8), .Y(n_386) );
BUFx5_ASAP7_75t_L g387 ( .A(n_216), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_46), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_163), .B(n_168), .Y(n_389) );
BUFx5_ASAP7_75t_L g390 ( .A(n_231), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_110), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_184), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_158), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_189), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_97), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_148), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_66), .Y(n_397) );
INVx2_ASAP7_75t_SL g398 ( .A(n_96), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_182), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_387), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_326), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_305), .A2(n_128), .B(n_127), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_387), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_319), .B(n_0), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_387), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_387), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_387), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_326), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_344), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_309), .B(n_4), .Y(n_412) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_320), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_309), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_322), .B(n_5), .Y(n_415) );
BUFx12f_ASAP7_75t_L g416 ( .A(n_377), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_344), .A2(n_10), .B1(n_7), .B2(n_9), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_322), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_387), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_369), .B(n_7), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_390), .Y(n_422) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_321), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_423) );
AND2x6_ASAP7_75t_L g424 ( .A(n_389), .B(n_129), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_326), .Y(n_425) );
AND2x2_ASAP7_75t_SL g426 ( .A(n_301), .B(n_270), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_326), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_328), .B(n_12), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_370), .Y(n_430) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_320), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_320), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_326), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_321), .A2(n_17), .B1(n_15), .B2(n_16), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_320), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_400), .Y(n_436) );
INVx5_ASAP7_75t_L g437 ( .A(n_424), .Y(n_437) );
BUFx3_ASAP7_75t_L g438 ( .A(n_424), .Y(n_438) );
INVx3_ASAP7_75t_L g439 ( .A(n_420), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_400), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_426), .A2(n_351), .B1(n_367), .B2(n_317), .Y(n_441) );
AND2x4_ASAP7_75t_L g442 ( .A(n_414), .B(n_313), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g443 ( .A(n_416), .B(n_373), .Y(n_443) );
NAND3xp33_ASAP7_75t_L g444 ( .A(n_401), .B(n_285), .C(n_281), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_401), .B(n_290), .C(n_288), .Y(n_445) );
OR2x6_ASAP7_75t_L g446 ( .A(n_411), .B(n_286), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_403), .Y(n_448) );
INVx4_ASAP7_75t_L g449 ( .A(n_424), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_414), .B(n_396), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_430), .Y(n_451) );
OR2x6_ASAP7_75t_L g452 ( .A(n_417), .B(n_398), .Y(n_452) );
NAND2xp33_ASAP7_75t_L g453 ( .A(n_424), .B(n_390), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_420), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_405), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_414), .B(n_298), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_405), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_420), .Y(n_458) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_405), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_407), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_407), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_407), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_408), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_410), .Y(n_465) );
INVx4_ASAP7_75t_L g466 ( .A(n_424), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_408), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_408), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_459), .B(n_426), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_451), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_454), .B(n_424), .Y(n_472) );
NOR2xp33_ASAP7_75t_SL g473 ( .A(n_449), .B(n_323), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_442), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_459), .B(n_412), .Y(n_475) );
OAI22xp5_ASAP7_75t_L g476 ( .A1(n_441), .A2(n_434), .B1(n_423), .B2(n_365), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_450), .B(n_429), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_456), .B(n_418), .Y(n_478) );
BUFx8_ASAP7_75t_L g479 ( .A(n_451), .Y(n_479) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_439), .B(n_424), .Y(n_480) );
AND2x6_ASAP7_75t_SL g481 ( .A(n_446), .B(n_404), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_449), .B(n_323), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_454), .B(n_415), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_442), .B(n_410), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_442), .B(n_410), .Y(n_485) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_439), .A2(n_409), .B(n_425), .C(n_406), .Y(n_486) );
INVx2_ASAP7_75t_SL g487 ( .A(n_443), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_439), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g489 ( .A(n_453), .B(n_466), .C(n_449), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_439), .B(n_294), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_458), .A2(n_406), .B1(n_427), .B2(n_425), .Y(n_491) );
AND2x4_ASAP7_75t_L g492 ( .A(n_458), .B(n_466), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_465), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_437), .B(n_314), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_436), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_440), .B(n_297), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_437), .B(n_342), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_466), .A2(n_433), .B(n_421), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_447), .B(n_342), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
INVx8_ASAP7_75t_L g502 ( .A(n_446), .Y(n_502) );
OR2x2_ASAP7_75t_L g503 ( .A(n_452), .B(n_327), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_448), .Y(n_504) );
AND2x4_ASAP7_75t_L g505 ( .A(n_446), .B(n_402), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_446), .A2(n_349), .B1(n_362), .B2(n_304), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_452), .B(n_402), .Y(n_507) );
OR2x6_ASAP7_75t_L g508 ( .A(n_452), .B(n_327), .Y(n_508) );
OR2x6_ASAP7_75t_L g509 ( .A(n_452), .B(n_275), .Y(n_509) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_438), .A2(n_444), .B1(n_445), .B2(n_455), .Y(n_510) );
NOR2x1p5_ASAP7_75t_L g511 ( .A(n_438), .B(n_397), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_455), .B(n_419), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_457), .B(n_273), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_457), .B(n_272), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_461), .B(n_274), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_461), .B(n_366), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_464), .B(n_276), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_468), .B(n_279), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_468), .B(n_345), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_460), .A2(n_362), .B1(n_349), .B2(n_296), .Y(n_521) );
NOR3xp33_ASAP7_75t_L g522 ( .A(n_462), .B(n_293), .C(n_278), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_462), .B(n_280), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_463), .B(n_275), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_467), .B(n_292), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_469), .B(n_419), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_469), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_487), .B(n_358), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_514), .B(n_361), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_480), .A2(n_422), .B(n_421), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_472), .A2(n_428), .B(n_422), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_472), .A2(n_428), .B(n_422), .Y(n_532) );
AO32x2_ASAP7_75t_L g533 ( .A1(n_476), .A2(n_390), .A3(n_386), .B1(n_431), .B2(n_413), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_499), .A2(n_428), .B(n_291), .Y(n_534) );
BUFx3_ASAP7_75t_L g535 ( .A(n_479), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_509), .A2(n_497), .B1(n_470), .B2(n_502), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_507), .A2(n_334), .B1(n_341), .B2(n_306), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_483), .A2(n_303), .B(n_299), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_488), .A2(n_308), .B(n_307), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_479), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_516), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_489), .A2(n_312), .B(n_311), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_502), .A2(n_347), .B1(n_350), .B2(n_346), .Y(n_543) );
INVx6_ASAP7_75t_L g544 ( .A(n_481), .Y(n_544) );
BUFx6f_ASAP7_75t_L g545 ( .A(n_492), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_492), .A2(n_318), .B(n_315), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_478), .A2(n_329), .B(n_325), .Y(n_547) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_486), .A2(n_331), .B(n_330), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_490), .A2(n_333), .B(n_332), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_473), .A2(n_354), .B1(n_355), .B2(n_352), .Y(n_550) );
OR2x6_ASAP7_75t_L g551 ( .A(n_502), .B(n_283), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_484), .A2(n_339), .B(n_337), .Y(n_552) );
BUFx3_ASAP7_75t_L g553 ( .A(n_516), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_485), .A2(n_343), .B(n_340), .Y(n_554) );
O2A1O1Ixp5_ASAP7_75t_L g555 ( .A1(n_505), .A2(n_371), .B(n_289), .C(n_282), .Y(n_555) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_506), .A2(n_508), .B1(n_476), .B2(n_503), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_513), .A2(n_353), .B(n_348), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_482), .B(n_300), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_525), .Y(n_559) );
AO22x1_ASAP7_75t_L g560 ( .A1(n_521), .A2(n_388), .B1(n_391), .B2(n_385), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_515), .A2(n_359), .B(n_357), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_525), .B(n_295), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g563 ( .A1(n_501), .A2(n_504), .B1(n_507), .B2(n_475), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_524), .Y(n_564) );
AOI21x1_ASAP7_75t_L g565 ( .A1(n_526), .A2(n_379), .B(n_368), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_511), .B(n_316), .Y(n_566) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_524), .A2(n_338), .B1(n_384), .B2(n_336), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_522), .B(n_338), .Y(n_568) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_524), .A2(n_384), .B1(n_324), .B2(n_363), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_517), .B(n_372), .Y(n_570) );
AND2x4_ASAP7_75t_L g571 ( .A(n_519), .B(n_382), .Y(n_571) );
INVx4_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_491), .A2(n_324), .B1(n_363), .B2(n_287), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_512), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_496), .B(n_310), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_518), .A2(n_393), .B(n_392), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_500), .B(n_335), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_520), .A2(n_399), .B(n_282), .C(n_284), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_523), .B(n_360), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_495), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g582 ( .A1(n_494), .A2(n_284), .B(n_302), .C(n_277), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_510), .A2(n_287), .B1(n_363), .B2(n_324), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_493), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_498), .B(n_374), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_527), .A2(n_324), .B1(n_363), .B2(n_287), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_480), .A2(n_378), .B(n_371), .Y(n_587) );
INVx1_ASAP7_75t_SL g588 ( .A(n_471), .Y(n_588) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_492), .Y(n_589) );
INVx3_ASAP7_75t_L g590 ( .A(n_492), .Y(n_590) );
AO21x1_ASAP7_75t_L g591 ( .A1(n_505), .A2(n_390), .B(n_413), .Y(n_591) );
INVx3_ASAP7_75t_SL g592 ( .A(n_509), .Y(n_592) );
AOI21xp5_ASAP7_75t_L g593 ( .A1(n_480), .A2(n_376), .B(n_375), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_480), .A2(n_381), .B(n_380), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_477), .B(n_383), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g596 ( .A1(n_509), .A2(n_364), .B1(n_395), .B2(n_356), .Y(n_596) );
BUFx3_ASAP7_75t_L g597 ( .A(n_479), .Y(n_597) );
BUFx12f_ASAP7_75t_L g598 ( .A(n_479), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_509), .A2(n_364), .B1(n_395), .B2(n_394), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_474), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_477), .B(n_395), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_509), .A2(n_356), .B1(n_432), .B2(n_431), .Y(n_602) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_487), .B(n_17), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_487), .B(n_18), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_509), .A2(n_435), .B1(n_432), .B2(n_21), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_473), .B(n_432), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_474), .Y(n_607) );
BUFx3_ASAP7_75t_L g608 ( .A(n_479), .Y(n_608) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_480), .A2(n_135), .B(n_133), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_509), .A2(n_435), .B1(n_21), .B2(n_19), .Y(n_610) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_509), .A2(n_435), .B1(n_23), .B2(n_20), .Y(n_611) );
AND2x4_ASAP7_75t_L g612 ( .A(n_509), .B(n_22), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_521), .B(n_22), .Y(n_613) );
AO31x2_ASAP7_75t_L g614 ( .A1(n_591), .A2(n_26), .A3(n_24), .B(n_25), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_601), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_532), .A2(n_139), .B(n_138), .Y(n_616) );
INVx8_ASAP7_75t_L g617 ( .A(n_540), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_535), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_575), .B(n_26), .Y(n_619) );
AO31x2_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_29), .A3(n_27), .B(n_28), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_597), .Y(n_621) );
AO21x2_ASAP7_75t_L g622 ( .A1(n_565), .A2(n_144), .B(n_142), .Y(n_622) );
AO31x2_ASAP7_75t_L g623 ( .A1(n_583), .A2(n_31), .A3(n_28), .B(n_30), .Y(n_623) );
BUFx3_ASAP7_75t_L g624 ( .A(n_608), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_530), .A2(n_150), .B(n_147), .Y(n_625) );
AO21x2_ASAP7_75t_L g626 ( .A1(n_563), .A2(n_152), .B(n_151), .Y(n_626) );
AO31x2_ASAP7_75t_L g627 ( .A1(n_582), .A2(n_34), .A3(n_32), .B(n_33), .Y(n_627) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_576), .A2(n_156), .B(n_153), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_562), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_578), .A2(n_159), .B(n_157), .Y(n_630) );
BUFx5_ASAP7_75t_L g631 ( .A(n_581), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_555), .A2(n_34), .B(n_32), .C(n_33), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_592), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_549), .A2(n_165), .B(n_162), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_560), .B(n_35), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_541), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_559), .Y(n_637) );
OA21x2_ASAP7_75t_L g638 ( .A1(n_609), .A2(n_170), .B(n_169), .Y(n_638) );
BUFx10_ASAP7_75t_L g639 ( .A(n_612), .Y(n_639) );
AO31x2_ASAP7_75t_L g640 ( .A1(n_537), .A2(n_39), .A3(n_36), .B(n_37), .Y(n_640) );
A2O1A1Ixp33_ASAP7_75t_L g641 ( .A1(n_557), .A2(n_561), .B(n_577), .C(n_579), .Y(n_641) );
BUFx2_ASAP7_75t_L g642 ( .A(n_612), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_538), .A2(n_44), .B(n_41), .C(n_42), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_563), .A2(n_44), .B1(n_41), .B2(n_42), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_595), .A2(n_173), .B(n_172), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_600), .Y(n_646) );
AO31x2_ASAP7_75t_L g647 ( .A1(n_596), .A2(n_48), .A3(n_45), .B(n_47), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_534), .A2(n_181), .B(n_178), .Y(n_648) );
AND2x4_ASAP7_75t_L g649 ( .A(n_590), .B(n_48), .Y(n_649) );
AO31x2_ASAP7_75t_L g650 ( .A1(n_567), .A2(n_50), .A3(n_51), .B(n_52), .Y(n_650) );
OAI21xp5_ASAP7_75t_SL g651 ( .A1(n_550), .A2(n_53), .B(n_54), .Y(n_651) );
AO31x2_ASAP7_75t_L g652 ( .A1(n_573), .A2(n_53), .A3(n_54), .B(n_55), .Y(n_652) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_564), .B(n_56), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_547), .A2(n_57), .B(n_58), .C(n_60), .Y(n_654) );
BUFx8_ASAP7_75t_L g655 ( .A(n_533), .Y(n_655) );
BUFx2_ASAP7_75t_SL g656 ( .A(n_572), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_607), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_552), .A2(n_196), .B(n_193), .Y(n_658) );
O2A1O1Ixp33_ASAP7_75t_SL g659 ( .A1(n_606), .A2(n_201), .B(n_267), .C(n_264), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_613), .Y(n_660) );
AOI21xp5_ASAP7_75t_L g661 ( .A1(n_554), .A2(n_199), .B(n_197), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_551), .B(n_65), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_551), .B(n_66), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_551), .B(n_70), .Y(n_664) );
AO31x2_ASAP7_75t_L g665 ( .A1(n_605), .A2(n_72), .A3(n_73), .B(n_74), .Y(n_665) );
OAI22xp33_ASAP7_75t_L g666 ( .A1(n_550), .A2(n_72), .B1(n_73), .B2(n_74), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_564), .A2(n_75), .B1(n_76), .B2(n_77), .Y(n_667) );
BUFx2_ASAP7_75t_L g668 ( .A(n_553), .Y(n_668) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_587), .A2(n_209), .B(n_262), .Y(n_669) );
NAND2x1p5_ASAP7_75t_L g670 ( .A(n_545), .B(n_78), .Y(n_670) );
AO31x2_ASAP7_75t_L g671 ( .A1(n_611), .A2(n_78), .A3(n_79), .B(n_80), .Y(n_671) );
AOI21xp5_ASAP7_75t_L g672 ( .A1(n_546), .A2(n_208), .B(n_260), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_543), .A2(n_79), .B(n_80), .C(n_82), .Y(n_673) );
AO21x1_ASAP7_75t_L g674 ( .A1(n_548), .A2(n_210), .B(n_258), .Y(n_674) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_580), .A2(n_207), .B(n_257), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_568), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_536), .A2(n_83), .B1(n_84), .B2(n_85), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_545), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_593), .A2(n_213), .B(n_254), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_568), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_566), .B(n_86), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_544), .A2(n_528), .B1(n_604), .B2(n_603), .Y(n_682) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_594), .A2(n_205), .B(n_249), .Y(n_683) );
BUFx2_ASAP7_75t_L g684 ( .A(n_545), .Y(n_684) );
AO31x2_ASAP7_75t_L g685 ( .A1(n_602), .A2(n_86), .A3(n_87), .B(n_88), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_589), .Y(n_686) );
AO21x2_ASAP7_75t_L g687 ( .A1(n_548), .A2(n_206), .B(n_248), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_542), .A2(n_87), .B(n_88), .C(n_89), .Y(n_688) );
OAI21xp5_ASAP7_75t_L g689 ( .A1(n_539), .A2(n_214), .B(n_247), .Y(n_689) );
BUFx2_ASAP7_75t_L g690 ( .A(n_589), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_571), .A2(n_90), .B1(n_91), .B2(n_92), .Y(n_691) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_571), .A2(n_90), .B1(n_92), .B2(n_93), .Y(n_692) );
BUFx3_ASAP7_75t_L g693 ( .A(n_589), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_529), .A2(n_95), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_694) );
AND2x4_ASAP7_75t_L g695 ( .A(n_584), .B(n_95), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_569), .Y(n_696) );
AOI221x1_ASAP7_75t_L g697 ( .A1(n_586), .A2(n_99), .B1(n_100), .B2(n_101), .C(n_102), .Y(n_697) );
AOI21xp5_ASAP7_75t_L g698 ( .A1(n_558), .A2(n_220), .B(n_244), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_585), .A2(n_215), .B(n_243), .Y(n_699) );
AO31x2_ASAP7_75t_L g700 ( .A1(n_586), .A2(n_101), .A3(n_102), .B(n_103), .Y(n_700) );
INVx5_ASAP7_75t_L g701 ( .A(n_533), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_570), .B(n_104), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_599), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_533), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_610), .Y(n_705) );
OR2x2_ASAP7_75t_L g706 ( .A(n_588), .B(n_109), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_574), .B(n_109), .Y(n_707) );
BUFx2_ASAP7_75t_L g708 ( .A(n_588), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_556), .A2(n_111), .B1(n_112), .B2(n_113), .Y(n_709) );
BUFx8_ASAP7_75t_L g710 ( .A(n_598), .Y(n_710) );
INVx1_ASAP7_75t_SL g711 ( .A(n_588), .Y(n_711) );
CKINVDCx11_ASAP7_75t_R g712 ( .A(n_598), .Y(n_712) );
INVx2_ASAP7_75t_L g713 ( .A(n_574), .Y(n_713) );
INVxp67_ASAP7_75t_L g714 ( .A(n_588), .Y(n_714) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_574), .A2(n_113), .B1(n_114), .B2(n_115), .Y(n_715) );
AO31x2_ASAP7_75t_L g716 ( .A1(n_591), .A2(n_116), .A3(n_117), .B(n_118), .Y(n_716) );
BUFx2_ASAP7_75t_L g717 ( .A(n_588), .Y(n_717) );
AOI21xp5_ASAP7_75t_SL g718 ( .A1(n_572), .A2(n_268), .B(n_228), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g719 ( .A1(n_531), .A2(n_226), .B(n_238), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_601), .Y(n_720) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_545), .Y(n_721) );
INVx1_ASAP7_75t_SL g722 ( .A(n_588), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_574), .B(n_121), .Y(n_723) );
AND2x4_ASAP7_75t_L g724 ( .A(n_713), .B(n_642), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_722), .B(n_122), .Y(n_725) );
NAND2x1p5_ASAP7_75t_L g726 ( .A(n_664), .B(n_123), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_717), .B(n_123), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_714), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_660), .B(n_124), .Y(n_729) );
INVxp67_ASAP7_75t_SL g730 ( .A(n_655), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_646), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g732 ( .A1(n_617), .A2(n_239), .B(n_232), .Y(n_732) );
OAI22x1_ASAP7_75t_L g733 ( .A1(n_664), .A2(n_204), .B1(n_233), .B2(n_236), .Y(n_733) );
OAI21xp5_ASAP7_75t_L g734 ( .A1(n_632), .A2(n_705), .B(n_619), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_657), .Y(n_735) );
AO21x2_ASAP7_75t_L g736 ( .A1(n_616), .A2(n_719), .B(n_648), .Y(n_736) );
AND2x4_ASAP7_75t_L g737 ( .A(n_676), .B(n_680), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_710), .Y(n_738) );
NAND2x1p5_ASAP7_75t_L g739 ( .A(n_695), .B(n_649), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_629), .B(n_637), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_723), .B(n_707), .Y(n_741) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_669), .A2(n_696), .B(n_702), .Y(n_742) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_695), .B(n_649), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_638), .A2(n_630), .B(n_628), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_710), .Y(n_745) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_712), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g747 ( .A1(n_679), .A2(n_683), .B(n_645), .Y(n_747) );
AO31x2_ASAP7_75t_L g748 ( .A1(n_697), .A2(n_644), .A3(n_688), .B(n_654), .Y(n_748) );
AO21x2_ASAP7_75t_L g749 ( .A1(n_622), .A2(n_689), .B(n_626), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_706), .Y(n_750) );
CKINVDCx11_ASAP7_75t_R g751 ( .A(n_618), .Y(n_751) );
AO21x2_ASAP7_75t_L g752 ( .A1(n_687), .A2(n_699), .B(n_625), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_636), .B(n_631), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_659), .A2(n_661), .B(n_658), .Y(n_754) );
BUFx3_ASAP7_75t_L g755 ( .A(n_617), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_631), .B(n_682), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_631), .B(n_709), .Y(n_757) );
AO31x2_ASAP7_75t_L g758 ( .A1(n_677), .A2(n_643), .A3(n_715), .B(n_634), .Y(n_758) );
OA21x2_ASAP7_75t_L g759 ( .A1(n_672), .A2(n_698), .B(n_675), .Y(n_759) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_701), .A2(n_653), .B1(n_670), .B2(n_694), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_678), .B(n_686), .Y(n_761) );
INVx1_ASAP7_75t_SL g762 ( .A(n_639), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_662), .B(n_663), .Y(n_763) );
AO21x2_ASAP7_75t_L g764 ( .A1(n_703), .A2(n_635), .B(n_666), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_640), .Y(n_765) );
AO31x2_ASAP7_75t_L g766 ( .A1(n_667), .A2(n_692), .A3(n_691), .B(n_655), .Y(n_766) );
OR2x2_ASAP7_75t_L g767 ( .A(n_624), .B(n_633), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_684), .B(n_690), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g769 ( .A1(n_673), .A2(n_718), .B(n_681), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_621), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_640), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_640), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_668), .B(n_693), .Y(n_773) );
OR2x6_ASAP7_75t_L g774 ( .A(n_656), .B(n_671), .Y(n_774) );
AO31x2_ASAP7_75t_L g775 ( .A1(n_614), .A2(n_716), .A3(n_627), .B(n_623), .Y(n_775) );
OAI21x1_ASAP7_75t_L g776 ( .A1(n_716), .A2(n_614), .B(n_627), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_650), .Y(n_777) );
AO31x2_ASAP7_75t_L g778 ( .A1(n_614), .A2(n_716), .A3(n_627), .B(n_623), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_620), .A2(n_623), .B(n_652), .Y(n_779) );
INVx4_ASAP7_75t_L g780 ( .A(n_647), .Y(n_780) );
OR2x6_ASAP7_75t_L g781 ( .A(n_671), .B(n_647), .Y(n_781) );
INVx2_ASAP7_75t_SL g782 ( .A(n_671), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_650), .B(n_665), .Y(n_783) );
AOI21x1_ASAP7_75t_L g784 ( .A1(n_652), .A2(n_665), .B(n_685), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_665), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g786 ( .A(n_700), .B(n_503), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_708), .B(n_717), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_713), .B(n_574), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_713), .Y(n_789) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_708), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_632), .A2(n_555), .B(n_641), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_713), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_713), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_713), .Y(n_794) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_708), .Y(n_795) );
OAI21xp5_ASAP7_75t_L g796 ( .A1(n_632), .A2(n_555), .B(n_641), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_713), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_713), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_713), .B(n_574), .Y(n_799) );
AO31x2_ASAP7_75t_L g800 ( .A1(n_704), .A2(n_674), .A3(n_591), .B(n_583), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_713), .B(n_574), .Y(n_801) );
INVx3_ASAP7_75t_L g802 ( .A(n_721), .Y(n_802) );
INVx1_ASAP7_75t_SL g803 ( .A(n_711), .Y(n_803) );
AO21x2_ASAP7_75t_L g804 ( .A1(n_704), .A2(n_632), .B(n_591), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_713), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_713), .B(n_574), .Y(n_806) );
INVx6_ASAP7_75t_L g807 ( .A(n_710), .Y(n_807) );
AO31x2_ASAP7_75t_L g808 ( .A1(n_704), .A2(n_674), .A3(n_591), .B(n_583), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_615), .A2(n_720), .B(n_641), .Y(n_809) );
AO21x2_ASAP7_75t_L g810 ( .A1(n_704), .A2(n_632), .B(n_591), .Y(n_810) );
OAI21x1_ASAP7_75t_SL g811 ( .A1(n_651), .A2(n_563), .B(n_572), .Y(n_811) );
BUFx3_ASAP7_75t_L g812 ( .A(n_710), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_704), .A2(n_632), .B(n_591), .Y(n_813) );
AO31x2_ASAP7_75t_L g814 ( .A1(n_704), .A2(n_674), .A3(n_591), .B(n_583), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g815 ( .A(n_714), .B(n_598), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_713), .B(n_574), .Y(n_816) );
AO21x2_ASAP7_75t_L g817 ( .A1(n_704), .A2(n_632), .B(n_591), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_713), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_785), .Y(n_819) );
AO21x1_ASAP7_75t_SL g820 ( .A1(n_756), .A2(n_753), .B(n_757), .Y(n_820) );
NOR2xp33_ASAP7_75t_SL g821 ( .A(n_738), .B(n_745), .Y(n_821) );
OR2x6_ASAP7_75t_L g822 ( .A(n_739), .B(n_743), .Y(n_822) );
AO21x2_ASAP7_75t_L g823 ( .A1(n_779), .A2(n_783), .B(n_784), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_731), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_735), .Y(n_825) );
BUFx3_ASAP7_75t_L g826 ( .A(n_812), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_786), .B(n_740), .Y(n_827) );
AND2x2_ASAP7_75t_L g828 ( .A(n_799), .B(n_793), .Y(n_828) );
INVx1_ASAP7_75t_L g829 ( .A(n_765), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_771), .Y(n_830) );
INVx1_ASAP7_75t_L g831 ( .A(n_772), .Y(n_831) );
OR2x6_ASAP7_75t_L g832 ( .A(n_743), .B(n_726), .Y(n_832) );
BUFx2_ASAP7_75t_L g833 ( .A(n_774), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_790), .Y(n_834) );
INVx1_ASAP7_75t_L g835 ( .A(n_789), .Y(n_835) );
OR2x2_ASAP7_75t_L g836 ( .A(n_730), .B(n_790), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_730), .B(n_788), .Y(n_837) );
AO21x2_ASAP7_75t_L g838 ( .A1(n_779), .A2(n_783), .B(n_776), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_777), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_782), .Y(n_840) );
BUFx3_ASAP7_75t_L g841 ( .A(n_807), .Y(n_841) );
AND2x2_ASAP7_75t_L g842 ( .A(n_805), .B(n_792), .Y(n_842) );
INVx4_ASAP7_75t_L g843 ( .A(n_726), .Y(n_843) );
AND2x2_ASAP7_75t_L g844 ( .A(n_794), .B(n_818), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_797), .B(n_798), .Y(n_845) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_728), .Y(n_846) );
BUFx2_ASAP7_75t_L g847 ( .A(n_774), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_788), .B(n_801), .Y(n_848) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_728), .Y(n_849) );
INVx1_ASAP7_75t_SL g850 ( .A(n_751), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_801), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_806), .B(n_816), .Y(n_852) );
OR2x6_ASAP7_75t_L g853 ( .A(n_811), .B(n_774), .Y(n_853) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_787), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_763), .B(n_781), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_727), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_750), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_781), .B(n_775), .Y(n_858) );
AO21x2_ASAP7_75t_L g859 ( .A1(n_791), .A2(n_796), .B(n_744), .Y(n_859) );
OR2x6_ASAP7_75t_L g860 ( .A(n_756), .B(n_733), .Y(n_860) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_795), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_775), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_781), .B(n_778), .Y(n_863) );
BUFx3_ASAP7_75t_L g864 ( .A(n_807), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_780), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g866 ( .A(n_807), .Y(n_866) );
INVx2_ASAP7_75t_SL g867 ( .A(n_767), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_780), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_753), .Y(n_869) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_791), .A2(n_796), .B(n_742), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_803), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_724), .B(n_734), .Y(n_872) );
BUFx12f_ASAP7_75t_L g873 ( .A(n_746), .Y(n_873) );
OR2x2_ASAP7_75t_L g874 ( .A(n_803), .B(n_768), .Y(n_874) );
AND2x2_ASAP7_75t_L g875 ( .A(n_724), .B(n_737), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_729), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_725), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_809), .Y(n_878) );
INVx2_ASAP7_75t_SL g879 ( .A(n_773), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_741), .B(n_766), .Y(n_880) );
AND2x2_ASAP7_75t_L g881 ( .A(n_766), .B(n_761), .Y(n_881) );
BUFx3_ASAP7_75t_L g882 ( .A(n_755), .Y(n_882) );
OR2x6_ASAP7_75t_L g883 ( .A(n_760), .B(n_757), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_768), .Y(n_884) );
BUFx3_ASAP7_75t_L g885 ( .A(n_802), .Y(n_885) );
AND2x4_ASAP7_75t_L g886 ( .A(n_802), .B(n_766), .Y(n_886) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_815), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_764), .A2(n_760), .B1(n_769), .B2(n_762), .Y(n_888) );
OR2x6_ASAP7_75t_L g889 ( .A(n_770), .B(n_754), .Y(n_889) );
AND2x2_ASAP7_75t_L g890 ( .A(n_880), .B(n_817), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_819), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_848), .B(n_762), .Y(n_892) );
AND2x2_ASAP7_75t_L g893 ( .A(n_880), .B(n_817), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_881), .B(n_804), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_848), .B(n_852), .Y(n_895) );
NOR2x1p5_ASAP7_75t_L g896 ( .A(n_866), .B(n_732), .Y(n_896) );
AND2x2_ASAP7_75t_L g897 ( .A(n_881), .B(n_804), .Y(n_897) );
AND2x2_ASAP7_75t_L g898 ( .A(n_855), .B(n_810), .Y(n_898) );
INVxp67_ASAP7_75t_SL g899 ( .A(n_837), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_837), .B(n_748), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_855), .B(n_810), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_819), .Y(n_902) );
AND2x2_ASAP7_75t_L g903 ( .A(n_858), .B(n_813), .Y(n_903) );
BUFx2_ASAP7_75t_L g904 ( .A(n_833), .Y(n_904) );
OR2x2_ASAP7_75t_L g905 ( .A(n_827), .B(n_748), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_839), .Y(n_906) );
OR2x2_ASAP7_75t_L g907 ( .A(n_836), .B(n_748), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_886), .B(n_749), .Y(n_908) );
INVxp67_ASAP7_75t_L g909 ( .A(n_867), .Y(n_909) );
INVx3_ASAP7_75t_L g910 ( .A(n_843), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_852), .B(n_758), .Y(n_911) );
NAND2xp5_ASAP7_75t_SL g912 ( .A(n_843), .B(n_747), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_829), .Y(n_913) );
BUFx2_ASAP7_75t_L g914 ( .A(n_833), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_829), .Y(n_915) );
OR2x2_ASAP7_75t_L g916 ( .A(n_836), .B(n_758), .Y(n_916) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_851), .Y(n_917) );
AND2x2_ASAP7_75t_L g918 ( .A(n_863), .B(n_758), .Y(n_918) );
HB1xp67_ASAP7_75t_L g919 ( .A(n_884), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_830), .Y(n_920) );
AND2x2_ASAP7_75t_L g921 ( .A(n_863), .B(n_869), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_846), .Y(n_922) );
INVxp67_ASAP7_75t_L g923 ( .A(n_867), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_831), .Y(n_924) );
HB1xp67_ASAP7_75t_L g925 ( .A(n_849), .Y(n_925) );
OR2x2_ASAP7_75t_L g926 ( .A(n_874), .B(n_814), .Y(n_926) );
AND2x2_ASAP7_75t_L g927 ( .A(n_844), .B(n_814), .Y(n_927) );
INVxp67_ASAP7_75t_L g928 ( .A(n_821), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_862), .Y(n_929) );
INVx1_ASAP7_75t_SL g930 ( .A(n_826), .Y(n_930) );
AND2x2_ASAP7_75t_L g931 ( .A(n_844), .B(n_808), .Y(n_931) );
AND2x2_ASAP7_75t_L g932 ( .A(n_845), .B(n_808), .Y(n_932) );
INVx3_ASAP7_75t_L g933 ( .A(n_843), .Y(n_933) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_826), .B(n_759), .Y(n_934) );
OR2x2_ASAP7_75t_L g935 ( .A(n_874), .B(n_814), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_882), .Y(n_936) );
OR2x2_ASAP7_75t_L g937 ( .A(n_834), .B(n_800), .Y(n_937) );
OR2x2_ASAP7_75t_L g938 ( .A(n_854), .B(n_800), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_872), .B(n_800), .Y(n_939) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_861), .Y(n_940) );
INVx4_ASAP7_75t_L g941 ( .A(n_832), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_828), .B(n_736), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_828), .B(n_752), .Y(n_943) );
BUFx3_ASAP7_75t_L g944 ( .A(n_882), .Y(n_944) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_879), .Y(n_945) );
BUFx3_ASAP7_75t_L g946 ( .A(n_866), .Y(n_946) );
INVx1_ASAP7_75t_L g947 ( .A(n_865), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_865), .Y(n_948) );
AND2x4_ASAP7_75t_L g949 ( .A(n_943), .B(n_853), .Y(n_949) );
OR2x2_ASAP7_75t_L g950 ( .A(n_900), .B(n_859), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_919), .Y(n_951) );
HB1xp67_ASAP7_75t_L g952 ( .A(n_945), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_922), .Y(n_953) );
INVxp67_ASAP7_75t_SL g954 ( .A(n_917), .Y(n_954) );
AND2x2_ASAP7_75t_L g955 ( .A(n_918), .B(n_868), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_918), .B(n_868), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_899), .B(n_857), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_895), .B(n_871), .Y(n_958) );
NOR2xp67_ASAP7_75t_L g959 ( .A(n_928), .B(n_887), .Y(n_959) );
OR2x2_ASAP7_75t_L g960 ( .A(n_900), .B(n_859), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_942), .B(n_859), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_925), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_892), .B(n_856), .Y(n_963) );
BUFx3_ASAP7_75t_L g964 ( .A(n_936), .Y(n_964) );
OR2x2_ASAP7_75t_L g965 ( .A(n_907), .B(n_823), .Y(n_965) );
NAND2x1_ASAP7_75t_L g966 ( .A(n_941), .B(n_853), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_940), .Y(n_967) );
OR2x2_ASAP7_75t_L g968 ( .A(n_907), .B(n_823), .Y(n_968) );
BUFx2_ASAP7_75t_L g969 ( .A(n_904), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_909), .B(n_876), .Y(n_970) );
INVx1_ASAP7_75t_L g971 ( .A(n_929), .Y(n_971) );
HB1xp67_ASAP7_75t_L g972 ( .A(n_923), .Y(n_972) );
AND2x4_ASAP7_75t_L g973 ( .A(n_943), .B(n_847), .Y(n_973) );
AND2x2_ASAP7_75t_L g974 ( .A(n_942), .B(n_820), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_921), .B(n_820), .Y(n_975) );
AND2x2_ASAP7_75t_L g976 ( .A(n_921), .B(n_823), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_891), .Y(n_977) );
AND2x4_ASAP7_75t_L g978 ( .A(n_908), .B(n_889), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_891), .Y(n_979) );
INVxp67_ASAP7_75t_SL g980 ( .A(n_934), .Y(n_980) );
OR2x2_ASAP7_75t_L g981 ( .A(n_916), .B(n_838), .Y(n_981) );
HB1xp67_ASAP7_75t_L g982 ( .A(n_944), .Y(n_982) );
INVx1_ASAP7_75t_L g983 ( .A(n_902), .Y(n_983) );
AND2x2_ASAP7_75t_L g984 ( .A(n_898), .B(n_838), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_927), .B(n_824), .Y(n_985) );
AND2x2_ASAP7_75t_L g986 ( .A(n_898), .B(n_870), .Y(n_986) );
INVx1_ASAP7_75t_SL g987 ( .A(n_930), .Y(n_987) );
BUFx3_ASAP7_75t_L g988 ( .A(n_946), .Y(n_988) );
AND2x2_ASAP7_75t_L g989 ( .A(n_901), .B(n_870), .Y(n_989) );
OR2x2_ASAP7_75t_L g990 ( .A(n_911), .B(n_840), .Y(n_990) );
INVx1_ASAP7_75t_L g991 ( .A(n_902), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_906), .Y(n_992) );
AND2x2_ASAP7_75t_SL g993 ( .A(n_941), .B(n_888), .Y(n_993) );
OR2x2_ASAP7_75t_L g994 ( .A(n_905), .B(n_883), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_926), .B(n_883), .Y(n_995) );
INVx1_ASAP7_75t_L g996 ( .A(n_913), .Y(n_996) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_931), .B(n_825), .Y(n_997) );
OR2x2_ASAP7_75t_L g998 ( .A(n_926), .B(n_883), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_913), .Y(n_999) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_935), .B(n_883), .Y(n_1000) );
INVx1_ASAP7_75t_SL g1001 ( .A(n_946), .Y(n_1001) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_932), .B(n_878), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_915), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1004 ( .A(n_920), .B(n_835), .Y(n_1004) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_951), .B(n_939), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1006 ( .A(n_953), .B(n_939), .Y(n_1006) );
INVx1_ASAP7_75t_SL g1007 ( .A(n_987), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1008 ( .A(n_950), .B(n_960), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_962), .B(n_947), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_967), .B(n_947), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_986), .B(n_903), .Y(n_1011) );
INVx1_ASAP7_75t_L g1012 ( .A(n_977), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_958), .B(n_948), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_985), .B(n_948), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_979), .Y(n_1015) );
AND2x2_ASAP7_75t_L g1016 ( .A(n_986), .B(n_903), .Y(n_1016) );
CKINVDCx20_ASAP7_75t_R g1017 ( .A(n_988), .Y(n_1017) );
INVx2_ASAP7_75t_L g1018 ( .A(n_971), .Y(n_1018) );
INVx1_ASAP7_75t_SL g1019 ( .A(n_1001), .Y(n_1019) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_964), .Y(n_1020) );
OR2x6_ASAP7_75t_L g1021 ( .A(n_966), .B(n_860), .Y(n_1021) );
NOR2xp33_ASAP7_75t_L g1022 ( .A(n_970), .B(n_850), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_997), .B(n_957), .Y(n_1023) );
AND2x2_ASAP7_75t_L g1024 ( .A(n_989), .B(n_894), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_989), .B(n_894), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_976), .B(n_961), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_983), .Y(n_1027) );
OR2x2_ASAP7_75t_L g1028 ( .A(n_950), .B(n_938), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1029 ( .A(n_976), .B(n_897), .Y(n_1029) );
AND2x2_ASAP7_75t_L g1030 ( .A(n_961), .B(n_897), .Y(n_1030) );
INVx1_ASAP7_75t_L g1031 ( .A(n_991), .Y(n_1031) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_984), .B(n_890), .Y(n_1032) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_965), .B(n_937), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_992), .Y(n_1034) );
NAND2x1p5_ASAP7_75t_L g1035 ( .A(n_966), .B(n_941), .Y(n_1035) );
INVx1_ASAP7_75t_L g1036 ( .A(n_996), .Y(n_1036) );
NAND2x1p5_ASAP7_75t_L g1037 ( .A(n_964), .B(n_910), .Y(n_1037) );
INVx1_ASAP7_75t_L g1038 ( .A(n_999), .Y(n_1038) );
INVx1_ASAP7_75t_L g1039 ( .A(n_1003), .Y(n_1039) );
AND2x2_ASAP7_75t_L g1040 ( .A(n_984), .B(n_890), .Y(n_1040) );
AND2x2_ASAP7_75t_L g1041 ( .A(n_955), .B(n_893), .Y(n_1041) );
NAND2xp5_ASAP7_75t_L g1042 ( .A(n_952), .B(n_924), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1009), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1010), .Y(n_1044) );
OR2x2_ASAP7_75t_L g1045 ( .A(n_1008), .B(n_968), .Y(n_1045) );
OR2x2_ASAP7_75t_L g1046 ( .A(n_1008), .B(n_968), .Y(n_1046) );
INVx2_ASAP7_75t_SL g1047 ( .A(n_1017), .Y(n_1047) );
OR2x2_ASAP7_75t_L g1048 ( .A(n_1026), .B(n_981), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1026), .B(n_1002), .Y(n_1049) );
AND2x4_ASAP7_75t_L g1050 ( .A(n_1021), .B(n_980), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g1051 ( .A(n_1030), .B(n_1002), .Y(n_1051) );
NOR2xp33_ASAP7_75t_L g1052 ( .A(n_1019), .B(n_972), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1053 ( .A(n_1024), .B(n_955), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1033), .B(n_981), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1018), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1056 ( .A(n_1017), .Y(n_1056) );
AND2x2_ASAP7_75t_L g1057 ( .A(n_1024), .B(n_956), .Y(n_1057) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1042), .Y(n_1058) );
AND2x2_ASAP7_75t_L g1059 ( .A(n_1025), .B(n_974), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_1032), .B(n_982), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_1040), .B(n_990), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_1040), .B(n_990), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1063 ( .A(n_1029), .B(n_963), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g1064 ( .A1(n_1047), .A2(n_959), .B1(n_1021), .B2(n_988), .Y(n_1064) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1047), .B(n_1007), .Y(n_1065) );
AND2x2_ASAP7_75t_L g1066 ( .A(n_1059), .B(n_1011), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1058), .B(n_1041), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1059), .B(n_1016), .Y(n_1068) );
INVxp67_ASAP7_75t_L g1069 ( .A(n_1052), .Y(n_1069) );
AOI222xp33_ASAP7_75t_L g1070 ( .A1(n_1043), .A2(n_1023), .B1(n_1022), .B2(n_1006), .C1(n_1005), .C2(n_1013), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1054), .Y(n_1071) );
AOI21xp5_ASAP7_75t_L g1072 ( .A1(n_1050), .A2(n_1021), .B(n_1035), .Y(n_1072) );
NAND2xp5_ASAP7_75t_L g1073 ( .A(n_1044), .B(n_1041), .Y(n_1073) );
NAND2xp5_ASAP7_75t_L g1074 ( .A(n_1053), .B(n_1029), .Y(n_1074) );
OA22x2_ASAP7_75t_L g1075 ( .A1(n_1056), .A2(n_1021), .B1(n_1020), .B2(n_860), .Y(n_1075) );
OAI22xp5_ASAP7_75t_L g1076 ( .A1(n_1056), .A2(n_1037), .B1(n_1035), .B2(n_860), .Y(n_1076) );
AOI211xp5_ASAP7_75t_L g1077 ( .A1(n_1050), .A2(n_975), .B(n_841), .C(n_864), .Y(n_1077) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_1045), .A2(n_1046), .B1(n_1035), .B2(n_1037), .C(n_1014), .Y(n_1078) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1068), .B(n_1053), .Y(n_1079) );
NAND2xp5_ASAP7_75t_L g1080 ( .A(n_1070), .B(n_1057), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1068), .B(n_1057), .Y(n_1081) );
AOI211xp5_ASAP7_75t_L g1082 ( .A1(n_1064), .A2(n_864), .B(n_1046), .C(n_1048), .Y(n_1082) );
OAI322xp33_ASAP7_75t_L g1083 ( .A1(n_1069), .A2(n_1060), .A3(n_1063), .B1(n_1062), .B2(n_1061), .C1(n_1049), .C2(n_1051), .Y(n_1083) );
INVxp67_ASAP7_75t_L g1084 ( .A(n_1065), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_1075), .A2(n_910), .B1(n_933), .B2(n_994), .Y(n_1085) );
OR2x2_ASAP7_75t_L g1086 ( .A(n_1071), .B(n_1028), .Y(n_1086) );
NOR2x1_ASAP7_75t_L g1087 ( .A(n_1078), .B(n_896), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1088 ( .A1(n_1065), .A2(n_1031), .B1(n_1012), .B2(n_1027), .C(n_1036), .Y(n_1088) );
OAI32xp33_ASAP7_75t_L g1089 ( .A1(n_1076), .A2(n_933), .A3(n_995), .B1(n_998), .B2(n_1000), .Y(n_1089) );
AOI211xp5_ASAP7_75t_L g1090 ( .A1(n_1072), .A2(n_912), .B(n_994), .C(n_1000), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1066), .B(n_978), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1092 ( .A1(n_1067), .A2(n_1015), .B1(n_1039), .B2(n_1038), .C(n_1034), .Y(n_1092) );
NAND3xp33_ASAP7_75t_SL g1093 ( .A(n_1077), .B(n_969), .C(n_914), .Y(n_1093) );
AOI21xp5_ASAP7_75t_L g1094 ( .A1(n_1073), .A2(n_993), .B(n_954), .Y(n_1094) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_1074), .A2(n_949), .B1(n_995), .B2(n_973), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_1075), .A2(n_949), .B1(n_978), .B2(n_973), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_1069), .B(n_873), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1070), .B(n_1055), .Y(n_1098) );
AOI211x1_ASAP7_75t_SL g1099 ( .A1(n_1098), .A2(n_1080), .B(n_1093), .C(n_1094), .Y(n_1099) );
NAND4xp25_ASAP7_75t_L g1100 ( .A(n_1097), .B(n_1087), .C(n_1082), .D(n_1096), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1084), .B(n_1081), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1102 ( .A(n_1092), .B(n_1088), .Y(n_1102) );
NOR3xp33_ASAP7_75t_SL g1103 ( .A(n_1085), .B(n_1089), .C(n_1083), .Y(n_1103) );
NOR3xp33_ASAP7_75t_L g1104 ( .A(n_1100), .B(n_1090), .C(n_1095), .Y(n_1104) );
NAND3x2_ASAP7_75t_L g1105 ( .A(n_1099), .B(n_1086), .C(n_1079), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1101), .B(n_1091), .Y(n_1106) );
NAND3xp33_ASAP7_75t_L g1107 ( .A(n_1103), .B(n_877), .C(n_832), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1106), .Y(n_1108) );
NAND2xp5_ASAP7_75t_L g1109 ( .A(n_1104), .B(n_1102), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1107), .Y(n_1110) );
XNOR2x1_ASAP7_75t_L g1111 ( .A(n_1109), .B(n_1105), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1110), .B(n_1108), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1113 ( .A(n_1112), .Y(n_1113) );
OR2x2_ASAP7_75t_L g1114 ( .A(n_1113), .B(n_1111), .Y(n_1114) );
AOI21xp5_ASAP7_75t_L g1115 ( .A1(n_1114), .A2(n_822), .B(n_1004), .Y(n_1115) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_1115), .B(n_842), .Y(n_1116) );
OR2x6_ASAP7_75t_L g1117 ( .A(n_1116), .B(n_885), .Y(n_1117) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_1117), .A2(n_875), .B1(n_889), .B2(n_973), .Y(n_1118) );
endmodule