module fake_jpeg_27023_n_28 (n_0, n_3, n_2, n_1, n_28);

input n_0;
input n_3;
input n_2;
input n_1;

output n_28;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_4;
wire n_16;
wire n_24;
wire n_26;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g4 ( 
.A(n_2),
.Y(n_4)
);

BUFx6f_ASAP7_75t_L g5 ( 
.A(n_3),
.Y(n_5)
);

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g7 ( 
.A(n_2),
.B(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_7),
.B(n_2),
.Y(n_8)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_4),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g9 ( 
.A(n_7),
.B(n_4),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_12),
.B(n_2),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_8),
.B(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_16),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_10),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_5),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_13),
.B1(n_5),
.B2(n_6),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_18),
.Y(n_22)
);

AO221x1_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_3),
.B1(n_6),
.B2(n_5),
.C(n_0),
.Y(n_21)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_20),
.C(n_0),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_SL g26 ( 
.A1(n_24),
.A2(n_25),
.B(n_0),
.C(n_1),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_21),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_26),
.A2(n_0),
.B(n_1),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_27),
.B(n_1),
.Y(n_28)
);


endmodule