module fake_aes_489_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
AND2x6_ASAP7_75t_L g11 ( .A(n_2), .B(n_3), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_5), .B(n_2), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_8), .B(n_1), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
BUFx12f_ASAP7_75t_L g15 ( .A(n_9), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
BUFx3_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_16), .B(n_0), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_12), .B(n_0), .C(n_6), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_16), .Y(n_21) );
NAND2xp33_ASAP7_75t_SL g22 ( .A(n_13), .B(n_10), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_19), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
BUFx3_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
BUFx3_ASAP7_75t_L g26 ( .A(n_18), .Y(n_26) );
AOI22xp33_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_19), .B1(n_11), .B2(n_22), .Y(n_27) );
OA21x2_ASAP7_75t_L g28 ( .A1(n_23), .A2(n_21), .B(n_20), .Y(n_28) );
AOI22xp33_ASAP7_75t_L g29 ( .A1(n_25), .A2(n_11), .B1(n_13), .B2(n_26), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_26), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_27), .Y(n_31) );
NOR2xp33_ASAP7_75t_L g32 ( .A(n_31), .B(n_25), .Y(n_32) );
NOR3xp33_ASAP7_75t_SL g33 ( .A(n_30), .B(n_11), .C(n_29), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_30), .Y(n_34) );
INVx1_ASAP7_75t_SL g35 ( .A(n_34), .Y(n_35) );
NOR2xp33_ASAP7_75t_R g36 ( .A(n_32), .B(n_11), .Y(n_36) );
INVx5_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
CKINVDCx16_ASAP7_75t_R g38 ( .A(n_36), .Y(n_38) );
NOR2x1_ASAP7_75t_L g39 ( .A(n_35), .B(n_11), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_39), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_41) );
endmodule