module real_aes_4744_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_1118, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_1119, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_1118;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_1119;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_1106;
wire n_522;
wire n_1092;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_1067;
wire n_518;
wire n_792;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_1091;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_1110;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_932;
wire n_399;
wire n_1021;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_948;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_1116;
wire n_573;
wire n_510;
wire n_1099;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_1108;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_1078;
wire n_495;
wire n_892;
wire n_994;
wire n_370;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_1098;
wire n_467;
wire n_875;
wire n_951;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_1049;
wire n_976;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1082;
wire n_468;
wire n_755;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_1025;
wire n_409;
wire n_860;
wire n_781;
wire n_748;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_1115;
wire n_504;
wire n_725;
wire n_455;
wire n_960;
wire n_1081;
wire n_671;
wire n_973;
wire n_1084;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_1100;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_1112;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1103;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1095;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_1080;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_334;
wire n_735;
wire n_569;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_853;
wire n_810;
wire n_1079;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1000;
wire n_1014;
wire n_1003;
wire n_366;
wire n_346;
wire n_1083;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_1085;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_1071;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_715;
wire n_959;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_359;
wire n_717;
wire n_1090;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_1114;
wire n_566;
wire n_719;
wire n_967;
wire n_837;
wire n_871;
wire n_1045;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1076;
wire n_396;
wire n_804;
wire n_1102;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_1104;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_797;
wire n_668;
wire n_862;
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_0), .A2(n_271), .B1(n_486), .B2(n_690), .Y(n_793) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1), .Y(n_1095) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_2), .A2(n_234), .B1(n_336), .B2(n_1109), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_3), .A2(n_212), .B1(n_486), .B2(n_498), .Y(n_654) );
INVx1_ASAP7_75t_L g521 ( .A(n_4), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_5), .A2(n_259), .B1(n_391), .B2(n_393), .Y(n_751) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_6), .A2(n_251), .B1(n_466), .B2(n_470), .Y(n_682) );
INVx1_ASAP7_75t_SL g923 ( .A(n_7), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_8), .A2(n_179), .B1(n_336), .B2(n_359), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_9), .A2(n_197), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g1098 ( .A(n_10), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_11), .A2(n_13), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_12), .A2(n_60), .B1(n_552), .B2(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g352 ( .A(n_14), .B(n_341), .Y(n_352) );
AOI21xp33_ASAP7_75t_L g598 ( .A1(n_15), .A2(n_599), .B(n_600), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g885 ( .A(n_16), .Y(n_885) );
INVx1_ASAP7_75t_L g1093 ( .A(n_17), .Y(n_1093) );
AOI221x1_ASAP7_75t_L g676 ( .A1(n_18), .A2(n_75), .B1(n_567), .B2(n_638), .C(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_19), .A2(n_292), .B1(n_535), .B2(n_540), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_20), .A2(n_245), .B1(n_537), .B2(n_552), .Y(n_646) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_21), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_22), .A2(n_27), .B1(n_371), .B2(n_588), .Y(n_752) );
INVx1_ASAP7_75t_L g575 ( .A(n_23), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g854 ( .A1(n_23), .A2(n_82), .B1(n_855), .B2(n_857), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_24), .A2(n_38), .B1(n_718), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_25), .A2(n_73), .B1(n_456), .B2(n_457), .Y(n_455) );
INVx1_ASAP7_75t_L g479 ( .A(n_26), .Y(n_479) );
AOI21xp33_ASAP7_75t_L g417 ( .A1(n_28), .A2(n_418), .B(n_419), .Y(n_417) );
INVx1_ASAP7_75t_L g798 ( .A(n_29), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_30), .A2(n_207), .B1(n_409), .B2(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_31), .A2(n_94), .B1(n_503), .B2(n_504), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_32), .A2(n_202), .B1(n_840), .B2(n_844), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_33), .B(n_572), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_34), .A2(n_260), .B1(n_393), .B2(n_590), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_35), .A2(n_45), .B1(n_371), .B2(n_375), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_36), .A2(n_191), .B1(n_336), .B2(n_540), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_37), .A2(n_254), .B1(n_453), .B2(n_725), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_39), .A2(n_112), .B1(n_503), .B2(n_504), .Y(n_789) );
INVx1_ASAP7_75t_L g883 ( .A(n_40), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_41), .A2(n_205), .B1(n_393), .B2(n_590), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_42), .A2(n_193), .B1(n_375), .B2(n_587), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_43), .A2(n_105), .B1(n_412), .B2(n_599), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g1100 ( .A1(n_44), .A2(n_295), .B1(n_484), .B2(n_1101), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_46), .A2(n_281), .B1(n_484), .B2(n_487), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_47), .A2(n_90), .B1(n_535), .B2(n_540), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_48), .B(n_490), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_49), .A2(n_119), .B1(n_678), .B2(n_771), .Y(n_770) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_50), .A2(n_307), .B1(n_379), .B2(n_386), .Y(n_611) );
OA22x2_ASAP7_75t_L g346 ( .A1(n_51), .A2(n_131), .B1(n_341), .B2(n_345), .Y(n_346) );
INVx1_ASAP7_75t_L g366 ( .A(n_51), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_52), .A2(n_159), .B1(n_412), .B2(n_616), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_53), .A2(n_268), .B1(n_495), .B2(n_501), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_54), .A2(n_93), .B1(n_409), .B2(n_412), .Y(n_408) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_55), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_56), .A2(n_301), .B1(n_336), .B2(n_500), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g390 ( .A1(n_57), .A2(n_185), .B1(n_391), .B2(n_393), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_58), .B(n_616), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_59), .A2(n_83), .B1(n_371), .B2(n_463), .Y(n_1071) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_61), .B(n_147), .Y(n_322) );
INVx1_ASAP7_75t_L g344 ( .A(n_61), .Y(n_344) );
OAI21xp33_ASAP7_75t_L g367 ( .A1(n_61), .A2(n_131), .B(n_368), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g804 ( .A1(n_62), .A2(n_213), .B1(n_458), .B2(n_463), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_63), .A2(n_211), .B1(n_779), .B2(n_781), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_64), .A2(n_222), .B1(n_379), .B2(n_386), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g1070 ( .A1(n_65), .A2(n_150), .B1(n_458), .B2(n_539), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_66), .A2(n_148), .B1(n_560), .B2(n_561), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_67), .A2(n_199), .B1(n_490), .B2(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g524 ( .A(n_68), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_69), .A2(n_187), .B1(n_539), .B2(n_555), .Y(n_554) );
AOI21xp33_ASAP7_75t_L g619 ( .A1(n_70), .A2(n_560), .B(n_620), .Y(n_619) );
XOR2x2_ASAP7_75t_L g505 ( .A(n_71), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g833 ( .A(n_72), .Y(n_833) );
AND2x4_ASAP7_75t_L g841 ( .A(n_72), .B(n_233), .Y(n_841) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_72), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_190), .B1(n_460), .B2(n_462), .Y(n_459) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_76), .A2(n_249), .B1(n_379), .B2(n_386), .Y(n_753) );
INVx1_ASAP7_75t_L g710 ( .A(n_77), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_78), .A2(n_126), .B1(n_397), .B2(n_725), .Y(n_809) );
INVx1_ASAP7_75t_L g528 ( .A(n_79), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_80), .A2(n_294), .B1(n_386), .B2(n_552), .Y(n_728) );
AO22x1_ASAP7_75t_L g608 ( .A1(n_81), .A2(n_267), .B1(n_463), .B2(n_609), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_84), .A2(n_100), .B1(n_466), .B2(n_470), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_85), .A2(n_122), .B1(n_397), .B2(n_399), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_86), .A2(n_188), .B1(n_397), .B2(n_412), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_87), .A2(n_118), .B1(n_371), .B2(n_475), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_88), .B(n_594), .Y(n_1064) );
INVx1_ASAP7_75t_L g800 ( .A(n_89), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_91), .A2(n_104), .B1(n_590), .B2(n_645), .Y(n_807) );
INVx1_ASAP7_75t_L g831 ( .A(n_92), .Y(n_831) );
AND2x4_ASAP7_75t_L g835 ( .A(n_92), .B(n_318), .Y(n_835) );
INVx1_ASAP7_75t_SL g856 ( .A(n_92), .Y(n_856) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_95), .B(n_594), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g731 ( .A1(n_96), .A2(n_99), .B1(n_539), .B2(n_555), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_97), .A2(n_171), .B1(n_473), .B2(n_475), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_98), .B(n_489), .Y(n_794) );
CKINVDCx16_ASAP7_75t_R g836 ( .A(n_101), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_102), .A2(n_121), .B1(n_829), .B2(n_894), .Y(n_893) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_103), .A2(n_224), .B1(n_590), .B2(n_1073), .Y(n_1072) );
INVx1_ASAP7_75t_L g580 ( .A(n_106), .Y(n_580) );
INVx1_ASAP7_75t_L g763 ( .A(n_107), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_108), .A2(n_272), .B1(n_495), .B2(n_498), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_109), .A2(n_226), .B1(n_497), .B2(n_498), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_110), .A2(n_225), .B1(n_537), .B2(n_552), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_111), .A2(n_136), .B1(n_465), .B2(n_468), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_113), .A2(n_219), .B1(n_573), .B2(n_638), .Y(n_637) );
AOI21xp5_ASAP7_75t_L g1066 ( .A1(n_114), .A2(n_560), .B(n_1067), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_115), .A2(n_221), .B1(n_494), .B2(n_497), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_116), .A2(n_164), .B1(n_572), .B2(n_573), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g635 ( .A1(n_117), .A2(n_196), .B1(n_526), .B2(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_120), .A2(n_285), .B1(n_774), .B2(n_775), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_123), .B(n_594), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_124), .A2(n_258), .B1(n_379), .B2(n_386), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_125), .A2(n_298), .B1(n_555), .B2(n_645), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_127), .A2(n_142), .B1(n_463), .B2(n_540), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_128), .A2(n_278), .B1(n_747), .B2(n_748), .Y(n_746) );
CKINVDCx6p67_ASAP7_75t_R g706 ( .A(n_129), .Y(n_706) );
INVx1_ASAP7_75t_L g358 ( .A(n_130), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_130), .B(n_182), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_130), .B(n_364), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_131), .B(n_242), .Y(n_321) );
XNOR2x1_ASAP7_75t_L g785 ( .A(n_132), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g332 ( .A(n_133), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_134), .A2(n_157), .B1(n_409), .B2(n_452), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_135), .A2(n_140), .B1(n_535), .B2(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_137), .B(n_418), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_138), .A2(n_155), .B1(n_500), .B2(n_501), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_139), .A2(n_218), .B1(n_460), .B2(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g1068 ( .A(n_141), .Y(n_1068) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_143), .A2(n_238), .B1(n_587), .B2(n_588), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g864 ( .A1(n_144), .A2(n_275), .B1(n_859), .B2(n_860), .Y(n_864) );
INVx1_ASAP7_75t_L g519 ( .A(n_145), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_146), .A2(n_162), .B1(n_515), .B2(n_517), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_147), .B(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_149), .A2(n_174), .B1(n_539), .B2(n_540), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_151), .A2(n_309), .B1(n_379), .B2(n_386), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_152), .A2(n_283), .B1(n_460), .B2(n_533), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_153), .A2(n_246), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_154), .A2(n_270), .B1(n_526), .B2(n_636), .Y(n_768) );
XNOR2x1_ASAP7_75t_L g630 ( .A(n_156), .B(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_158), .A2(n_290), .B1(n_453), .B2(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g838 ( .A(n_160), .Y(n_838) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_161), .A2(n_257), .B1(n_460), .B2(n_533), .Y(n_729) );
INVx1_ASAP7_75t_L g420 ( .A(n_163), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_165), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_166), .A2(n_195), .B1(n_379), .B2(n_386), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_167), .B(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_168), .A2(n_300), .B1(n_494), .B2(n_500), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_169), .A2(n_311), .B1(n_397), .B2(n_399), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_170), .A2(n_255), .B1(n_829), .B2(n_850), .Y(n_869) );
INVx1_ASAP7_75t_L g1088 ( .A(n_172), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_173), .A2(n_302), .B1(n_418), .B2(n_517), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_175), .A2(n_287), .B1(n_855), .B2(n_857), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_176), .A2(n_241), .B1(n_844), .B2(n_868), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_177), .A2(n_239), .B1(n_497), .B2(n_501), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_178), .A2(n_253), .B1(n_465), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_180), .A2(n_237), .B1(n_483), .B2(n_500), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_181), .A2(n_293), .B1(n_503), .B2(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g342 ( .A(n_182), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_183), .B(n_634), .Y(n_769) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_184), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g496 ( .A1(n_186), .A2(n_291), .B1(n_497), .B2(n_498), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_189), .A2(n_201), .B1(n_848), .B2(n_868), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_192), .A2(n_210), .B1(n_460), .B2(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g569 ( .A(n_194), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_198), .B(n_634), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g811 ( .A1(n_200), .A2(n_216), .B1(n_560), .B2(n_567), .C(n_812), .Y(n_811) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_203), .A2(n_434), .B(n_439), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_204), .A2(n_279), .B1(n_447), .B2(n_449), .Y(n_446) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_206), .A2(n_297), .B1(n_418), .B2(n_487), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_208), .A2(n_229), .B1(n_829), .B2(n_850), .Y(n_849) );
OAI21x1_ASAP7_75t_L g603 ( .A1(n_209), .A2(n_604), .B(n_623), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_209), .B(n_607), .Y(n_626) );
INVx1_ASAP7_75t_L g440 ( .A(n_214), .Y(n_440) );
INVx1_ASAP7_75t_L g720 ( .A(n_215), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_217), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g601 ( .A(n_220), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g1104 ( .A1(n_223), .A2(n_252), .B1(n_391), .B2(n_393), .Y(n_1104) );
INVx1_ASAP7_75t_L g509 ( .A(n_227), .Y(n_509) );
INVx1_ASAP7_75t_L g813 ( .A(n_228), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_230), .A2(n_247), .B1(n_840), .B2(n_848), .Y(n_847) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_231), .A2(n_565), .B(n_568), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_232), .A2(n_263), .B1(n_555), .B2(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_233), .Y(n_323) );
AND2x4_ASAP7_75t_L g832 ( .A(n_233), .B(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_235), .A2(n_240), .B1(n_495), .B2(n_501), .Y(n_661) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_236), .Y(n_691) );
INVx1_ASAP7_75t_L g356 ( .A(n_242), .Y(n_356) );
INVxp67_ASAP7_75t_L g407 ( .A(n_242), .Y(n_407) );
INVx1_ASAP7_75t_L g621 ( .A(n_243), .Y(n_621) );
INVx1_ASAP7_75t_L g712 ( .A(n_244), .Y(n_712) );
INVxp67_ASAP7_75t_R g842 ( .A(n_248), .Y(n_842) );
INVx2_ASAP7_75t_L g318 ( .A(n_250), .Y(n_318) );
INVx1_ASAP7_75t_SL g675 ( .A(n_255), .Y(n_675) );
NOR3xp33_ASAP7_75t_L g702 ( .A(n_255), .B(n_703), .C(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g1090 ( .A(n_256), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_261), .A2(n_262), .B1(n_486), .B2(n_487), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g796 ( .A1(n_264), .A2(n_483), .B(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_265), .A2(n_273), .B1(n_483), .B2(n_484), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_266), .A2(n_276), .B1(n_412), .B2(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g716 ( .A(n_269), .Y(n_716) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_274), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g1059 ( .A(n_275), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_275), .A2(n_1080), .B1(n_1110), .B2(n_1112), .Y(n_1079) );
INVx1_ASAP7_75t_L g881 ( .A(n_277), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_280), .A2(n_284), .B1(n_412), .B2(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g754 ( .A(n_282), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_286), .A2(n_306), .B1(n_489), .B2(n_490), .Y(n_488) );
AND2x2_ASAP7_75t_L g677 ( .A(n_288), .B(n_678), .Y(n_677) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_289), .A2(n_304), .B1(n_532), .B2(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g1080 ( .A1(n_296), .A2(n_1081), .B1(n_1082), .B2(n_1083), .Y(n_1080) );
CKINVDCx5p33_ASAP7_75t_R g1081 ( .A(n_296), .Y(n_1081) );
INVx1_ASAP7_75t_L g924 ( .A(n_299), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_303), .A2(n_310), .B1(n_597), .B2(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g722 ( .A(n_305), .Y(n_722) );
XOR2x2_ASAP7_75t_L g430 ( .A(n_308), .B(n_431), .Y(n_430) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_324), .B(n_819), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
BUFx4_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .C(n_323), .Y(n_315) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_316), .B(n_1077), .Y(n_1076) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_316), .B(n_1078), .Y(n_1111) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_316), .A2(n_323), .B(n_856), .Y(n_1116) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AO21x1_ASAP7_75t_L g1113 ( .A1(n_317), .A2(n_1114), .B(n_1116), .Y(n_1113) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g830 ( .A(n_318), .B(n_831), .Y(n_830) );
AND3x4_ASAP7_75t_L g855 ( .A(n_318), .B(n_832), .C(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g1077 ( .A(n_319), .B(n_1078), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_320), .A2(n_424), .B(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g1078 ( .A(n_323), .Y(n_1078) );
XNOR2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_542), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_427), .B2(n_428), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
XNOR2x1_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
CKINVDCx5p33_ASAP7_75t_R g331 ( .A(n_332), .Y(n_331) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_395), .Y(n_333) );
NAND4xp25_ASAP7_75t_L g334 ( .A(n_335), .B(n_370), .C(n_378), .D(n_390), .Y(n_334) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_337), .Y(n_463) );
BUFx6f_ASAP7_75t_L g535 ( .A(n_337), .Y(n_535) );
BUFx3_ASAP7_75t_L g774 ( .A(n_337), .Y(n_774) );
AND2x4_ASAP7_75t_L g337 ( .A(n_338), .B(n_347), .Y(n_337) );
AND2x2_ASAP7_75t_L g372 ( .A(n_338), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g398 ( .A(n_338), .B(n_384), .Y(n_398) );
AND2x2_ASAP7_75t_L g418 ( .A(n_338), .B(n_388), .Y(n_418) );
AND2x2_ASAP7_75t_L g438 ( .A(n_338), .B(n_388), .Y(n_438) );
AND2x2_ASAP7_75t_L g461 ( .A(n_338), .B(n_373), .Y(n_461) );
AND2x4_ASAP7_75t_L g486 ( .A(n_338), .B(n_384), .Y(n_486) );
AND2x4_ASAP7_75t_L g494 ( .A(n_338), .B(n_369), .Y(n_494) );
AND2x4_ASAP7_75t_L g500 ( .A(n_338), .B(n_373), .Y(n_500) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_346), .Y(n_338) );
INVx1_ASAP7_75t_L g382 ( .A(n_339), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
NAND2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx2_ASAP7_75t_L g345 ( .A(n_341), .Y(n_345) );
INVx3_ASAP7_75t_L g351 ( .A(n_341), .Y(n_351) );
NAND2xp33_ASAP7_75t_L g357 ( .A(n_341), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g368 ( .A(n_341), .Y(n_368) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_341), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_342), .B(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OAI21xp5_ASAP7_75t_L g406 ( .A1(n_344), .A2(n_368), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
AND2x2_ASAP7_75t_L g405 ( .A(n_346), .B(n_406), .Y(n_405) );
AND2x2_ASAP7_75t_L g411 ( .A(n_346), .B(n_382), .Y(n_411) );
AND2x4_ASAP7_75t_L g498 ( .A(n_347), .B(n_381), .Y(n_498) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g369 ( .A(n_348), .Y(n_369) );
OR2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_353), .Y(n_348) );
AND2x4_ASAP7_75t_L g373 ( .A(n_349), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g384 ( .A(n_349), .B(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
AND2x2_ASAP7_75t_L g401 ( .A(n_349), .B(n_402), .Y(n_401) );
AND2x4_ASAP7_75t_L g349 ( .A(n_350), .B(n_352), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_351), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g364 ( .A(n_351), .Y(n_364) );
NAND3xp33_ASAP7_75t_L g425 ( .A(n_352), .B(n_363), .C(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g385 ( .A(n_354), .Y(n_385) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g458 ( .A(n_360), .Y(n_458) );
INVx5_ASAP7_75t_L g609 ( .A(n_360), .Y(n_609) );
INVx1_ASAP7_75t_L g643 ( .A(n_360), .Y(n_643) );
INVx1_ASAP7_75t_L g775 ( .A(n_360), .Y(n_775) );
INVx3_ASAP7_75t_L g1109 ( .A(n_360), .Y(n_1109) );
INVx6_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx12f_ASAP7_75t_L g540 ( .A(n_361), .Y(n_540) );
AND2x4_ASAP7_75t_L g361 ( .A(n_362), .B(n_369), .Y(n_361) );
AND2x4_ASAP7_75t_L g377 ( .A(n_362), .B(n_373), .Y(n_377) );
AND2x4_ASAP7_75t_L g413 ( .A(n_362), .B(n_388), .Y(n_413) );
AND2x4_ASAP7_75t_L g487 ( .A(n_362), .B(n_388), .Y(n_487) );
AND2x4_ASAP7_75t_L g495 ( .A(n_362), .B(n_369), .Y(n_495) );
AND2x4_ASAP7_75t_L g501 ( .A(n_362), .B(n_373), .Y(n_501) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x4_ASAP7_75t_L g394 ( .A(n_369), .B(n_381), .Y(n_394) );
BUFx4f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_372), .Y(n_587) );
AND2x4_ASAP7_75t_L g392 ( .A(n_373), .B(n_381), .Y(n_392) );
AND2x4_ASAP7_75t_L g497 ( .A(n_373), .B(n_381), .Y(n_497) );
INVx2_ASAP7_75t_SL g375 ( .A(n_376), .Y(n_375) );
INVx4_ASAP7_75t_L g475 ( .A(n_376), .Y(n_475) );
INVx4_ASAP7_75t_L g533 ( .A(n_376), .Y(n_533) );
INVx4_ASAP7_75t_L g588 ( .A(n_376), .Y(n_588) );
INVx1_ASAP7_75t_L g648 ( .A(n_376), .Y(n_648) );
INVx1_ASAP7_75t_L g781 ( .A(n_376), .Y(n_781) );
INVx2_ASAP7_75t_L g1073 ( .A(n_376), .Y(n_1073) );
INVx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx12f_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx3_ASAP7_75t_L g467 ( .A(n_380), .Y(n_467) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_380), .Y(n_552) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
AND2x2_ASAP7_75t_L g387 ( .A(n_381), .B(n_388), .Y(n_387) );
AND2x4_ASAP7_75t_L g503 ( .A(n_381), .B(n_384), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_381), .B(n_388), .Y(n_504) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x4_ASAP7_75t_L g410 ( .A(n_384), .B(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g483 ( .A(n_384), .B(n_411), .Y(n_483) );
AND2x4_ASAP7_75t_L g388 ( .A(n_385), .B(n_389), .Y(n_388) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g471 ( .A(n_387), .Y(n_471) );
BUFx5_ASAP7_75t_L g537 ( .A(n_387), .Y(n_537) );
AND2x4_ASAP7_75t_L g416 ( .A(n_388), .B(n_411), .Y(n_416) );
AND2x2_ASAP7_75t_L g489 ( .A(n_388), .B(n_411), .Y(n_489) );
INVx1_ASAP7_75t_L g474 ( .A(n_391), .Y(n_474) );
BUFx12f_ASAP7_75t_L g532 ( .A(n_391), .Y(n_532) );
BUFx12f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_392), .Y(n_555) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_392), .Y(n_590) );
BUFx3_ASAP7_75t_L g456 ( .A(n_393), .Y(n_456) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_394), .Y(n_539) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_394), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_396), .B(n_408), .C(n_414), .D(n_417), .Y(n_395) );
INVx3_ASAP7_75t_L g1091 ( .A(n_397), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
BUFx3_ASAP7_75t_L g453 ( .A(n_398), .Y(n_453) );
INVx2_ASAP7_75t_L g563 ( .A(n_398), .Y(n_563) );
INVx2_ASAP7_75t_SL g441 ( .A(n_399), .Y(n_441) );
BUFx4f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx5_ASAP7_75t_L g516 ( .A(n_400), .Y(n_516) );
BUFx2_ASAP7_75t_L g725 ( .A(n_400), .Y(n_725) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_405), .Y(n_400) );
AND2x2_ASAP7_75t_L g484 ( .A(n_401), .B(n_405), .Y(n_484) );
AND2x4_ASAP7_75t_L g690 ( .A(n_401), .B(n_405), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g424 ( .A(n_403), .Y(n_424) );
BUFx3_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g527 ( .A(n_410), .Y(n_527) );
BUFx6f_ASAP7_75t_L g560 ( .A(n_410), .Y(n_560) );
BUFx3_ASAP7_75t_L g745 ( .A(n_410), .Y(n_745) );
INVx3_ASAP7_75t_L g1096 ( .A(n_412), .Y(n_1096) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_413), .Y(n_450) );
INVx3_ASAP7_75t_L g574 ( .A(n_413), .Y(n_574) );
INVx2_ASAP7_75t_L g520 ( .A(n_415), .Y(n_520) );
BUFx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g448 ( .A(n_416), .Y(n_448) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_416), .Y(n_599) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_416), .Y(n_616) );
BUFx8_ASAP7_75t_SL g638 ( .A(n_416), .Y(n_638) );
INVx2_ASAP7_75t_L g719 ( .A(n_416), .Y(n_719) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_421), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g748 ( .A(n_421), .Y(n_748) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g490 ( .A(n_422), .Y(n_490) );
INVx2_ASAP7_75t_SL g517 ( .A(n_422), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g797 ( .A(n_422), .B(n_798), .Y(n_797) );
BUFx6f_ASAP7_75t_L g814 ( .A(n_422), .Y(n_814) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx3_ASAP7_75t_L g445 ( .A(n_423), .Y(n_445) );
INVx2_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
AO22x2_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_476), .B2(n_541), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_432), .B(n_454), .Y(n_431) );
NAND3xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_446), .C(n_451), .Y(n_432) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g567 ( .A(n_437), .Y(n_567) );
INVx2_ASAP7_75t_L g594 ( .A(n_437), .Y(n_594) );
INVx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g513 ( .A(n_438), .Y(n_513) );
BUFx3_ASAP7_75t_L g747 ( .A(n_438), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_441), .B(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_444), .B(n_601), .Y(n_600) );
INVx4_ASAP7_75t_L g640 ( .A(n_444), .Y(n_640) );
INVx4_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_L g679 ( .A(n_445), .Y(n_679) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g572 ( .A(n_448), .Y(n_572) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx4_ASAP7_75t_L g522 ( .A(n_450), .Y(n_522) );
BUFx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g529 ( .A(n_453), .Y(n_529) );
NAND4xp25_ASAP7_75t_L g454 ( .A(n_455), .B(n_459), .C(n_464), .D(n_472), .Y(n_454) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx8_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g780 ( .A(n_461), .Y(n_780) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx4f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_470), .Y(n_553) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g541 ( .A(n_476), .Y(n_541) );
XNOR2x1_ASAP7_75t_L g476 ( .A(n_477), .B(n_505), .Y(n_476) );
INVx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
XNOR2x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
OR2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
NAND4xp25_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .C(n_488), .D(n_491), .Y(n_481) );
INVx2_ASAP7_75t_L g695 ( .A(n_483), .Y(n_695) );
INVx2_ASAP7_75t_L g697 ( .A(n_486), .Y(n_697) );
INVx2_ASAP7_75t_L g692 ( .A(n_487), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g492 ( .A(n_493), .B(n_496), .C(n_499), .D(n_502), .Y(n_492) );
NAND2x1_ASAP7_75t_L g506 ( .A(n_507), .B(n_530), .Y(n_506) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_518), .C(n_523), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_510), .B(n_514), .Y(n_508) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx2_ASAP7_75t_L g634 ( .A(n_512), .Y(n_634) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_516), .A2(n_569), .B(n_570), .Y(n_568) );
INVx4_ASAP7_75t_L g597 ( .A(n_516), .Y(n_597) );
INVx2_ASAP7_75t_L g771 ( .A(n_516), .Y(n_771) );
INVx2_ASAP7_75t_L g1063 ( .A(n_516), .Y(n_1063) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_518) );
OAI22xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_528), .B2(n_529), .Y(n_523) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND4x1_ASAP7_75t_L g530 ( .A(n_531), .B(n_534), .C(n_536), .D(n_538), .Y(n_530) );
XOR2xp5_ASAP7_75t_L g542 ( .A(n_543), .B(n_665), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B1(n_628), .B2(n_664), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
OA22x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_576), .B2(n_577), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_575), .Y(n_548) );
NOR2x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_558), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .C(n_556), .D(n_557), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_564), .C(n_571), .Y(n_558) );
INVx4_ASAP7_75t_L g711 ( .A(n_560), .Y(n_711) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g636 ( .A(n_562), .Y(n_636) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g714 ( .A(n_563), .Y(n_714) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g723 ( .A(n_567), .Y(n_723) );
INVx3_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
OAI22xp5_ASAP7_75t_L g715 ( .A1(n_574), .A2(n_716), .B1(n_717), .B2(n_720), .Y(n_715) );
INVx2_ASAP7_75t_L g767 ( .A(n_574), .Y(n_767) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_602), .B1(n_603), .B2(n_627), .Y(n_578) );
INVx1_ASAP7_75t_L g627 ( .A(n_579), .Y(n_627) );
XNOR2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
NOR4xp75_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .C(n_591), .D(n_595), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g595 ( .A(n_596), .B(n_598), .Y(n_595) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_613), .Y(n_604) );
NOR3xp33_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .C(n_610), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g625 ( .A(n_608), .B(n_618), .C(n_626), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_610), .B(n_614), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_618), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
INVx2_ASAP7_75t_L g1094 ( .A(n_616), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g664 ( .A(n_628), .Y(n_664) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AO22x2_ASAP7_75t_L g629 ( .A1(n_630), .A2(n_649), .B1(n_662), .B2(n_663), .Y(n_629) );
INVx2_ASAP7_75t_L g662 ( .A(n_630), .Y(n_662) );
OR2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_641), .Y(n_631) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .C(n_637), .D(n_639), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .C(n_646), .D(n_647), .Y(n_641) );
INVx1_ASAP7_75t_L g663 ( .A(n_649), .Y(n_663) );
INVxp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_657), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .C(n_655), .D(n_656), .Y(n_652) );
NAND4xp25_ASAP7_75t_L g657 ( .A(n_658), .B(n_659), .C(n_660), .D(n_661), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_759), .B2(n_760), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AO22x2_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_734), .B1(n_755), .B2(n_756), .Y(n_667) );
INVx2_ASAP7_75t_L g755 ( .A(n_668), .Y(n_755) );
OAI22xp5_ASAP7_75t_SL g668 ( .A1(n_669), .A2(n_670), .B1(n_705), .B2(n_733), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2x1_ASAP7_75t_L g671 ( .A(n_672), .B(n_698), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_673), .B(n_680), .C(n_684), .Y(n_672) );
OAI22xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_676), .B2(n_1118), .Y(n_673) );
INVx1_ASAP7_75t_L g703 ( .A(n_674), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g680 ( .A(n_675), .B(n_681), .Y(n_680) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_675), .A2(n_685), .B1(n_686), .B2(n_1119), .Y(n_684) );
INVx1_ASAP7_75t_L g700 ( .A(n_676), .Y(n_700) );
INVx4_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_681), .B(n_699), .C(n_702), .Y(n_698) );
AND2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
INVx1_ASAP7_75t_L g704 ( .A(n_685), .Y(n_704) );
INVx1_ASAP7_75t_L g701 ( .A(n_686), .Y(n_701) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_687), .B(n_693), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_691), .B2(n_692), .Y(n_687) );
INVx4_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_696), .B2(n_697), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_705), .Y(n_733) );
XNOR2x1_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_706), .A2(n_828), .B1(n_834), .B2(n_836), .Y(n_827) );
NAND2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_726), .Y(n_707) );
NOR3xp33_ASAP7_75t_SL g708 ( .A(n_709), .B(n_715), .C(n_721), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_711), .B1(n_712), .B2(n_713), .Y(n_709) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
OAI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_724), .Y(n_721) );
NOR2x1_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g758 ( .A(n_737), .Y(n_758) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
XOR2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_754), .Y(n_739) );
NOR2x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_749), .Y(n_740) );
NAND4xp25_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .C(n_744), .D(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g1089 ( .A(n_745), .Y(n_1089) );
INVx2_ASAP7_75t_L g1099 ( .A(n_747), .Y(n_1099) );
NAND4xp25_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .C(n_752), .D(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_782), .B1(n_816), .B2(n_817), .Y(n_760) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g816 ( .A(n_762), .Y(n_816) );
XNOR2x1_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_763), .A2(n_834), .B1(n_880), .B2(n_881), .Y(n_879) );
OR2x2_ASAP7_75t_L g764 ( .A(n_765), .B(n_772), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .C(n_769), .D(n_770), .Y(n_765) );
NAND4xp25_ASAP7_75t_L g772 ( .A(n_773), .B(n_776), .C(n_777), .D(n_778), .Y(n_772) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx3_ASAP7_75t_L g818 ( .A(n_783), .Y(n_818) );
AO22x2_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_785), .B1(n_799), .B2(n_815), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
OR2x2_ASAP7_75t_L g786 ( .A(n_787), .B(n_792), .Y(n_786) );
NAND4xp25_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .C(n_790), .D(n_791), .Y(n_787) );
NAND4xp25_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .C(n_795), .D(n_796), .Y(n_792) );
INVx1_ASAP7_75t_L g815 ( .A(n_799), .Y(n_815) );
XNOR2x1_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .C(n_808), .D(n_811), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_L g805 ( .A(n_806), .B(n_807), .Y(n_805) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_814), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g1067 ( .A(n_814), .B(n_1068), .Y(n_1067) );
INVx1_ASAP7_75t_L g1101 ( .A(n_814), .Y(n_1101) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_1052), .B1(n_1054), .B2(n_1075), .C(n_1079), .Y(n_819) );
AOI211xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_965), .B(n_1013), .C(n_1038), .Y(n_820) );
NAND5xp2_ASAP7_75t_L g821 ( .A(n_822), .B(n_900), .C(n_929), .D(n_938), .E(n_958), .Y(n_821) );
NOR3xp33_ASAP7_75t_SL g822 ( .A(n_823), .B(n_870), .C(n_888), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_825), .B(n_851), .Y(n_824) );
INVx1_ASAP7_75t_L g950 ( .A(n_825), .Y(n_950) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_825), .A2(n_967), .B1(n_969), .B2(n_970), .C(n_971), .Y(n_966) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_825), .B(n_897), .Y(n_978) );
NAND2xp5_ASAP7_75t_L g1032 ( .A(n_825), .B(n_877), .Y(n_1032) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_845), .Y(n_825) );
AND2x2_ASAP7_75t_L g887 ( .A(n_826), .B(n_846), .Y(n_887) );
INVx2_ASAP7_75t_L g904 ( .A(n_826), .Y(n_904) );
INVx3_ASAP7_75t_L g911 ( .A(n_826), .Y(n_911) );
OR2x2_ASAP7_75t_L g940 ( .A(n_826), .B(n_846), .Y(n_940) );
NOR2xp33_ASAP7_75t_L g957 ( .A(n_826), .B(n_878), .Y(n_957) );
OR2x2_ASAP7_75t_L g826 ( .A(n_827), .B(n_837), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g922 ( .A1(n_828), .A2(n_834), .B1(n_923), .B2(n_924), .C(n_925), .Y(n_922) );
INVx3_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_830), .B(n_832), .Y(n_829) );
AND2x4_ASAP7_75t_L g840 ( .A(n_830), .B(n_841), .Y(n_840) );
AND2x2_ASAP7_75t_L g859 ( .A(n_830), .B(n_841), .Y(n_859) );
AND2x2_ASAP7_75t_L g868 ( .A(n_830), .B(n_841), .Y(n_868) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_832), .B(n_835), .Y(n_834) );
AND2x4_ASAP7_75t_L g850 ( .A(n_832), .B(n_835), .Y(n_850) );
AND2x4_ASAP7_75t_L g857 ( .A(n_832), .B(n_835), .Y(n_857) );
AND2x4_ASAP7_75t_L g844 ( .A(n_835), .B(n_841), .Y(n_844) );
AND2x2_ASAP7_75t_L g848 ( .A(n_835), .B(n_841), .Y(n_848) );
AND2x2_ASAP7_75t_L g860 ( .A(n_835), .B(n_841), .Y(n_860) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_839), .B1(n_842), .B2(n_843), .Y(n_837) );
INVx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g1053 ( .A(n_840), .Y(n_1053) );
INVx2_ASAP7_75t_L g843 ( .A(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_845), .B(n_890), .Y(n_889) );
INVx3_ASAP7_75t_L g920 ( .A(n_845), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_845), .B(n_891), .Y(n_1030) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_845), .B(n_891), .Y(n_1051) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
AND2x2_ASAP7_75t_L g910 ( .A(n_846), .B(n_911), .Y(n_910) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_846), .B(n_891), .Y(n_1026) );
AND2x2_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .Y(n_846) );
O2A1O1Ixp33_ASAP7_75t_L g974 ( .A1(n_851), .A2(n_964), .B(n_975), .C(n_977), .Y(n_974) );
AOI222xp33_ASAP7_75t_L g1023 ( .A1(n_851), .A2(n_1024), .B1(n_1026), .B2(n_1027), .C1(n_1028), .C2(n_1031), .Y(n_1023) );
NAND2xp5_ASAP7_75t_L g1025 ( .A(n_851), .B(n_877), .Y(n_1025) );
AND2x2_ASAP7_75t_L g851 ( .A(n_852), .B(n_861), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_852), .B(n_872), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_852), .B(n_874), .Y(n_932) );
AND2x2_ASAP7_75t_SL g937 ( .A(n_852), .B(n_907), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g961 ( .A(n_852), .B(n_962), .Y(n_961) );
AND2x2_ASAP7_75t_L g968 ( .A(n_852), .B(n_877), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g987 ( .A(n_852), .B(n_878), .Y(n_987) );
AND2x2_ASAP7_75t_L g999 ( .A(n_852), .B(n_865), .Y(n_999) );
A2O1A1Ixp33_ASAP7_75t_L g1033 ( .A1(n_852), .A2(n_1034), .B(n_1035), .C(n_1036), .Y(n_1033) );
CKINVDCx6p67_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
AND2x2_ASAP7_75t_L g899 ( .A(n_853), .B(n_861), .Y(n_899) );
AND2x2_ASAP7_75t_L g906 ( .A(n_853), .B(n_907), .Y(n_906) );
INVx1_ASAP7_75t_L g915 ( .A(n_853), .Y(n_915) );
OR2x2_ASAP7_75t_L g984 ( .A(n_853), .B(n_862), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_853), .B(n_874), .Y(n_1003) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_853), .B(n_969), .Y(n_1035) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_853), .B(n_862), .Y(n_1043) );
AND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_858), .Y(n_853) );
INVx1_ASAP7_75t_L g880 ( .A(n_855), .Y(n_880) );
INVx2_ASAP7_75t_SL g895 ( .A(n_857), .Y(n_895) );
INVx1_ASAP7_75t_L g886 ( .A(n_859), .Y(n_886) );
INVx1_ASAP7_75t_L g884 ( .A(n_860), .Y(n_884) );
INVx1_ASAP7_75t_L g1011 ( .A(n_861), .Y(n_1011) );
OR2x2_ASAP7_75t_L g1034 ( .A(n_861), .B(n_907), .Y(n_1034) );
AND2x2_ASAP7_75t_L g861 ( .A(n_862), .B(n_865), .Y(n_861) );
AND2x2_ASAP7_75t_L g872 ( .A(n_862), .B(n_866), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g875 ( .A(n_862), .Y(n_875) );
AND2x4_ASAP7_75t_SL g862 ( .A(n_863), .B(n_864), .Y(n_862) );
AND2x2_ASAP7_75t_L g874 ( .A(n_865), .B(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g913 ( .A(n_865), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g941 ( .A(n_865), .B(n_914), .Y(n_941) );
AND2x2_ASAP7_75t_L g956 ( .A(n_865), .B(n_914), .Y(n_956) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
AND2x2_ASAP7_75t_L g907 ( .A(n_866), .B(n_875), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_867), .B(n_869), .Y(n_866) );
AOI21xp33_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_873), .B(n_876), .Y(n_870) );
INVx1_ASAP7_75t_L g1019 ( .A(n_871), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1045 ( .A(n_871), .B(n_1046), .Y(n_1045) );
AND2x2_ASAP7_75t_L g952 ( .A(n_872), .B(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g962 ( .A(n_872), .Y(n_962) );
AND2x2_ASAP7_75t_L g969 ( .A(n_872), .B(n_878), .Y(n_969) );
AND2x2_ASAP7_75t_L g1021 ( .A(n_872), .B(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
AND2x2_ASAP7_75t_L g948 ( .A(n_874), .B(n_878), .Y(n_948) );
OAI321xp33_ASAP7_75t_L g986 ( .A1(n_874), .A2(n_912), .A3(n_951), .B1(n_985), .B2(n_987), .C(n_988), .Y(n_986) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_874), .B(n_953), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g918 ( .A(n_875), .B(n_914), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g876 ( .A(n_877), .B(n_887), .Y(n_876) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_877), .B(n_918), .Y(n_917) );
AND2x2_ASAP7_75t_L g953 ( .A(n_877), .B(n_914), .Y(n_953) );
NOR2x1p5_ASAP7_75t_L g983 ( .A(n_877), .B(n_984), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_877), .B(n_920), .Y(n_997) );
INVx1_ASAP7_75t_L g1008 ( .A(n_877), .Y(n_1008) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_877), .B(n_911), .Y(n_1049) );
CKINVDCx6p67_ASAP7_75t_R g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g898 ( .A(n_878), .Y(n_898) );
AND2x2_ASAP7_75t_L g905 ( .A(n_878), .B(n_906), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_878), .B(n_941), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g989 ( .A(n_878), .B(n_911), .Y(n_989) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_878), .B(n_1011), .Y(n_1010) );
OR2x6_ASAP7_75t_SL g878 ( .A(n_879), .B(n_882), .Y(n_878) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B1(n_885), .B2(n_886), .Y(n_882) );
INVx1_ASAP7_75t_L g972 ( .A(n_887), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_887), .B(n_891), .Y(n_1037) );
NOR2xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_896), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g930 ( .A(n_889), .B(n_897), .Y(n_930) );
INVx1_ASAP7_75t_L g1044 ( .A(n_889), .Y(n_1044) );
NOR2xp33_ASAP7_75t_L g927 ( .A(n_890), .B(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g945 ( .A(n_890), .Y(n_945) );
HB1xp67_ASAP7_75t_L g990 ( .A(n_890), .Y(n_990) );
INVx3_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g934 ( .A(n_891), .Y(n_934) );
AND2x2_ASAP7_75t_L g964 ( .A(n_891), .B(n_939), .Y(n_964) );
AND2x4_ASAP7_75t_L g891 ( .A(n_892), .B(n_893), .Y(n_891) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_897), .B(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_897), .B(n_937), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g1018 ( .A(n_897), .B(n_956), .Y(n_1018) );
INVx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g1046 ( .A(n_899), .Y(n_1046) );
OAI21xp33_ASAP7_75t_L g900 ( .A1(n_901), .A2(n_908), .B(n_926), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g902 ( .A(n_903), .B(n_905), .Y(n_902) );
INVx2_ASAP7_75t_L g970 ( .A(n_903), .Y(n_970) );
BUFx2_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_904), .B(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g993 ( .A(n_904), .Y(n_993) );
AND2x2_ASAP7_75t_L g1020 ( .A(n_904), .B(n_1021), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g1042 ( .A(n_904), .B(n_1043), .Y(n_1042) );
AND2x2_ASAP7_75t_L g967 ( .A(n_907), .B(n_968), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_912), .B1(n_916), .B2(n_919), .C(n_921), .Y(n_908) );
INVx1_ASAP7_75t_L g1000 ( .A(n_910), .Y(n_1000) );
O2A1O1Ixp33_ASAP7_75t_L g1014 ( .A1(n_910), .A2(n_1015), .B(n_1019), .C(n_1020), .Y(n_1014) );
INVx1_ASAP7_75t_L g982 ( .A(n_911), .Y(n_982) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_911), .B(n_945), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1039 ( .A(n_911), .B(n_952), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_912), .B(n_932), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g977 ( .A(n_912), .B(n_978), .Y(n_977) );
O2A1O1Ixp33_ASAP7_75t_L g1006 ( .A1(n_912), .A2(n_1007), .B(n_1009), .C(n_1012), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
AND2x2_ASAP7_75t_L g994 ( .A(n_914), .B(n_948), .Y(n_994) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_917), .B(n_1017), .Y(n_1016) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_918), .A2(n_997), .B1(n_998), .B2(n_1000), .Y(n_996) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_919), .B(n_955), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g971 ( .A1(n_919), .A2(n_928), .B1(n_960), .B2(n_972), .C(n_973), .Y(n_971) );
INVx3_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g946 ( .A1(n_920), .A2(n_947), .B1(n_949), .B2(n_951), .Y(n_946) );
INVx1_ASAP7_75t_L g985 ( .A(n_920), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_920), .A2(n_943), .B1(n_1039), .B2(n_1040), .C(n_1041), .Y(n_1038) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
BUFx3_ASAP7_75t_L g928 ( .A(n_922), .Y(n_928) );
INVx1_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
AOI22xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_931), .B1(n_933), .B2(n_935), .Y(n_929) );
INVx1_ASAP7_75t_L g1012 ( .A(n_933), .Y(n_1012) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
AOI311xp33_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_941), .A3(n_942), .B(n_946), .C(n_954), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_941), .B(n_957), .Y(n_973) );
OAI211xp5_ASAP7_75t_L g1013 ( .A1(n_942), .A2(n_1014), .B(n_1023), .C(n_1033), .Y(n_1013) );
INVx3_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_943), .B(n_950), .Y(n_949) );
INVx3_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g1048 ( .A(n_944), .B(n_1049), .Y(n_1048) );
INVx3_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_952), .B(n_993), .Y(n_1040) );
AOI21xp33_ASAP7_75t_L g1050 ( .A1(n_955), .A2(n_1003), .B(n_1051), .Y(n_1050) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_956), .B(n_957), .Y(n_955) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_960), .B(n_963), .Y(n_959) );
INVx1_ASAP7_75t_L g960 ( .A(n_961), .Y(n_960) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
NAND5xp2_ASAP7_75t_L g965 ( .A(n_966), .B(n_974), .C(n_979), .D(n_991), .E(n_995), .Y(n_965) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_978), .B(n_1048), .Y(n_1047) );
A2O1A1Ixp33_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_985), .B(n_986), .C(n_990), .Y(n_979) );
INVx1_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
INVx1_ASAP7_75t_L g1022 ( .A(n_987), .Y(n_1022) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1001 ( .A(n_990), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_992), .B(n_994), .Y(n_991) );
INVx1_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_993), .B(n_1029), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_1001), .B1(n_1002), .B2(n_1004), .C(n_1006), .Y(n_995) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
CKINVDCx14_ASAP7_75t_R g1007 ( .A(n_1008), .Y(n_1007) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
INVxp67_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1044), .B1(n_1045), .B2(n_1047), .C(n_1050), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_1053), .Y(n_1052) );
INVxp67_ASAP7_75t_SL g1054 ( .A(n_1055), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_1058), .Y(n_1057) );
XNOR2xp5_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .Y(n_1058) );
NOR2xp67_ASAP7_75t_L g1060 ( .A(n_1061), .B(n_1069), .Y(n_1060) );
NAND4xp25_ASAP7_75t_L g1061 ( .A(n_1062), .B(n_1064), .C(n_1065), .D(n_1066), .Y(n_1061) );
NAND4xp25_ASAP7_75t_SL g1069 ( .A(n_1070), .B(n_1071), .C(n_1072), .D(n_1074), .Y(n_1069) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
HB1xp67_ASAP7_75t_L g1083 ( .A(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NAND2xp5_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1102), .Y(n_1085) );
NOR3xp33_ASAP7_75t_SL g1086 ( .A(n_1087), .B(n_1092), .C(n_1097), .Y(n_1086) );
OAI22xp5_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1089), .B1(n_1090), .B2(n_1091), .Y(n_1087) );
OAI22xp5_ASAP7_75t_L g1092 ( .A1(n_1093), .A2(n_1094), .B1(n_1095), .B2(n_1096), .Y(n_1092) );
OAI21xp33_ASAP7_75t_L g1097 ( .A1(n_1098), .A2(n_1099), .B(n_1100), .Y(n_1097) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1106), .Y(n_1102) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1105), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
HB1xp67_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g1114 ( .A(n_1115), .Y(n_1114) );
endmodule