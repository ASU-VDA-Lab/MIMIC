module fake_netlist_5_1169_n_715 (n_137, n_91, n_82, n_122, n_10, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_715);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_715;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_139;
wire n_280;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_606;
wire n_640;
wire n_275;
wire n_559;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_692;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_570;
wire n_457;
wire n_514;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_140;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_691;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_50),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_125),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_73),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_64),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_2),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_62),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_35),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_95),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_34),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_10),
.Y(n_156)
);

BUFx2_ASAP7_75t_SL g157 ( 
.A(n_28),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_14),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_60),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_54),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_29),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_6),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_69),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_8),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_101),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_74),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_84),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_99),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_63),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_87),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_137),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_102),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_21),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_116),
.B(n_58),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_133),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_72),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_71),
.Y(n_190)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_174),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_147),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_0),
.Y(n_196)
);

OAI21x1_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_59),
.B(n_138),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_0),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_143),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_166),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_156),
.B(n_3),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_155),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_187),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_141),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_170),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_139),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

OAI22x1_ASAP7_75t_L g218 ( 
.A1(n_178),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_218)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_148),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_139),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_153),
.B(n_15),
.Y(n_226)
);

CKINVDCx11_ASAP7_75t_R g227 ( 
.A(n_140),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_218),
.B(n_140),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_216),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_227),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_224),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_160),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_208),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_192),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_206),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_R g248 ( 
.A(n_210),
.B(n_152),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_161),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_200),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_222),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_222),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_163),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_190),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_222),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVxp33_ASAP7_75t_SL g261 ( 
.A(n_205),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_212),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_201),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_226),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

NOR3xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_198),
.C(n_196),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_243),
.B(n_173),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_199),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_246),
.B(n_185),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_223),
.Y(n_276)
);

AO221x1_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_204),
.B1(n_209),
.B2(n_203),
.C(n_202),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_264),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_235),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_240),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_213),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_262),
.Y(n_283)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_260),
.Y(n_284)
);

NOR3xp33_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_223),
.C(n_213),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_237),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_199),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_261),
.B(n_226),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_199),
.Y(n_292)
);

OR2x6_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_203),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_242),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_256),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_263),
.B(n_219),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_246),
.B(n_219),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_191),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_252),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_234),
.Y(n_302)
);

BUFx6f_ASAP7_75t_SL g303 ( 
.A(n_231),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_247),
.B(n_219),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_257),
.B(n_191),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_242),
.B(n_191),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_233),
.Y(n_308)
);

BUFx6f_ASAP7_75t_SL g309 ( 
.A(n_230),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_255),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_165),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_238),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_236),
.B(n_191),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_L g315 ( 
.A(n_239),
.B(n_228),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_260),
.B(n_195),
.Y(n_316)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_260),
.Y(n_317)
);

AOI221xp5_ASAP7_75t_L g318 ( 
.A1(n_250),
.A2(n_195),
.B1(n_182),
.B2(n_181),
.C(n_188),
.Y(n_318)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_235),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_241),
.B(n_207),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_284),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_271),
.A2(n_207),
.B1(n_194),
.B2(n_197),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_194),
.Y(n_325)
);

INVx6_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_311),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_317),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_194),
.B1(n_186),
.B2(n_179),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_287),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_295),
.A2(n_176),
.B1(n_171),
.B2(n_167),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_311),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_311),
.Y(n_334)
);

AND2x4_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_16),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

INVx6_ASAP7_75t_L g337 ( 
.A(n_293),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_5),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_319),
.B(n_7),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_17),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_283),
.B(n_8),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_281),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_18),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_19),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_20),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_294),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_269),
.B(n_22),
.Y(n_347)
);

AOI22xp33_ASAP7_75t_L g348 ( 
.A1(n_277),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_319),
.B(n_9),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_290),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_309),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_279),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_13),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_282),
.B(n_23),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_288),
.Y(n_358)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_313),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_294),
.B(n_24),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_286),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_270),
.B(n_25),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_270),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

AND2x4_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_26),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_299),
.B(n_30),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_273),
.B(n_31),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_301),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_296),
.B(n_32),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_272),
.B(n_33),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_286),
.B(n_36),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_286),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_297),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_315),
.B(n_40),
.Y(n_377)
);

O2A1O1Ixp5_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_44),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_275),
.B(n_45),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_347),
.A2(n_304),
.B(n_312),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_331),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_341),
.B(n_315),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_357),
.B1(n_356),
.B2(n_347),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_358),
.B(n_46),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

NAND3xp33_ASAP7_75t_SL g390 ( 
.A(n_350),
.B(n_303),
.C(n_309),
.Y(n_390)
);

BUFx8_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

OAI22x1_ASAP7_75t_L g393 ( 
.A1(n_328),
.A2(n_303),
.B1(n_48),
.B2(n_49),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_323),
.A2(n_47),
.B(n_51),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_52),
.B(n_53),
.C(n_55),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_327),
.A2(n_56),
.B(n_61),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

BUFx8_ASAP7_75t_L g400 ( 
.A(n_359),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_333),
.A2(n_65),
.B(n_66),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_371),
.B(n_68),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_335),
.B(n_70),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_376),
.Y(n_404)
);

NOR2xp67_ASAP7_75t_SL g405 ( 
.A(n_380),
.B(n_75),
.Y(n_405)
);

INVx2_ASAP7_75t_SL g406 ( 
.A(n_326),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_335),
.B(n_77),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_78),
.B(n_79),
.C(n_80),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_332),
.B(n_81),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_82),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_83),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_85),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_337),
.B(n_340),
.Y(n_414)
);

OR2x6_ASAP7_75t_L g415 ( 
.A(n_337),
.B(n_88),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_334),
.A2(n_89),
.B(n_92),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_353),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_345),
.B(n_98),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_340),
.B(n_100),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_339),
.B(n_103),
.Y(n_420)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_366),
.B(n_106),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_352),
.Y(n_422)
);

NOR3xp33_ASAP7_75t_SL g423 ( 
.A(n_373),
.B(n_107),
.C(n_109),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_336),
.A2(n_110),
.B(n_111),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_363),
.A2(n_112),
.B(n_113),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_114),
.Y(n_426)
);

O2A1O1Ixp33_ASAP7_75t_L g427 ( 
.A1(n_348),
.A2(n_117),
.B(n_120),
.C(n_121),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_363),
.A2(n_122),
.B(n_123),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

OAI21x1_ASAP7_75t_L g431 ( 
.A1(n_426),
.A2(n_374),
.B(n_360),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_366),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_372),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_389),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_403),
.A2(n_362),
.B(n_374),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g438 ( 
.A1(n_411),
.A2(n_360),
.B(n_402),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_385),
.Y(n_439)
);

BUFx2_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_385),
.Y(n_441)
);

CKINVDCx11_ASAP7_75t_R g442 ( 
.A(n_415),
.Y(n_442)
);

BUFx12f_ASAP7_75t_L g443 ( 
.A(n_391),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_383),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_384),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_387),
.A2(n_324),
.B(n_378),
.Y(n_449)
);

INVx2_ASAP7_75t_SL g450 ( 
.A(n_399),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_410),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_382),
.A2(n_344),
.B(n_343),
.Y(n_452)
);

AO21x2_ASAP7_75t_L g453 ( 
.A1(n_386),
.A2(n_325),
.B(n_367),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_407),
.A2(n_344),
.B(n_367),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_404),
.Y(n_455)
);

BUFx2_ASAP7_75t_SL g456 ( 
.A(n_404),
.Y(n_456)
);

NAND2x1p5_ASAP7_75t_L g457 ( 
.A(n_405),
.B(n_377),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_415),
.Y(n_459)
);

CKINVDCx6p67_ASAP7_75t_R g460 ( 
.A(n_393),
.Y(n_460)
);

AO21x2_ASAP7_75t_L g461 ( 
.A1(n_418),
.A2(n_379),
.B(n_355),
.Y(n_461)
);

BUFx5_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_422),
.Y(n_463)
);

AO21x2_ASAP7_75t_L g464 ( 
.A1(n_396),
.A2(n_365),
.B(n_377),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_429),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_425),
.A2(n_375),
.B(n_329),
.Y(n_466)
);

INVx1_ASAP7_75t_SL g467 ( 
.A(n_392),
.Y(n_467)
);

AND2x4_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_406),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_388),
.Y(n_469)
);

AO21x2_ASAP7_75t_L g470 ( 
.A1(n_423),
.A2(n_362),
.B(n_128),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_413),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_428),
.A2(n_124),
.B(n_129),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_463),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_460),
.A2(n_409),
.B1(n_420),
.B2(n_390),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_444),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_448),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_451),
.Y(n_478)
);

BUFx6f_ASAP7_75t_SL g479 ( 
.A(n_436),
.Y(n_479)
);

BUFx12f_ASAP7_75t_L g480 ( 
.A(n_443),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_436),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_447),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_449),
.A2(n_408),
.B(n_424),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_443),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

OR2x6_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_417),
.Y(n_486)
);

OR2x6_ASAP7_75t_L g487 ( 
.A(n_434),
.B(n_427),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_437),
.A2(n_416),
.B(n_401),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_442),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_462),
.B(n_397),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_465),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_465),
.Y(n_492)
);

INVx6_ASAP7_75t_L g493 ( 
.A(n_455),
.Y(n_493)
);

BUFx8_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

INVx6_ASAP7_75t_L g496 ( 
.A(n_455),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_430),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_445),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_439),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_445),
.Y(n_500)
);

OAI22xp33_ASAP7_75t_L g501 ( 
.A1(n_460),
.A2(n_394),
.B1(n_131),
.B2(n_132),
.Y(n_501)
);

CKINVDCx11_ASAP7_75t_R g502 ( 
.A(n_435),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_440),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_469),
.A2(n_130),
.B1(n_134),
.B2(n_136),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_434),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_439),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_435),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_467),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_432),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_477),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_493),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_R g514 ( 
.A(n_484),
.B(n_434),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_509),
.Y(n_515)
);

OA21x2_ASAP7_75t_L g516 ( 
.A1(n_488),
.A2(n_452),
.B(n_431),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_474),
.A2(n_471),
.B1(n_459),
.B2(n_457),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_474),
.A2(n_468),
.B1(n_442),
.B2(n_462),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_475),
.Y(n_519)
);

NAND2x1p5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_439),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_476),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_477),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_502),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_509),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_487),
.A2(n_468),
.B1(n_462),
.B2(n_470),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

NAND2xp33_ASAP7_75t_R g527 ( 
.A(n_486),
.B(n_468),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_R g528 ( 
.A(n_486),
.B(n_433),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g529 ( 
.A(n_480),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_505),
.B(n_458),
.Y(n_530)
);

OAI21xp33_ASAP7_75t_SL g531 ( 
.A1(n_506),
.A2(n_466),
.B(n_454),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_491),
.Y(n_532)
);

OR2x6_ASAP7_75t_L g533 ( 
.A(n_487),
.B(n_457),
.Y(n_533)
);

OR2x6_ASAP7_75t_L g534 ( 
.A(n_487),
.B(n_457),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_502),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_478),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_491),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_481),
.B(n_447),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_490),
.A2(n_466),
.B(n_472),
.Y(n_539)
);

INVx4_ASAP7_75t_R g540 ( 
.A(n_510),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_481),
.B(n_458),
.Y(n_541)
);

NOR3xp33_ASAP7_75t_SL g542 ( 
.A(n_501),
.B(n_441),
.C(n_450),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_492),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_473),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_493),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_501),
.A2(n_462),
.B1(n_470),
.B2(n_464),
.Y(n_547)
);

NAND2xp33_ASAP7_75t_R g548 ( 
.A(n_486),
.B(n_433),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_R g549 ( 
.A(n_485),
.B(n_433),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_494),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_504),
.B(n_462),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_498),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_488),
.A2(n_452),
.B(n_472),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_500),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_R g556 ( 
.A(n_479),
.B(n_439),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_519),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_512),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_495),
.Y(n_559)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_461),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_552),
.B(n_508),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_554),
.A2(n_431),
.B(n_438),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_538),
.B(n_462),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_521),
.B(n_508),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_522),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_532),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_536),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_537),
.B(n_545),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_553),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_518),
.A2(n_506),
.B1(n_462),
.B2(n_489),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_555),
.B(n_503),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_549),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_511),
.B(n_503),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_551),
.Y(n_575)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_530),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_533),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_533),
.B(n_534),
.Y(n_579)
);

INVx5_ASAP7_75t_SL g580 ( 
.A(n_533),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_539),
.B(n_461),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_534),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_534),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_517),
.B(n_482),
.Y(n_585)
);

OAI22xp33_ASAP7_75t_L g586 ( 
.A1(n_527),
.A2(n_450),
.B1(n_496),
.B2(n_493),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_513),
.B(n_446),
.Y(n_588)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_539),
.Y(n_589)
);

OAI221xp5_ASAP7_75t_L g590 ( 
.A1(n_542),
.A2(n_547),
.B1(n_525),
.B2(n_531),
.C(n_528),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_520),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_513),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_573),
.B(n_515),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_589),
.B(n_547),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_524),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_546),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_531),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_560),
.Y(n_600)
);

OAI21xp33_ASAP7_75t_L g601 ( 
.A1(n_590),
.A2(n_535),
.B(n_523),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_461),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_569),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_560),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_579),
.Y(n_605)
);

BUFx2_ASAP7_75t_L g606 ( 
.A(n_572),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_569),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_546),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_587),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_579),
.B(n_550),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_568),
.B(n_526),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_568),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_585),
.B(n_529),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_574),
.B(n_520),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_582),
.B(n_483),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_583),
.B(n_578),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_586),
.B(n_570),
.Y(n_617)
);

NAND3xp33_ASAP7_75t_L g618 ( 
.A(n_584),
.B(n_548),
.C(n_514),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_563),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_583),
.B(n_591),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_595),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_596),
.B(n_606),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_619),
.B(n_600),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_599),
.B(n_580),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_599),
.B(n_580),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_612),
.B(n_564),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_598),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_603),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_610),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_580),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_610),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_600),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_603),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_620),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_607),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_607),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_604),
.B(n_580),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_622),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_636),
.Y(n_639)
);

OAI32xp33_ASAP7_75t_L g640 ( 
.A1(n_623),
.A2(n_613),
.A3(n_617),
.B1(n_601),
.B2(n_618),
.Y(n_640)
);

NOR2x1p5_ASAP7_75t_SL g641 ( 
.A(n_637),
.B(n_581),
.Y(n_641)
);

OAI22xp33_ASAP7_75t_L g642 ( 
.A1(n_629),
.A2(n_617),
.B1(n_605),
.B2(n_594),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_636),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_629),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_628),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_633),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_631),
.B(n_620),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_632),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_640),
.B(n_610),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_642),
.A2(n_594),
.B1(n_605),
.B2(n_631),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_638),
.A2(n_605),
.B1(n_629),
.B2(n_593),
.Y(n_651)
);

AOI211xp5_ASAP7_75t_SL g652 ( 
.A1(n_647),
.A2(n_625),
.B(n_624),
.C(n_609),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_648),
.Y(n_653)
);

NAND2x1p5_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_648),
.Y(n_654)
);

AOI21xp33_ASAP7_75t_SL g655 ( 
.A1(n_649),
.A2(n_611),
.B(n_644),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_650),
.Y(n_656)
);

OAI22xp33_ASAP7_75t_L g657 ( 
.A1(n_652),
.A2(n_629),
.B1(n_634),
.B2(n_626),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_651),
.B(n_621),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_657),
.B(n_647),
.Y(n_659)
);

NAND4xp25_ASAP7_75t_L g660 ( 
.A(n_658),
.B(n_608),
.C(n_577),
.D(n_592),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_655),
.B(n_656),
.Y(n_661)
);

NOR2xp67_ASAP7_75t_L g662 ( 
.A(n_654),
.B(n_646),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_661),
.B(n_592),
.C(n_627),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_662),
.A2(n_659),
.B1(n_625),
.B2(n_624),
.Y(n_664)
);

O2A1O1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_660),
.A2(n_645),
.B(n_632),
.C(n_639),
.Y(n_665)
);

AOI321xp33_ASAP7_75t_L g666 ( 
.A1(n_664),
.A2(n_597),
.A3(n_574),
.B1(n_630),
.B2(n_615),
.C(n_620),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_663),
.B(n_665),
.Y(n_667)
);

NOR4xp25_ASAP7_75t_L g668 ( 
.A(n_664),
.B(n_540),
.C(n_643),
.D(n_635),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_663),
.B(n_641),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_667),
.Y(n_670)
);

AND2x4_ASAP7_75t_L g671 ( 
.A(n_669),
.B(n_634),
.Y(n_671)
);

NOR2x1_ASAP7_75t_L g672 ( 
.A(n_668),
.B(n_446),
.Y(n_672)
);

NOR2x1_ASAP7_75t_L g673 ( 
.A(n_666),
.B(n_446),
.Y(n_673)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_667),
.A2(n_597),
.B1(n_479),
.B2(n_630),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_669),
.Y(n_676)
);

INVx1_ASAP7_75t_SL g677 ( 
.A(n_670),
.Y(n_677)
);

NAND4xp25_ASAP7_75t_L g678 ( 
.A(n_675),
.B(n_597),
.C(n_616),
.D(n_614),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_676),
.B(n_564),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_671),
.Y(n_680)
);

NAND3x2_ASAP7_75t_L g681 ( 
.A(n_672),
.B(n_674),
.C(n_673),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_670),
.B(n_556),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_672),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_676),
.B(n_588),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_677),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_680),
.B(n_561),
.Y(n_686)
);

HB1xp67_ASAP7_75t_L g687 ( 
.A(n_683),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_682),
.B(n_588),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

NAND4xp25_ASAP7_75t_SL g690 ( 
.A(n_681),
.B(n_602),
.C(n_591),
.D(n_561),
.Y(n_690)
);

NOR3xp33_ASAP7_75t_L g691 ( 
.A(n_678),
.B(n_588),
.C(n_571),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_684),
.Y(n_692)
);

NOR2x1_ASAP7_75t_L g693 ( 
.A(n_685),
.B(n_692),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_687),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_690),
.A2(n_684),
.B1(n_571),
.B2(n_602),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_686),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_689),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_691),
.Y(n_699)
);

AOI22xp5_ASAP7_75t_L g700 ( 
.A1(n_693),
.A2(n_499),
.B1(n_496),
.B2(n_446),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_694),
.B(n_559),
.Y(n_701)
);

BUFx2_ASAP7_75t_L g702 ( 
.A(n_698),
.Y(n_702)
);

AOI211xp5_ASAP7_75t_SL g703 ( 
.A1(n_697),
.A2(n_446),
.B(n_496),
.C(n_559),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_699),
.Y(n_704)
);

OAI31xp33_ASAP7_75t_SL g705 ( 
.A1(n_696),
.A2(n_566),
.A3(n_565),
.B(n_558),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_702),
.Y(n_706)
);

XOR2xp5_ASAP7_75t_L g707 ( 
.A(n_704),
.B(n_700),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_701),
.Y(n_708)
);

OA22x2_ASAP7_75t_L g709 ( 
.A1(n_706),
.A2(n_695),
.B1(n_703),
.B2(n_705),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_708),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_707),
.A2(n_499),
.B1(n_470),
.B2(n_483),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_710),
.A2(n_499),
.B1(n_566),
.B2(n_565),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_709),
.B1(n_711),
.B2(n_453),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_713),
.B(n_438),
.Y(n_714)
);

AOI211xp5_ASAP7_75t_L g715 ( 
.A1(n_714),
.A2(n_558),
.B(n_453),
.C(n_562),
.Y(n_715)
);


endmodule