module real_jpeg_28451_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_19),
.Y(n_41)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_0),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_1),
.A2(n_19),
.B1(n_21),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_39),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_32),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_3),
.A2(n_50),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_3),
.A2(n_24),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_24),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_40),
.B1(n_103),
.B2(n_107),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_4),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_5),
.A2(n_19),
.B1(n_21),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_5),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_19),
.B1(n_21),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_6),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_18)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_7),
.A2(n_21),
.A3(n_24),
.B1(n_88),
.B2(n_89),
.Y(n_87)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_11),
.A2(n_27),
.B1(n_50),
.B2(n_51),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_11),
.A2(n_19),
.B1(n_21),
.B2(n_27),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_79),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_77),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_45),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_15),
.B(n_45),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_30),
.C(n_37),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_16),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_26),
.B2(n_28),
.Y(n_16)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_17),
.A2(n_18),
.B1(n_26),
.B2(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_23),
.Y(n_17)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_18),
.B(n_56),
.Y(n_104)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_19),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_19),
.B(n_109),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_25),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_24),
.B(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_25),
.A2(n_34),
.A3(n_50),
.B1(n_55),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_48)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_36),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_37),
.B(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_38),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_42),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_40),
.A2(n_44),
.B1(n_97),
.B2(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_41),
.A2(n_71),
.B1(n_96),
.B2(n_98),
.Y(n_95)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_44),
.B(n_56),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_65),
.B1(n_75),
.B2(n_76),
.Y(n_45)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_65),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.Y(n_65)
);

INVx5_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_93),
.B(n_112),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_90),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_99)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_85),
.Y(n_88)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_100),
.B(n_111),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_99),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_105),
.B(n_110),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);


endmodule