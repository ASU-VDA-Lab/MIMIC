module fake_netlist_1_3074_n_671 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_671);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_90;
wire n_245;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_515;
wire n_253;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_65), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_61), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_55), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_17), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_40), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_48), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_25), .Y(n_85) );
BUFx3_ASAP7_75t_L g86 ( .A(n_74), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_69), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_58), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_11), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_18), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_70), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_4), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_13), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_75), .Y(n_97) );
INVxp67_ASAP7_75t_SL g98 ( .A(n_29), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_11), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_13), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_64), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_46), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_14), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_21), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_38), .Y(n_106) );
BUFx3_ASAP7_75t_L g107 ( .A(n_34), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_27), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_6), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_60), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_18), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_14), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVxp67_ASAP7_75t_SL g114 ( .A(n_20), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_45), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_52), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_37), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_22), .Y(n_119) );
BUFx3_ASAP7_75t_L g120 ( .A(n_71), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_16), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_10), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_54), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_107), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_77), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_107), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_80), .B(n_0), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_90), .B(n_0), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_84), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_77), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_84), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_111), .B(n_1), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_79), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_81), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_111), .B(n_2), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_82), .B(n_2), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_90), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_120), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_100), .B(n_3), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_100), .B(n_3), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_120), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_83), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_97), .Y(n_147) );
AND2x2_ASAP7_75t_L g148 ( .A(n_89), .B(n_4), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_99), .B(n_5), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_89), .B(n_5), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_83), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_104), .B(n_109), .Y(n_152) );
AND2x4_ASAP7_75t_L g153 ( .A(n_95), .B(n_6), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_85), .Y(n_154) );
CKINVDCx6p67_ASAP7_75t_R g155 ( .A(n_85), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_112), .B(n_7), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_88), .Y(n_157) );
HB1xp67_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_78), .B(n_7), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_96), .B(n_8), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_88), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_91), .B(n_92), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_91), .Y(n_163) );
HB1xp67_ASAP7_75t_L g164 ( .A(n_96), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_113), .B(n_8), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_124), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_155), .B(n_87), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_124), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_127), .B(n_87), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_127), .B(n_117), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_160), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_155), .B(n_117), .Y(n_173) );
BUFx2_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
OAI221xp5_ASAP7_75t_L g175 ( .A1(n_158), .A2(n_122), .B1(n_121), .B2(n_118), .C(n_101), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_132), .B(n_93), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_132), .B(n_93), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_135), .B(n_118), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_124), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_135), .B(n_122), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_164), .B(n_121), .Y(n_183) );
CKINVDCx8_ASAP7_75t_R g184 ( .A(n_135), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_147), .Y(n_185) );
OR2x2_ASAP7_75t_L g186 ( .A(n_130), .B(n_123), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_139), .B(n_123), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_152), .B(n_110), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_146), .Y(n_189) );
AND2x2_ASAP7_75t_SL g190 ( .A(n_135), .B(n_119), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_134), .B(n_105), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_146), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_138), .B(n_119), .Y(n_193) );
AND2x6_ASAP7_75t_L g194 ( .A(n_138), .B(n_92), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_160), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_139), .B(n_94), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_160), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_124), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_134), .B(n_116), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_143), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_136), .B(n_94), .Y(n_201) );
INVxp33_ASAP7_75t_SL g202 ( .A(n_144), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_136), .B(n_114), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_154), .Y(n_205) );
BUFx2_ASAP7_75t_L g206 ( .A(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_137), .B(n_108), .Y(n_207) );
INVx2_ASAP7_75t_SL g208 ( .A(n_162), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_124), .Y(n_209) );
INVx4_ASAP7_75t_SL g210 ( .A(n_162), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_138), .B(n_115), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_125), .Y(n_212) );
AO22x2_ASAP7_75t_L g213 ( .A1(n_160), .A2(n_106), .B1(n_103), .B2(n_102), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_137), .B(n_98), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_140), .B(n_42), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_154), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_140), .B(n_9), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_154), .Y(n_218) );
BUFx3_ASAP7_75t_L g219 ( .A(n_125), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_161), .B(n_9), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_161), .B(n_12), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_163), .B(n_15), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_125), .Y(n_223) );
BUFx3_ASAP7_75t_L g224 ( .A(n_125), .Y(n_224) );
AND2x6_ASAP7_75t_SL g225 ( .A(n_183), .B(n_153), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_190), .B(n_153), .Y(n_226) );
CKINVDCx11_ASAP7_75t_R g227 ( .A(n_174), .Y(n_227) );
CKINVDCx16_ASAP7_75t_R g228 ( .A(n_174), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_192), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_192), .Y(n_230) );
BUFx3_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_202), .B(n_163), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_171), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_192), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_184), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_188), .B(n_162), .Y(n_236) );
BUFx3_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_192), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_192), .Y(n_239) );
AND2x4_ASAP7_75t_L g240 ( .A(n_179), .B(n_153), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_177), .B(n_162), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_205), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_171), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_171), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_205), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
BUFx12f_ASAP7_75t_L g247 ( .A(n_185), .Y(n_247) );
AND3x2_ASAP7_75t_SL g248 ( .A(n_213), .B(n_151), .C(n_157), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_205), .Y(n_249) );
BUFx6f_ASAP7_75t_L g250 ( .A(n_198), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_178), .B(n_162), .Y(n_251) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_184), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_205), .Y(n_253) );
BUFx6f_ASAP7_75t_L g254 ( .A(n_198), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_203), .B(n_162), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_187), .B(n_148), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_190), .A2(n_148), .B1(n_150), .B2(n_162), .Y(n_257) );
BUFx3_ASAP7_75t_L g258 ( .A(n_194), .Y(n_258) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_212), .Y(n_259) );
BUFx2_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_203), .B(n_150), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_186), .B(n_151), .Y(n_262) );
INVx2_ASAP7_75t_SL g263 ( .A(n_190), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_167), .Y(n_264) );
INVx2_ASAP7_75t_SL g265 ( .A(n_179), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_195), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_195), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_186), .B(n_157), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_212), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_187), .B(n_129), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_195), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_196), .B(n_159), .Y(n_272) );
BUFx12f_ASAP7_75t_L g273 ( .A(n_185), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_205), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_218), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_197), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_156), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_183), .B(n_165), .Y(n_278) );
BUFx3_ASAP7_75t_L g279 ( .A(n_194), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_197), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_194), .A2(n_149), .B1(n_154), .B2(n_131), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_201), .B(n_133), .Y(n_283) );
AND2x6_ASAP7_75t_L g284 ( .A(n_193), .B(n_145), .Y(n_284) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_179), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_201), .B(n_133), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_231), .Y(n_288) );
BUFx12f_ASAP7_75t_L g289 ( .A(n_227), .Y(n_289) );
INVx2_ASAP7_75t_SL g290 ( .A(n_231), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_233), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_278), .B(n_200), .Y(n_292) );
BUFx2_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_233), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g295 ( .A1(n_226), .A2(n_213), .B1(n_194), .B2(n_206), .Y(n_295) );
OAI22xp5_ASAP7_75t_L g296 ( .A1(n_257), .A2(n_206), .B1(n_193), .B2(n_213), .Y(n_296) );
AOI22x1_ASAP7_75t_L g297 ( .A1(n_234), .A2(n_213), .B1(n_223), .B2(n_166), .Y(n_297) );
INVx3_ASAP7_75t_L g298 ( .A(n_237), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_243), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_243), .Y(n_300) );
BUFx4_ASAP7_75t_SL g301 ( .A(n_225), .Y(n_301) );
OAI222xp33_ASAP7_75t_L g302 ( .A1(n_228), .A2(n_175), .B1(n_179), .B2(n_182), .C1(n_222), .C2(n_193), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_237), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_228), .Y(n_304) );
NOR2x1_ASAP7_75t_L g305 ( .A(n_237), .B(n_217), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_244), .Y(n_306) );
INVx1_ASAP7_75t_SL g307 ( .A(n_282), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_244), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_258), .B(n_197), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_257), .A2(n_193), .B1(n_211), .B2(n_182), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_262), .Y(n_311) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_263), .A2(n_182), .B1(n_211), .B2(n_222), .Y(n_312) );
INVxp67_ASAP7_75t_L g313 ( .A(n_232), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_264), .B(n_173), .Y(n_314) );
NAND2x1_ASAP7_75t_L g315 ( .A(n_284), .B(n_182), .Y(n_315) );
BUFx6f_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_263), .A2(n_211), .B1(n_170), .B2(n_169), .Y(n_317) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_247), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_266), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_278), .B(n_214), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_266), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_256), .B(n_211), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_SL g323 ( .A1(n_241), .A2(n_220), .B(n_221), .C(n_199), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_268), .B(n_191), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_267), .Y(n_325) );
INVx5_ASAP7_75t_L g326 ( .A(n_284), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_247), .Y(n_327) );
BUFx3_ASAP7_75t_L g328 ( .A(n_258), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_267), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_256), .B(n_207), .Y(n_330) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_271), .A2(n_215), .B(n_224), .C(n_219), .Y(n_331) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_235), .Y(n_332) );
NAND2xp33_ASAP7_75t_L g333 ( .A(n_265), .B(n_208), .Y(n_333) );
INVx4_ASAP7_75t_L g334 ( .A(n_279), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_279), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_240), .A2(n_125), .B1(n_126), .B2(n_128), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_311), .B(n_277), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_307), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_292), .A2(n_240), .B1(n_286), .B2(n_265), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_324), .A2(n_240), .B(n_286), .C(n_255), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_292), .B(n_283), .Y(n_341) );
BUFx2_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_326), .Y(n_343) );
INVxp67_ASAP7_75t_SL g344 ( .A(n_310), .Y(n_344) );
OA21x2_ASAP7_75t_L g345 ( .A1(n_331), .A2(n_181), .B(n_223), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_294), .Y(n_346) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_289), .A2(n_273), .B1(n_252), .B2(n_248), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_313), .A2(n_273), .B1(n_279), .B2(n_270), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_316), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_291), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_296), .A2(n_240), .B1(n_270), .B2(n_260), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g352 ( .A1(n_320), .A2(n_260), .B1(n_280), .B2(n_271), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_295), .A2(n_248), .B1(n_287), .B2(n_283), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_320), .A2(n_280), .B1(n_276), .B2(n_261), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_291), .Y(n_355) );
O2A1O1Ixp33_ASAP7_75t_SL g356 ( .A1(n_315), .A2(n_251), .B(n_276), .C(n_236), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_323), .A2(n_272), .B(n_208), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_300), .Y(n_358) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_295), .A2(n_248), .B1(n_281), .B2(n_126), .Y(n_359) );
O2A1O1Ixp33_ASAP7_75t_L g360 ( .A1(n_302), .A2(n_172), .B(n_176), .C(n_180), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_326), .Y(n_361) );
AND2x4_ASAP7_75t_L g362 ( .A(n_322), .B(n_284), .Y(n_362) );
OAI221xp5_ASAP7_75t_L g363 ( .A1(n_314), .A2(n_225), .B1(n_219), .B2(n_224), .C(n_254), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_294), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_299), .Y(n_365) );
OAI22xp33_ASAP7_75t_L g366 ( .A1(n_289), .A2(n_285), .B1(n_246), .B2(n_269), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_300), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g368 ( .A1(n_344), .A2(n_308), .B1(n_306), .B2(n_319), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_340), .A2(n_312), .B(n_330), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_337), .B(n_332), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_338), .B(n_318), .Y(n_372) );
AOI322xp5_ASAP7_75t_L g373 ( .A1(n_341), .A2(n_327), .A3(n_318), .B1(n_322), .B2(n_301), .C1(n_317), .C2(n_315), .Y(n_373) );
AOI21xp5_ASAP7_75t_L g374 ( .A1(n_356), .A2(n_308), .B(n_319), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_321), .B1(n_306), .B2(n_325), .C(n_299), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_357), .A2(n_321), .B(n_297), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_338), .B(n_325), .Y(n_377) );
AOI221xp5_ASAP7_75t_SL g378 ( .A1(n_348), .A2(n_329), .B1(n_145), .B2(n_126), .C(n_142), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_353), .A2(n_329), .B1(n_297), .B2(n_305), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_351), .A2(n_293), .B1(n_309), .B2(n_303), .Y(n_380) );
AOI222xp33_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_284), .B1(n_293), .B2(n_326), .C1(n_305), .C2(n_334), .Y(n_381) );
AOI221xp5_ASAP7_75t_L g382 ( .A1(n_339), .A2(n_336), .B1(n_145), .B2(n_142), .C(n_128), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_347), .A2(n_284), .B1(n_126), .B2(n_128), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_342), .B(n_309), .Y(n_384) );
NOR2xp33_ASAP7_75t_R g385 ( .A(n_343), .B(n_326), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_359), .A2(n_309), .B1(n_328), .B2(n_303), .Y(n_386) );
BUFx3_ASAP7_75t_L g387 ( .A(n_346), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_359), .A2(n_284), .B1(n_128), .B2(n_142), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_346), .Y(n_389) );
INVx3_ASAP7_75t_L g390 ( .A(n_343), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g391 ( .A1(n_354), .A2(n_336), .B1(n_290), .B2(n_334), .C(n_288), .Y(n_391) );
AND2x6_ASAP7_75t_L g392 ( .A(n_346), .B(n_303), .Y(n_392) );
OAI211xp5_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_326), .B(n_128), .C(n_126), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_362), .A2(n_284), .B1(n_290), .B2(n_334), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_389), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_370), .A2(n_352), .B1(n_350), .B2(n_358), .C(n_355), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_377), .B(n_364), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_371), .A2(n_367), .B1(n_358), .B2(n_350), .C(n_355), .Y(n_398) );
OAI31xp33_ASAP7_75t_L g399 ( .A1(n_380), .A2(n_366), .A3(n_362), .B(n_367), .Y(n_399) );
INVx4_ASAP7_75t_SL g400 ( .A(n_392), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_384), .B(n_365), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_365), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_373), .B(n_145), .C(n_142), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_368), .B(n_365), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_375), .A2(n_364), .B(n_343), .C(n_360), .Y(n_405) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_383), .A2(n_364), .B(n_345), .C(n_326), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_368), .A2(n_362), .B1(n_361), .B2(n_328), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_372), .B(n_362), .Y(n_409) );
NAND3xp33_ASAP7_75t_SL g410 ( .A(n_383), .B(n_189), .C(n_172), .Y(n_410) );
OAI221xp5_ASAP7_75t_L g411 ( .A1(n_388), .A2(n_361), .B1(n_345), .B2(n_334), .C(n_335), .Y(n_411) );
BUFx3_ASAP7_75t_L g412 ( .A(n_392), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_328), .B1(n_349), .B2(n_316), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_386), .A2(n_316), .B1(n_349), .B2(n_288), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_378), .B(n_349), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_381), .A2(n_345), .B1(n_142), .B2(n_145), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_382), .B(n_345), .C(n_218), .Y(n_417) );
OA21x2_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_181), .B(n_168), .Y(n_418) );
NOR3xp33_ASAP7_75t_L g419 ( .A(n_390), .B(n_166), .C(n_168), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_379), .B(n_218), .C(n_209), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx5_ASAP7_75t_SL g422 ( .A(n_385), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_392), .Y(n_423) );
AOI31xp33_ASAP7_75t_L g424 ( .A1(n_379), .A2(n_15), .A3(n_16), .B(n_17), .Y(n_424) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_392), .A2(n_349), .B1(n_316), .B2(n_288), .Y(n_425) );
INVx4_ASAP7_75t_L g426 ( .A(n_392), .Y(n_426) );
BUFx3_ASAP7_75t_L g427 ( .A(n_394), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_374), .B(n_218), .C(n_209), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_397), .B(n_349), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
OAI31xp33_ASAP7_75t_L g431 ( .A1(n_403), .A2(n_405), .A3(n_399), .B(n_396), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_404), .B(n_349), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_397), .B(n_385), .Y(n_433) );
BUFx3_ASAP7_75t_L g434 ( .A(n_412), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_404), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_426), .B(n_316), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
NOR3xp33_ASAP7_75t_L g438 ( .A(n_424), .B(n_393), .C(n_391), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_401), .B(n_219), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_398), .B(n_224), .C(n_189), .D(n_216), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_400), .B(n_19), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_427), .B(n_180), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_402), .B(n_23), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_418), .Y(n_444) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_395), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_395), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_400), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_418), .Y(n_448) );
AND3x1_ASAP7_75t_L g449 ( .A(n_406), .B(n_288), .C(n_335), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_423), .Y(n_450) );
OAI211xp5_ASAP7_75t_SL g451 ( .A1(n_409), .A2(n_204), .B(n_216), .C(n_176), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_423), .Y(n_452) );
NAND3xp33_ASAP7_75t_SL g453 ( .A(n_416), .B(n_204), .C(n_275), .Y(n_453) );
AND2x4_ASAP7_75t_SL g454 ( .A(n_426), .B(n_335), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_427), .B(n_421), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_426), .B(n_24), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_405), .B(n_285), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
OAI31xp33_ASAP7_75t_SL g460 ( .A1(n_407), .A2(n_408), .A3(n_414), .B(n_420), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_400), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_412), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_416), .B(n_26), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_417), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g465 ( .A1(n_410), .A2(n_218), .B(n_250), .C(n_285), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
OAI31xp33_ASAP7_75t_L g467 ( .A1(n_413), .A2(n_298), .A3(n_275), .B(n_274), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_422), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_422), .B(n_30), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_428), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_422), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_425), .B(n_31), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_419), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_402), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_415), .A2(n_333), .B(n_298), .Y(n_475) );
AOI21xp33_ASAP7_75t_L g476 ( .A1(n_403), .A2(n_254), .B(n_285), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_404), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_435), .B(n_33), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_435), .B(n_36), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_477), .B(n_39), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_430), .B(n_41), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_445), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_477), .B(n_43), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_446), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_446), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_474), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_474), .B(n_44), .Y(n_487) );
AOI222xp33_ASAP7_75t_L g488 ( .A1(n_466), .A2(n_298), .B1(n_285), .B2(n_269), .C1(n_259), .C2(n_254), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_432), .B(n_47), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_455), .B(n_49), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_429), .B(n_50), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_455), .B(n_53), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_462), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_433), .B(n_56), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_429), .B(n_57), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_432), .B(n_59), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_462), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_466), .B(n_62), .Y(n_499) );
OR2x6_ASAP7_75t_L g500 ( .A(n_434), .B(n_269), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_443), .B(n_66), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_438), .A2(n_269), .B1(n_259), .B2(n_254), .Y(n_502) );
NOR3xp33_ASAP7_75t_L g503 ( .A(n_440), .B(n_242), .C(n_274), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_450), .B(n_67), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_443), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_452), .B(n_68), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_461), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_450), .B(n_72), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_450), .B(n_76), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_452), .B(n_246), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_456), .B(n_246), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_434), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_456), .B(n_246), .Y(n_515) );
BUFx2_ASAP7_75t_SL g516 ( .A(n_471), .Y(n_516) );
OAI33xp33_ASAP7_75t_L g517 ( .A1(n_473), .A2(n_275), .A3(n_274), .B1(n_245), .B2(n_234), .B3(n_238), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_442), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_456), .B(n_269), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_447), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_440), .A2(n_245), .B(n_242), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_459), .B(n_259), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_439), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_459), .B(n_259), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_431), .B(n_259), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_437), .B(n_444), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_469), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_437), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_464), .B(n_254), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_441), .B(n_250), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_431), .B(n_250), .Y(n_531) );
OAI211xp5_ASAP7_75t_SL g532 ( .A1(n_473), .A2(n_242), .B(n_245), .C(n_238), .Y(n_532) );
AOI221x1_ASAP7_75t_L g533 ( .A1(n_441), .A2(n_250), .B1(n_246), .B2(n_238), .C(n_234), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g534 ( .A(n_486), .B(n_441), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_528), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_514), .B(n_460), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_482), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_518), .B(n_460), .Y(n_539) );
OAI21xp5_ASAP7_75t_SL g540 ( .A1(n_527), .A2(n_468), .B(n_469), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_523), .A2(n_449), .B1(n_471), .B2(n_463), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_498), .Y(n_542) );
INVxp67_ASAP7_75t_SL g543 ( .A(n_528), .Y(n_543) );
AOI211xp5_ASAP7_75t_SL g544 ( .A1(n_505), .A2(n_441), .B(n_457), .C(n_472), .Y(n_544) );
OR2x2_ASAP7_75t_L g545 ( .A(n_492), .B(n_484), .Y(n_545) );
INVxp33_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_485), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_520), .B(n_439), .Y(n_548) );
NAND2x1_ASAP7_75t_L g549 ( .A(n_500), .B(n_457), .Y(n_549) );
INVx3_ASAP7_75t_L g550 ( .A(n_526), .Y(n_550) );
NAND2x1_ASAP7_75t_L g551 ( .A(n_500), .B(n_472), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_507), .B(n_458), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_510), .Y(n_553) );
AOI32xp33_ASAP7_75t_L g554 ( .A1(n_487), .A2(n_449), .A3(n_463), .B1(n_471), .B2(n_465), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_513), .B(n_491), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_513), .B(n_464), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_526), .B(n_458), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_480), .B(n_444), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_530), .B(n_470), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_491), .B(n_436), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_516), .Y(n_561) );
INVx2_ASAP7_75t_SL g562 ( .A(n_500), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_480), .B(n_444), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_489), .B(n_448), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_529), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_483), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_497), .B(n_436), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_478), .B(n_448), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_478), .B(n_448), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_483), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_497), .B(n_436), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_479), .B(n_437), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_502), .B(n_465), .C(n_467), .D(n_451), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_479), .B(n_470), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_499), .B(n_453), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_483), .Y(n_577) );
OAI22xp5_ASAP7_75t_L g578 ( .A1(n_495), .A2(n_454), .B1(n_475), .B2(n_476), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_512), .B(n_470), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_489), .B(n_467), .Y(n_580) );
NOR3xp33_ASAP7_75t_L g581 ( .A(n_525), .B(n_476), .C(n_229), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_531), .B(n_454), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_536), .B(n_524), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_550), .B(n_512), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g585 ( .A(n_561), .B(n_496), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_545), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_555), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_539), .B(n_524), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g589 ( .A1(n_576), .A2(n_502), .B1(n_490), .B2(n_493), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_537), .B(n_522), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_553), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_538), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_542), .Y(n_593) );
INVxp33_ASAP7_75t_L g594 ( .A(n_549), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_547), .B(n_522), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_550), .B(n_515), .Y(n_596) );
INVx2_ASAP7_75t_SL g597 ( .A(n_550), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_551), .A2(n_517), .B(n_481), .Y(n_598) );
AND3x1_ASAP7_75t_L g599 ( .A(n_544), .B(n_501), .C(n_508), .Y(n_599) );
INVx1_ASAP7_75t_SL g600 ( .A(n_560), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_567), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g602 ( .A1(n_540), .A2(n_530), .B(n_506), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_548), .Y(n_603) );
AO21x1_ASAP7_75t_L g604 ( .A1(n_543), .A2(n_506), .B(n_509), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_557), .B(n_511), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_535), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_543), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_556), .B(n_506), .Y(n_608) );
AOI21xp5_ASAP7_75t_SL g609 ( .A1(n_534), .A2(n_530), .B(n_533), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_554), .A2(n_541), .B(n_546), .Y(n_610) );
AOI21xp5_ASAP7_75t_L g611 ( .A1(n_574), .A2(n_508), .B(n_504), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_535), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_552), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_565), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_576), .A2(n_488), .B(n_503), .C(n_532), .Y(n_615) );
AOI322xp5_ASAP7_75t_L g616 ( .A1(n_567), .A2(n_509), .A3(n_504), .B1(n_519), .B2(n_454), .C1(n_521), .C2(n_253), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_559), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_546), .B(n_250), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_562), .A2(n_229), .B(n_230), .C(n_239), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_565), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_562), .B(n_230), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_579), .B(n_239), .Y(n_622) );
INVxp67_ASAP7_75t_L g623 ( .A(n_582), .Y(n_623) );
NAND2xp33_ASAP7_75t_L g624 ( .A(n_566), .B(n_249), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_578), .B(n_249), .C(n_253), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_580), .B(n_210), .Y(n_626) );
XNOR2x1_ASAP7_75t_L g627 ( .A(n_568), .B(n_210), .Y(n_627) );
INVx3_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
NAND2xp5_ASAP7_75t_SL g629 ( .A(n_581), .B(n_210), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_575), .B(n_210), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_582), .A2(n_571), .B1(n_577), .B2(n_572), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_564), .Y(n_632) );
XNOR2xp5_ASAP7_75t_L g633 ( .A(n_569), .B(n_570), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_569), .B(n_573), .Y(n_634) );
XNOR2xp5_ASAP7_75t_L g635 ( .A(n_558), .B(n_563), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_581), .A2(n_536), .B(n_539), .C(n_424), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_610), .B(n_583), .Y(n_637) );
AOI221xp5_ASAP7_75t_L g638 ( .A1(n_636), .A2(n_603), .B1(n_623), .B2(n_613), .C(n_599), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_594), .A2(n_585), .B1(n_600), .B2(n_602), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_588), .B(n_586), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_591), .Y(n_641) );
OAI21xp5_ASAP7_75t_SL g642 ( .A1(n_594), .A2(n_615), .B(n_611), .Y(n_642) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_593), .A2(n_592), .B1(n_601), .B2(n_597), .C(n_587), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_598), .A2(n_597), .B(n_604), .C(n_625), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_589), .A2(n_618), .B(n_626), .Y(n_645) );
O2A1O1Ixp33_ASAP7_75t_L g646 ( .A1(n_604), .A2(n_629), .B(n_621), .C(n_607), .Y(n_646) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_609), .A2(n_631), .B(n_616), .C(n_617), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_632), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_634), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_649), .B(n_633), .Y(n_650) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_642), .A2(n_624), .B(n_628), .C(n_617), .Y(n_651) );
OAI31xp33_ASAP7_75t_L g652 ( .A1(n_647), .A2(n_627), .A3(n_628), .B(n_635), .Y(n_652) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_638), .A2(n_609), .B(n_608), .C(n_590), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_637), .B(n_620), .Y(n_654) );
INVx2_ASAP7_75t_L g655 ( .A(n_641), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_648), .B(n_614), .Y(n_656) );
NOR3xp33_ASAP7_75t_L g657 ( .A(n_644), .B(n_619), .C(n_622), .Y(n_657) );
NOR2xp67_ASAP7_75t_L g658 ( .A(n_653), .B(n_639), .Y(n_658) );
OR3x1_ASAP7_75t_L g659 ( .A(n_652), .B(n_645), .C(n_646), .Y(n_659) );
AOI211xp5_ASAP7_75t_L g660 ( .A1(n_651), .A2(n_643), .B(n_640), .C(n_596), .Y(n_660) );
OAI222xp33_ASAP7_75t_L g661 ( .A1(n_654), .A2(n_634), .B1(n_584), .B2(n_596), .C1(n_595), .C2(n_605), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_658), .A2(n_657), .B1(n_654), .B2(n_650), .Y(n_662) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_659), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_660), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_663), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
OAI222xp33_ASAP7_75t_L g668 ( .A1(n_666), .A2(n_664), .B1(n_662), .B2(n_655), .C1(n_656), .C2(n_661), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_667), .A2(n_630), .B1(n_606), .B2(n_612), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_669), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_667), .B1(n_668), .B2(n_584), .Y(n_671) );
endmodule