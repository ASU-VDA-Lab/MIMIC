module fake_jpeg_6261_n_333 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_5),
.B(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_20),
.B(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_35),
.A2(n_29),
.B(n_28),
.C(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_44),
.Y(n_51)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_41),
.B1(n_27),
.B2(n_19),
.Y(n_63)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_54),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_39),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_18),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_23),
.B1(n_32),
.B2(n_17),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_35),
.Y(n_55)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_58),
.Y(n_88)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_34),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_28),
.B1(n_19),
.B2(n_30),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_34),
.B1(n_23),
.B2(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_35),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_70),
.B(n_73),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_81),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_37),
.B1(n_44),
.B2(n_41),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_44),
.B1(n_36),
.B2(n_37),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_63),
.Y(n_118)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_80),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_51),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_91),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_90),
.B1(n_95),
.B2(n_98),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_55),
.A2(n_37),
.B1(n_42),
.B2(n_36),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_62),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_36),
.Y(n_93)
);

NAND3xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_94),
.C(n_25),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_32),
.Y(n_94)
);

AO22x1_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_41),
.B1(n_40),
.B2(n_42),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_21),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_45),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_71),
.C(n_68),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_102),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_76),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_53),
.B(n_41),
.C(n_40),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_122),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_107),
.Y(n_131)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_113),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_53),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_114),
.Y(n_129)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_66),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_119),
.Y(n_143)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_95),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_125),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_40),
.B(n_16),
.C(n_27),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_88),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_97),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_127),
.A2(n_86),
.B1(n_25),
.B2(n_24),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_140),
.Y(n_162)
);

AOI32xp33_ASAP7_75t_L g133 ( 
.A1(n_103),
.A2(n_86),
.A3(n_93),
.B1(n_73),
.B2(n_83),
.Y(n_133)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_16),
.B(n_21),
.C(n_46),
.D(n_62),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_135),
.Y(n_160)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_93),
.B1(n_73),
.B2(n_64),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_150),
.B1(n_78),
.B2(n_77),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_89),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_141),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_56),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_149),
.Y(n_164)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_64),
.B1(n_60),
.B2(n_45),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_156),
.B1(n_100),
.B2(n_120),
.Y(n_180)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_59),
.B1(n_92),
.B2(n_91),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_110),
.Y(n_151)
);

INVx13_ASAP7_75t_L g170 ( 
.A(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_123),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_153),
.B(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_67),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_101),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_155),
.A2(n_102),
.B(n_115),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_97),
.B1(n_82),
.B2(n_57),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_99),
.C(n_108),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_159),
.B(n_172),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_108),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_181),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_168),
.Y(n_198)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_144),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_169),
.Y(n_195)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_124),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_72),
.Y(n_173)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_130),
.B(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_129),
.Y(n_178)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_128),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_179),
.B(n_192),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_193),
.B1(n_190),
.B2(n_188),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_104),
.B(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_100),
.C(n_145),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_187),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_126),
.B1(n_111),
.B2(n_122),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_17),
.B1(n_25),
.B2(n_24),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_186),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_155),
.A2(n_48),
.B(n_67),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_150),
.Y(n_188)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_189),
.B(n_183),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_191),
.A2(n_148),
.B1(n_158),
.B2(n_132),
.Y(n_197)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_197),
.A2(n_170),
.B1(n_22),
.B2(n_72),
.Y(n_247)
);

XOR2x2_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_133),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_204),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_191),
.A2(n_137),
.B1(n_146),
.B2(n_139),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_203),
.A2(n_193),
.B1(n_166),
.B2(n_168),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_152),
.Y(n_204)
);

AOI221xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_147),
.B1(n_151),
.B2(n_149),
.C(n_132),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_213),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_153),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_208),
.A2(n_211),
.B(n_167),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g211 ( 
.A1(n_162),
.A2(n_0),
.B(n_1),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_172),
.B(n_46),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_180),
.A2(n_24),
.B1(n_22),
.B2(n_17),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_189),
.B(n_170),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_217),
.B(n_182),
.C(n_171),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_230),
.C(n_235),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_192),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_174),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_239),
.B1(n_244),
.B2(n_245),
.Y(n_259)
);

AOI22x1_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_199),
.B1(n_197),
.B2(n_187),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_228),
.A2(n_229),
.B1(n_201),
.B2(n_22),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_185),
.B1(n_186),
.B2(n_169),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_178),
.C(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_162),
.Y(n_231)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_231),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_184),
.Y(n_232)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_232),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_198),
.A2(n_163),
.B(n_160),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_161),
.C(n_164),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_202),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_236),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_237),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_238),
.B(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_203),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_241),
.B(n_247),
.CI(n_215),
.CON(n_248),
.SN(n_248)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_242),
.Y(n_250)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_218),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_209),
.B(n_210),
.Y(n_245)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_211),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_265),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_194),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_253),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_194),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_256),
.C(n_262),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_219),
.C(n_221),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_226),
.C(n_228),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_204),
.C(n_212),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.C(n_268),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_195),
.C(n_201),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_241),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_240),
.B(n_46),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_261),
.B(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_227),
.B1(n_231),
.B2(n_232),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_284),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_243),
.B1(n_240),
.B2(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_273),
.A2(n_282),
.B1(n_283),
.B2(n_257),
.Y(n_291)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_274),
.B(n_275),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_234),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_276),
.Y(n_286)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_263),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_277),
.B(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_46),
.B1(n_1),
.B2(n_2),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_0),
.B(n_1),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_8),
.B(n_15),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_267),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_285),
.B(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

OAI221xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_267),
.B1(n_248),
.B2(n_266),
.C(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_255),
.C(n_254),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_295),
.C(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_252),
.C(n_256),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_271),
.B(n_253),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_272),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_21),
.C(n_2),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_0),
.C(n_3),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_3),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_273),
.B1(n_278),
.B2(n_281),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_300),
.A2(n_303),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_283),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_308),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_282),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_311),
.C(n_298),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_8),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_290),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_289),
.A2(n_3),
.B(n_4),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_9),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_288),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_299),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_313),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_316),
.B(n_318),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_294),
.C(n_10),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_7),
.A3(n_12),
.B1(n_11),
.B2(n_13),
.C1(n_6),
.C2(n_5),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_11),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_304),
.A2(n_3),
.B(n_4),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_11),
.Y(n_326)
);

AOI31xp33_ASAP7_75t_L g323 ( 
.A1(n_315),
.A2(n_300),
.A3(n_309),
.B(n_310),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_324),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_317),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_327),
.A2(n_328),
.B(n_325),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_321),
.A2(n_313),
.B(n_306),
.Y(n_328)
);

OAI221xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_329),
.B1(n_322),
.B2(n_319),
.C(n_13),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_5),
.B1(n_6),
.B2(n_324),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_5),
.Y(n_333)
);


endmodule