module fake_jpeg_20859_n_331 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_19),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.C(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_71),
.C(n_19),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_35),
.C(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_53),
.B(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_45),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_33),
.B1(n_34),
.B2(n_22),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_62),
.B1(n_21),
.B2(n_30),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_34),
.B1(n_33),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_58),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_35),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_91),
.Y(n_117)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_75),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_18),
.B1(n_26),
.B2(n_31),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_19),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_78),
.B(n_102),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_79),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_89),
.B1(n_107),
.B2(n_106),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_52),
.B(n_47),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_83),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_51),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_84),
.Y(n_136)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_46),
.B1(n_39),
.B2(n_41),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

INVx4_ASAP7_75t_SL g91 ( 
.A(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_94),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_25),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_26),
.B1(n_32),
.B2(n_28),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_100),
.B(n_101),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_55),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_103),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g104 ( 
.A(n_57),
.B(n_41),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_69),
.Y(n_125)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_111),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_47),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_58),
.A2(n_46),
.B1(n_39),
.B2(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_110),
.A2(n_114),
.B1(n_69),
.B2(n_70),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_11),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_68),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_118),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_68),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_122),
.A2(n_145),
.B1(n_103),
.B2(n_88),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_125),
.B(n_16),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_63),
.B1(n_30),
.B2(n_20),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_128),
.A2(n_131),
.B1(n_84),
.B2(n_87),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_45),
.B1(n_27),
.B2(n_17),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_82),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_134),
.B(n_136),
.Y(n_165)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_113),
.Y(n_137)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_27),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_141),
.Y(n_151)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_89),
.Y(n_146)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_27),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_149),
.Y(n_164)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_150),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_152),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_85),
.Y(n_153)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_104),
.C(n_100),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_154),
.B(n_168),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_107),
.B1(n_80),
.B2(n_91),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_155),
.A2(n_166),
.B1(n_144),
.B2(n_136),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_142),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_157),
.B(n_158),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_109),
.C(n_108),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_162),
.C(n_175),
.Y(n_187)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_161),
.A2(n_176),
.B(n_178),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_88),
.C(n_77),
.Y(n_162)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_98),
.B1(n_96),
.B2(n_77),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_116),
.B(n_111),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_169),
.A2(n_172),
.B1(n_176),
.B2(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_93),
.Y(n_170)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_25),
.B(n_29),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_181),
.B(n_120),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_125),
.A2(n_146),
.B1(n_121),
.B2(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_119),
.B(n_86),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_174),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_118),
.B(n_27),
.C(n_17),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_123),
.B(n_17),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_115),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_0),
.Y(n_213)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_0),
.B(n_1),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_122),
.B(n_16),
.C(n_29),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_182),
.B(n_140),
.C(n_117),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_185),
.A2(n_190),
.B1(n_178),
.B2(n_161),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_197),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_159),
.B(n_147),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_188),
.B(n_2),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_193),
.B1(n_196),
.B2(n_210),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_191),
.B(n_195),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_156),
.A2(n_140),
.B1(n_134),
.B2(n_133),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_133),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_163),
.A2(n_141),
.B1(n_137),
.B2(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_176),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_165),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_215),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_171),
.A2(n_132),
.B1(n_135),
.B2(n_127),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_206),
.B(n_213),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_202),
.A2(n_155),
.B1(n_177),
.B2(n_160),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_166),
.Y(n_204)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_204),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_181),
.A2(n_25),
.B(n_29),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_135),
.C(n_139),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_212),
.C(n_164),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_163),
.A2(n_136),
.B1(n_132),
.B2(n_139),
.Y(n_210)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_173),
.A2(n_16),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_214),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_13),
.C(n_12),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_158),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_202),
.A2(n_183),
.B(n_169),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_218),
.A2(n_216),
.B(n_231),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g220 ( 
.A1(n_185),
.A2(n_154),
.B(n_179),
.C(n_153),
.D(n_182),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_231),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_175),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_216),
.B(n_208),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_224),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_184),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_157),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_227),
.B(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_194),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_188),
.C(n_201),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_235),
.C(n_190),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_234),
.B1(n_213),
.B2(n_205),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_214),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_177),
.B1(n_3),
.B2(n_6),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_12),
.C(n_11),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_195),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_10),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_196),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_240),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_2),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_241),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_10),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_236),
.A2(n_192),
.B(n_208),
.C(n_211),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_251),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_223),
.C(n_239),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_199),
.B1(n_197),
.B2(n_189),
.Y(n_245)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_261),
.B1(n_234),
.B2(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_218),
.A2(n_206),
.B1(n_193),
.B2(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_219),
.B1(n_233),
.B2(n_237),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_213),
.B1(n_201),
.B2(n_212),
.Y(n_251)
);

XOR2x1_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_205),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_252),
.B(n_238),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_235),
.Y(n_265)
);

AOI22x1_ASAP7_75t_L g259 ( 
.A1(n_232),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_261),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_11),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_253),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_264),
.B(n_269),
.C(n_270),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_246),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_222),
.C(n_221),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_222),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_267),
.B1(n_274),
.B2(n_243),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_252),
.A2(n_217),
.B1(n_226),
.B2(n_221),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_229),
.B(n_228),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_275),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_217),
.C(n_241),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_260),
.C(n_251),
.Y(n_277)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_279),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_254),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_280),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_282),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_271),
.A2(n_258),
.B(n_263),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_268),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_280),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_279),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_275),
.Y(n_293)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_293),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_278),
.A2(n_245),
.B(n_248),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_294),
.B(n_281),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_286),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_269),
.C(n_264),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_301),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_300),
.B(n_291),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_270),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_304),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_295),
.C(n_277),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_265),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_283),
.B(n_263),
.C(n_276),
.Y(n_306)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_308),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_289),
.C(n_285),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_311),
.A2(n_313),
.B(n_314),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_312),
.A2(n_310),
.B1(n_314),
.B2(n_309),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_298),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_306),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_307),
.A2(n_287),
.B1(n_303),
.B2(n_294),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_316),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_308),
.A2(n_287),
.B1(n_303),
.B2(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_312),
.A2(n_296),
.B1(n_250),
.B2(n_256),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_320),
.B(n_259),
.CI(n_262),
.CON(n_323),
.SN(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_318),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_324),
.A2(n_325),
.B(n_315),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_321),
.B(n_317),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_322),
.B(n_316),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_319),
.C(n_259),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_8),
.C(n_9),
.Y(n_329)
);

HAxp5_ASAP7_75t_SL g330 ( 
.A(n_329),
.B(n_8),
.CON(n_330),
.SN(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_330),
.Y(n_331)
);


endmodule