module real_aes_8888_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_503;
wire n_287;
wire n_357;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_183;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_L g292 ( .A1(n_0), .A2(n_217), .B(n_219), .C(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_1), .A2(n_243), .B(n_244), .Y(n_242) );
AOI22xp33_ASAP7_75t_L g124 ( .A1(n_2), .A2(n_77), .B1(n_125), .B2(n_132), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_3), .B(n_254), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_4), .A2(n_53), .B1(n_175), .B2(n_176), .Y(n_174) );
INVx1_ASAP7_75t_L g176 ( .A(n_4), .Y(n_176) );
INVx1_ASAP7_75t_L g193 ( .A(n_5), .Y(n_193) );
AND2x6_ASAP7_75t_L g217 ( .A(n_5), .B(n_191), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_5), .B(n_522), .Y(n_521) );
OAI22xp5_ASAP7_75t_SL g169 ( .A1(n_6), .A2(n_170), .B1(n_171), .B2(n_180), .Y(n_169) );
INVx1_ASAP7_75t_L g180 ( .A(n_6), .Y(n_180) );
INVx1_ASAP7_75t_L g318 ( .A(n_7), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_8), .B(n_227), .Y(n_295) );
AO22x2_ASAP7_75t_L g91 ( .A1(n_9), .A2(n_29), .B1(n_92), .B2(n_93), .Y(n_91) );
INVx1_ASAP7_75t_L g209 ( .A(n_10), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g81 ( .A1(n_11), .A2(n_50), .B1(n_82), .B2(n_83), .Y(n_81) );
INVx1_ASAP7_75t_L g83 ( .A(n_11), .Y(n_83) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_11), .A2(n_262), .B(n_303), .C(n_305), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_12), .B(n_254), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_13), .A2(n_74), .B1(n_148), .B2(n_151), .Y(n_147) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_14), .A2(n_31), .B1(n_92), .B2(n_96), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_15), .B(n_350), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g171 ( .A1(n_16), .A2(n_172), .B1(n_173), .B2(n_179), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_16), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g115 ( .A1(n_17), .A2(n_56), .B1(n_116), .B2(n_121), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_18), .A2(n_248), .B(n_279), .C(n_282), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_19), .B(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_20), .B(n_227), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g211 ( .A(n_21), .Y(n_211) );
INVx1_ASAP7_75t_L g260 ( .A(n_22), .Y(n_260) );
AOI22xp5_ASAP7_75t_SL g518 ( .A1(n_22), .A2(n_84), .B1(n_85), .B2(n_260), .Y(n_518) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_23), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_24), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_25), .A2(n_39), .B1(n_139), .B2(n_143), .Y(n_138) );
INVx1_ASAP7_75t_L g347 ( .A(n_26), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_27), .A2(n_63), .B1(n_155), .B2(n_159), .Y(n_154) );
INVx2_ASAP7_75t_L g215 ( .A(n_28), .Y(n_215) );
CKINVDCx20_ASAP7_75t_R g297 ( .A(n_30), .Y(n_297) );
OAI221xp5_ASAP7_75t_L g184 ( .A1(n_31), .A2(n_42), .B1(n_51), .B2(n_185), .C(n_186), .Y(n_184) );
INVxp67_ASAP7_75t_L g187 ( .A(n_31), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_32), .A2(n_248), .B(n_249), .C(n_251), .Y(n_247) );
INVxp67_ASAP7_75t_L g348 ( .A(n_33), .Y(n_348) );
CKINVDCx14_ASAP7_75t_R g245 ( .A(n_34), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_35), .A2(n_219), .B(n_259), .C(n_266), .Y(n_258) );
INVx1_ASAP7_75t_L g527 ( .A(n_35), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g315 ( .A1(n_36), .A2(n_229), .B(n_316), .C(n_317), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g268 ( .A(n_37), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_38), .Y(n_344) );
INVx1_ASAP7_75t_L g277 ( .A(n_40), .Y(n_277) );
XOR2xp5_ASAP7_75t_L g528 ( .A(n_41), .B(n_84), .Y(n_528) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_42), .A2(n_67), .B1(n_92), .B2(n_96), .Y(n_99) );
INVxp67_ASAP7_75t_L g188 ( .A(n_42), .Y(n_188) );
CKINVDCx14_ASAP7_75t_R g314 ( .A(n_43), .Y(n_314) );
INVx1_ASAP7_75t_L g191 ( .A(n_44), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_45), .Y(n_102) );
INVx1_ASAP7_75t_L g208 ( .A(n_46), .Y(n_208) );
INVx1_ASAP7_75t_SL g250 ( .A(n_47), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_48), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_49), .B(n_254), .Y(n_284) );
INVx1_ASAP7_75t_L g82 ( .A(n_50), .Y(n_82) );
AO22x2_ASAP7_75t_L g101 ( .A1(n_51), .A2(n_71), .B1(n_92), .B2(n_93), .Y(n_101) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_52), .A2(n_57), .B1(n_104), .B2(n_110), .Y(n_103) );
INVx1_ASAP7_75t_L g175 ( .A(n_53), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_54), .A2(n_243), .B(n_313), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_55), .A2(n_75), .B1(n_163), .B2(n_166), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_58), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_59), .A2(n_243), .B(n_300), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_60), .A2(n_342), .B(n_343), .Y(n_341) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_61), .Y(n_257) );
INVx1_ASAP7_75t_L g301 ( .A(n_62), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_64), .A2(n_174), .B1(n_177), .B2(n_178), .Y(n_173) );
INVx1_ASAP7_75t_L g177 ( .A(n_64), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_65), .A2(n_243), .B(n_276), .Y(n_275) );
INVx1_ASAP7_75t_L g304 ( .A(n_66), .Y(n_304) );
INVx2_ASAP7_75t_L g206 ( .A(n_68), .Y(n_206) );
INVx1_ASAP7_75t_L g294 ( .A(n_69), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_70), .A2(n_219), .B(n_222), .C(n_231), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_72), .B(n_204), .Y(n_319) );
INVx1_ASAP7_75t_L g92 ( .A(n_73), .Y(n_92) );
INVx1_ASAP7_75t_L g94 ( .A(n_73), .Y(n_94) );
INVx2_ASAP7_75t_L g280 ( .A(n_76), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_181), .B1(n_194), .B2(n_514), .C(n_517), .Y(n_78) );
XNOR2xp5_ASAP7_75t_L g79 ( .A(n_80), .B(n_169), .Y(n_79) );
AOI22xp5_ASAP7_75t_L g80 ( .A1(n_81), .A2(n_84), .B1(n_85), .B2(n_168), .Y(n_80) );
CKINVDCx14_ASAP7_75t_R g168 ( .A(n_81), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g222 ( .A1(n_82), .A2(n_223), .B(n_226), .C(n_228), .Y(n_222) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NAND2x1_ASAP7_75t_L g85 ( .A(n_86), .B(n_136), .Y(n_85) );
NOR2xp33_ASAP7_75t_L g86 ( .A(n_87), .B(n_114), .Y(n_86) );
OAI21xp5_ASAP7_75t_SL g87 ( .A1(n_88), .A2(n_102), .B(n_103), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x6_ASAP7_75t_L g89 ( .A(n_90), .B(n_97), .Y(n_89) );
AND2x4_ASAP7_75t_L g121 ( .A(n_90), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_95), .Y(n_90) );
AND2x2_ASAP7_75t_L g109 ( .A(n_91), .B(n_99), .Y(n_109) );
INVx2_ASAP7_75t_L g131 ( .A(n_91), .Y(n_131) );
INVx1_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_94), .Y(n_96) );
INVx2_ASAP7_75t_L g108 ( .A(n_95), .Y(n_108) );
INVx1_ASAP7_75t_L g120 ( .A(n_95), .Y(n_120) );
OR2x2_ASAP7_75t_L g130 ( .A(n_95), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g135 ( .A(n_95), .B(n_131), .Y(n_135) );
AND2x6_ASAP7_75t_L g150 ( .A(n_97), .B(n_129), .Y(n_150) );
AND2x4_ASAP7_75t_L g152 ( .A(n_97), .B(n_135), .Y(n_152) );
AND2x2_ASAP7_75t_L g158 ( .A(n_97), .B(n_142), .Y(n_158) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_100), .Y(n_97) );
AND2x2_ASAP7_75t_L g128 ( .A(n_98), .B(n_101), .Y(n_128) );
INVx2_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
AND2x2_ASAP7_75t_L g141 ( .A(n_99), .B(n_123), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_99), .B(n_101), .Y(n_146) );
INVx1_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g107 ( .A(n_101), .Y(n_107) );
INVx1_ASAP7_75t_L g123 ( .A(n_101), .Y(n_123) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x4_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
AND2x2_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g113 ( .A(n_107), .Y(n_113) );
AND2x2_ASAP7_75t_L g142 ( .A(n_108), .B(n_131), .Y(n_142) );
AND2x4_ASAP7_75t_L g112 ( .A(n_109), .B(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g118 ( .A(n_109), .B(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_124), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x6_ASAP7_75t_L g167 ( .A(n_120), .B(n_146), .Y(n_167) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx4_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
AND2x6_ASAP7_75t_L g134 ( .A(n_128), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g161 ( .A(n_128), .B(n_142), .Y(n_161) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_SL g132 ( .A(n_133), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g165 ( .A(n_135), .B(n_141), .Y(n_165) );
NOR2x1_ASAP7_75t_L g136 ( .A(n_137), .B(n_153), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_147), .Y(n_137) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
AND2x4_ASAP7_75t_L g144 ( .A(n_142), .B(n_145), .Y(n_144) );
BUFx2_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx11_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_162), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx8_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g170 ( .A(n_171), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_173), .Y(n_179) );
INVx1_ASAP7_75t_L g178 ( .A(n_174), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_183), .Y(n_182) );
AND3x1_ASAP7_75t_SL g183 ( .A(n_184), .B(n_189), .C(n_192), .Y(n_183) );
INVxp67_ASAP7_75t_L g522 ( .A(n_184), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
INVx1_ASAP7_75t_SL g523 ( .A(n_189), .Y(n_523) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_189), .A2(n_219), .B(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g532 ( .A(n_189), .Y(n_532) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_190), .B(n_193), .Y(n_526) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OR2x2_ASAP7_75t_SL g531 ( .A(n_192), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_196), .B(n_469), .Y(n_195) );
NOR4xp25_ASAP7_75t_L g196 ( .A(n_197), .B(n_406), .C(n_440), .D(n_456), .Y(n_196) );
NAND4xp25_ASAP7_75t_SL g197 ( .A(n_198), .B(n_332), .C(n_370), .D(n_386), .Y(n_197) );
AOI222xp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_269), .B1(n_307), .B2(n_320), .C1(n_325), .C2(n_331), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI31xp33_ASAP7_75t_L g502 ( .A1(n_200), .A2(n_503), .A3(n_504), .B(n_506), .Y(n_502) );
OR2x2_ASAP7_75t_L g200 ( .A(n_201), .B(n_237), .Y(n_200) );
AND2x2_ASAP7_75t_L g477 ( .A(n_201), .B(n_239), .Y(n_477) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_SL g324 ( .A(n_202), .Y(n_324) );
AND2x2_ASAP7_75t_L g331 ( .A(n_202), .B(n_255), .Y(n_331) );
AND2x2_ASAP7_75t_L g391 ( .A(n_202), .B(n_240), .Y(n_391) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_210), .B(n_233), .Y(n_202) );
INVx3_ASAP7_75t_L g254 ( .A(n_203), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_203), .B(n_268), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g296 ( .A(n_203), .B(n_297), .Y(n_296) );
INVx4_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
BUFx6f_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g340 ( .A(n_205), .Y(n_340) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
AND2x2_ASAP7_75t_SL g236 ( .A(n_206), .B(n_207), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_212), .A2(n_236), .B(n_257), .C(n_258), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g290 ( .A1(n_212), .A2(n_291), .B(n_292), .Y(n_290) );
NAND2x1p5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
AND2x4_ASAP7_75t_L g243 ( .A(n_213), .B(n_217), .Y(n_243) );
AND2x2_ASAP7_75t_L g213 ( .A(n_214), .B(n_216), .Y(n_213) );
INVx1_ASAP7_75t_L g265 ( .A(n_214), .Y(n_265) );
INVx1_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g220 ( .A(n_215), .Y(n_220) );
INVx1_ASAP7_75t_L g283 ( .A(n_215), .Y(n_283) );
INVx1_ASAP7_75t_L g221 ( .A(n_216), .Y(n_221) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_216), .Y(n_225) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_216), .Y(n_227) );
INVx3_ASAP7_75t_L g262 ( .A(n_216), .Y(n_262) );
INVx4_ASAP7_75t_SL g232 ( .A(n_217), .Y(n_232) );
BUFx3_ASAP7_75t_L g266 ( .A(n_217), .Y(n_266) );
INVx5_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
AND2x2_ASAP7_75t_L g516 ( .A(n_219), .B(n_266), .Y(n_516) );
AND2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
BUFx3_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_220), .Y(n_252) );
O2A1O1Ixp5_ASAP7_75t_L g293 ( .A1(n_223), .A2(n_228), .B(n_294), .C(n_295), .Y(n_293) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx4_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
INVx4_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
INVx2_ASAP7_75t_L g316 ( .A(n_227), .Y(n_316) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g305 ( .A(n_230), .Y(n_305) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_232), .A2(n_245), .B(n_246), .C(n_247), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g276 ( .A1(n_232), .A2(n_246), .B(n_277), .C(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_SL g300 ( .A1(n_232), .A2(n_246), .B(n_301), .C(n_302), .Y(n_300) );
O2A1O1Ixp33_ASAP7_75t_SL g313 ( .A1(n_232), .A2(n_246), .B(n_314), .C(n_315), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_SL g343 ( .A1(n_232), .A2(n_246), .B(n_344), .C(n_345), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g350 ( .A(n_235), .Y(n_350) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g289 ( .A(n_236), .Y(n_289) );
OA21x2_ASAP7_75t_L g311 ( .A1(n_236), .A2(n_312), .B(n_319), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_237), .B(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_238), .B(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_238), .B(n_335), .Y(n_381) );
AND2x2_ASAP7_75t_L g474 ( .A(n_238), .B(n_414), .Y(n_474) );
OAI321xp33_ASAP7_75t_L g508 ( .A1(n_238), .A2(n_324), .A3(n_481), .B1(n_509), .B2(n_511), .C(n_512), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g512 ( .A(n_238), .B(n_310), .C(n_421), .D(n_513), .Y(n_512) );
AND2x4_ASAP7_75t_L g238 ( .A(n_239), .B(n_255), .Y(n_238) );
AND2x2_ASAP7_75t_L g376 ( .A(n_239), .B(n_322), .Y(n_376) );
AND2x2_ASAP7_75t_L g395 ( .A(n_239), .B(n_324), .Y(n_395) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g323 ( .A(n_240), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g351 ( .A(n_240), .B(n_255), .Y(n_351) );
AND2x2_ASAP7_75t_L g437 ( .A(n_240), .B(n_322), .Y(n_437) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_242), .B(n_253), .Y(n_240) );
OA21x2_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_275), .B(n_284), .Y(n_274) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_241), .A2(n_299), .B(n_306), .Y(n_298) );
BUFx2_ASAP7_75t_L g342 ( .A(n_243), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_248), .B(n_250), .Y(n_249) );
INVx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx3_ASAP7_75t_SL g322 ( .A(n_255), .Y(n_322) );
AND2x2_ASAP7_75t_L g369 ( .A(n_255), .B(n_356), .Y(n_369) );
OR2x2_ASAP7_75t_L g402 ( .A(n_255), .B(n_324), .Y(n_402) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_255), .Y(n_409) );
AND2x2_ASAP7_75t_L g438 ( .A(n_255), .B(n_323), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_255), .B(n_411), .Y(n_453) );
AND2x2_ASAP7_75t_L g485 ( .A(n_255), .B(n_477), .Y(n_485) );
AND2x2_ASAP7_75t_L g494 ( .A(n_255), .B(n_336), .Y(n_494) );
OR2x6_ASAP7_75t_L g255 ( .A(n_256), .B(n_267), .Y(n_255) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_261), .B(n_263), .C(n_264), .Y(n_259) );
OAI22xp33_ASAP7_75t_L g346 ( .A1(n_261), .A2(n_281), .B1(n_347), .B2(n_348), .Y(n_346) );
INVx5_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_262), .B(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g345 ( .A(n_265), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_285), .Y(n_270) );
INVx1_ASAP7_75t_SL g462 ( .A(n_271), .Y(n_462) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g327 ( .A(n_272), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g309 ( .A(n_273), .B(n_287), .Y(n_309) );
AND2x2_ASAP7_75t_L g398 ( .A(n_273), .B(n_311), .Y(n_398) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g368 ( .A(n_274), .B(n_298), .Y(n_368) );
OR2x2_ASAP7_75t_L g379 ( .A(n_274), .B(n_311), .Y(n_379) );
AND2x2_ASAP7_75t_L g405 ( .A(n_274), .B(n_311), .Y(n_405) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_274), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_281), .B(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_285), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_285), .B(n_462), .Y(n_461) );
INVx2_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g378 ( .A(n_286), .B(n_379), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g464 ( .A1(n_286), .A2(n_368), .A3(n_374), .B1(n_405), .B2(n_455), .C1(n_465), .C2(n_467), .Y(n_464) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_298), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_287), .B(n_310), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_287), .B(n_311), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_287), .B(n_328), .Y(n_385) );
AND2x2_ASAP7_75t_L g439 ( .A(n_287), .B(n_405), .Y(n_439) );
INVx1_ASAP7_75t_L g443 ( .A(n_287), .Y(n_443) );
AND2x2_ASAP7_75t_L g455 ( .A(n_287), .B(n_298), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_287), .B(n_327), .Y(n_487) );
INVx4_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g352 ( .A(n_288), .B(n_298), .Y(n_352) );
BUFx3_ASAP7_75t_L g366 ( .A(n_288), .Y(n_366) );
AND3x2_ASAP7_75t_L g448 ( .A(n_288), .B(n_428), .C(n_449), .Y(n_448) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_290), .B(n_296), .Y(n_288) );
NAND3xp33_ASAP7_75t_L g308 ( .A(n_298), .B(n_309), .C(n_310), .Y(n_308) );
INVx1_ASAP7_75t_SL g328 ( .A(n_298), .Y(n_328) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_298), .Y(n_433) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g427 ( .A(n_309), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g434 ( .A(n_309), .Y(n_434) );
AND2x2_ASAP7_75t_L g472 ( .A(n_310), .B(n_450), .Y(n_472) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx3_ASAP7_75t_L g353 ( .A(n_311), .Y(n_353) );
AND2x2_ASAP7_75t_L g428 ( .A(n_311), .B(n_328), .Y(n_428) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
OR2x2_ASAP7_75t_L g372 ( .A(n_322), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g491 ( .A(n_322), .B(n_391), .Y(n_491) );
AND2x2_ASAP7_75t_L g505 ( .A(n_322), .B(n_324), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_323), .B(n_336), .Y(n_446) );
AND2x2_ASAP7_75t_L g493 ( .A(n_323), .B(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g356 ( .A(n_324), .B(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g373 ( .A(n_324), .B(n_336), .Y(n_373) );
INVx1_ASAP7_75t_L g383 ( .A(n_324), .Y(n_383) );
AND2x2_ASAP7_75t_L g414 ( .A(n_324), .B(n_336), .Y(n_414) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g456 ( .A1(n_326), .A2(n_457), .B1(n_461), .B2(n_463), .C(n_464), .Y(n_456) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_327), .B(n_329), .Y(n_326) );
AND2x2_ASAP7_75t_L g360 ( .A(n_327), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_330), .B(n_367), .Y(n_510) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_352), .A3(n_353), .B1(n_354), .B2(n_360), .C1(n_362), .C2(n_369), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_351), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_335), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_335), .B(n_401), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g424 ( .A1(n_335), .A2(n_351), .B(n_425), .C(n_426), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_335), .B(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_335), .B(n_395), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_335), .B(n_477), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_335), .B(n_505), .Y(n_504) );
BUFx3_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_336), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_336), .B(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g466 ( .A(n_336), .B(n_353), .Y(n_466) );
OA21x2_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_341), .B(n_349), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_338), .A2(n_358), .B(n_359), .Y(n_357) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g358 ( .A(n_341), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_349), .Y(n_359) );
INVx1_ASAP7_75t_L g441 ( .A(n_351), .Y(n_441) );
OAI31xp33_ASAP7_75t_L g451 ( .A1(n_351), .A2(n_376), .A3(n_452), .B(n_454), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_351), .B(n_357), .Y(n_503) );
INVx1_ASAP7_75t_SL g364 ( .A(n_352), .Y(n_364) );
AND2x2_ASAP7_75t_L g397 ( .A(n_352), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g478 ( .A(n_352), .B(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g363 ( .A(n_353), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g388 ( .A(n_353), .Y(n_388) );
AND2x2_ASAP7_75t_L g415 ( .A(n_353), .B(n_368), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_353), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g507 ( .A(n_353), .B(n_455), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_355), .B(n_425), .Y(n_498) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g394 ( .A(n_357), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g412 ( .A(n_357), .Y(n_412) );
NAND2xp33_ASAP7_75t_SL g362 ( .A(n_363), .B(n_365), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g406 ( .A1(n_364), .A2(n_407), .B(n_413), .C(n_429), .Y(n_406) );
OR2x2_ASAP7_75t_L g481 ( .A(n_364), .B(n_462), .Y(n_481) );
OR2x2_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
CKINVDCx16_ASAP7_75t_R g418 ( .A(n_366), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_366), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g387 ( .A(n_368), .B(n_388), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_374), .B(n_377), .C(n_380), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g421 ( .A(n_373), .Y(n_421) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_376), .B(n_414), .Y(n_419) );
INVx1_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OR2x2_ASAP7_75t_L g384 ( .A(n_379), .B(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g417 ( .A(n_379), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g479 ( .A(n_379), .Y(n_479) );
AOI21xp33_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_382), .B(n_384), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_382), .A2(n_393), .B(n_396), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_389), .B(n_392), .C(n_399), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_387), .B(n_443), .Y(n_442) );
INVx1_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_390), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g403 ( .A(n_391), .Y(n_403) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_393), .A2(n_459), .B(n_460), .Y(n_458) );
INVx1_ASAP7_75t_SL g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_398), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g423 ( .A(n_398), .Y(n_423) );
AOI21xp33_ASAP7_75t_SL g399 ( .A1(n_400), .A2(n_403), .B(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g454 ( .A(n_405), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_411), .B(n_437), .Y(n_463) );
AND2x2_ASAP7_75t_L g476 ( .A(n_411), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g490 ( .A(n_411), .B(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g500 ( .A(n_411), .B(n_438), .Y(n_500) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_416), .C(n_424), .Y(n_413) );
INVx1_ASAP7_75t_L g460 ( .A(n_414), .Y(n_460) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_420), .B2(n_422), .Y(n_416) );
OR2x2_ASAP7_75t_L g422 ( .A(n_418), .B(n_423), .Y(n_422) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_418), .B(n_479), .Y(n_501) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g495 ( .A(n_428), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_435), .B1(n_438), .B2(n_439), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
INVx1_ASAP7_75t_L g513 ( .A(n_433), .Y(n_513) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g459 ( .A(n_437), .Y(n_459) );
OAI211xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_442), .B(n_444), .C(n_451), .Y(n_440) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVxp67_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_459), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR5xp2_ASAP7_75t_L g469 ( .A(n_470), .B(n_488), .C(n_496), .D(n_502), .E(n_508), .Y(n_469) );
OAI211xp5_ASAP7_75t_SL g470 ( .A1(n_471), .A2(n_473), .B(n_475), .C(n_482), .Y(n_470) );
INVxp67_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B(n_480), .Y(n_475) );
OAI21xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_485), .B(n_486), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_485), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AOI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_495), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_SL g511 ( .A(n_491), .Y(n_511) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_499), .B(n_501), .Y(n_496) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_515), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_516), .Y(n_515) );
OAI322xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .A3(n_523), .B1(n_524), .B2(n_527), .C1(n_528), .C2(n_529), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_531), .Y(n_530) );
endmodule