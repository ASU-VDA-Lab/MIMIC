module fake_ariane_1578_n_3690 (n_295, n_356, n_556, n_170, n_190, n_698, n_695, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_691, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_694, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_699, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_693, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_696, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_692, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_697, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_3690);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_698;
input n_695;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_691;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_694;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_699;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_693;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_696;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_692;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_697;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_3690;

wire n_2752;
wire n_3527;
wire n_913;
wire n_1681;
wire n_2163;
wire n_3432;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_3619;
wire n_2484;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_3152;
wire n_2346;
wire n_3434;
wire n_1469;
wire n_1353;
wire n_3056;
wire n_3500;
wire n_3480;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_3268;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_3181;
wire n_850;
wire n_2993;
wire n_1916;
wire n_2879;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_2818;
wire n_3578;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_3487;
wire n_1238;
wire n_2694;
wire n_3668;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_3352;
wire n_3517;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_3561;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_3526;
wire n_2042;
wire n_2123;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_3154;
wire n_2646;
wire n_1298;
wire n_737;
wire n_2653;
wire n_2873;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_3115;
wire n_2278;
wire n_3330;
wire n_3514;
wire n_1088;
wire n_1424;
wire n_766;
wire n_2976;
wire n_1835;
wire n_3383;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_3416;
wire n_870;
wire n_2547;
wire n_3382;
wire n_1453;
wire n_958;
wire n_945;
wire n_2554;
wire n_3145;
wire n_2248;
wire n_3665;
wire n_3063;
wire n_813;
wire n_3281;
wire n_3535;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_2908;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_3220;
wire n_2960;
wire n_754;
wire n_903;
wire n_3270;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_3348;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_3261;
wire n_1761;
wire n_829;
wire n_1062;
wire n_738;
wire n_3679;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_2906;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_3283;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_3657;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_3451;
wire n_2322;
wire n_2746;
wire n_3419;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_1944;
wire n_2370;
wire n_2663;
wire n_2233;
wire n_2914;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_3545;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_2878;
wire n_1241;
wire n_821;
wire n_770;
wire n_3252;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_3315;
wire n_1145;
wire n_3523;
wire n_971;
wire n_3144;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_3606;
wire n_786;
wire n_1404;
wire n_3347;
wire n_3420;
wire n_868;
wire n_3474;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_3150;
wire n_2950;
wire n_1542;
wire n_3552;
wire n_1314;
wire n_3639;
wire n_3254;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_3121;
wire n_2847;
wire n_884;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_3209;
wire n_3324;
wire n_3015;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_2988;
wire n_1636;
wire n_3482;
wire n_823;
wire n_1900;
wire n_1074;
wire n_3230;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_3207;
wire n_3641;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_3073;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_3183;
wire n_3571;
wire n_1013;
wire n_1495;
wire n_3607;
wire n_1637;
wire n_3297;
wire n_2571;
wire n_2427;
wire n_3325;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2874;
wire n_3003;
wire n_3049;
wire n_3136;
wire n_2867;
wire n_3634;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_2899;
wire n_1548;
wire n_3066;
wire n_1811;
wire n_2045;
wire n_3274;
wire n_3013;
wire n_3612;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_2902;
wire n_1544;
wire n_3271;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_3164;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2956;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_3652;
wire n_3449;
wire n_2788;
wire n_1443;
wire n_1021;
wire n_3089;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_3084;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_3458;
wire n_2727;
wire n_942;
wire n_3580;
wire n_1437;
wire n_3511;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_2909;
wire n_1416;
wire n_3554;
wire n_1461;
wire n_2717;
wire n_3012;
wire n_1391;
wire n_2981;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_3472;
wire n_2527;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_3126;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_2038;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_3485;
wire n_1594;
wire n_1935;
wire n_2806;
wire n_3191;
wire n_1716;
wire n_1872;
wire n_3562;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3119;
wire n_1108;
wire n_3588;
wire n_851;
wire n_1590;
wire n_1351;
wire n_3280;
wire n_3234;
wire n_3413;
wire n_2216;
wire n_1274;
wire n_3539;
wire n_2426;
wire n_1819;
wire n_3095;
wire n_947;
wire n_2134;
wire n_1260;
wire n_930;
wire n_1179;
wire n_3284;
wire n_2703;
wire n_2926;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_3391;
wire n_3506;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_3678;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_2791;
wire n_2683;
wire n_3212;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_3529;
wire n_2970;
wire n_3159;
wire n_992;
wire n_966;
wire n_955;
wire n_3549;
wire n_3624;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_3192;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_3306;
wire n_3250;
wire n_3029;
wire n_2398;
wire n_3538;
wire n_1376;
wire n_1292;
wire n_1972;
wire n_2015;
wire n_1178;
wire n_2925;
wire n_1435;
wire n_3407;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_3460;
wire n_3544;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2952;
wire n_3530;
wire n_2415;
wire n_2693;
wire n_2877;
wire n_3120;
wire n_2922;
wire n_3000;
wire n_2871;
wire n_2930;
wire n_3193;
wire n_3240;
wire n_2745;
wire n_2087;
wire n_1491;
wire n_931;
wire n_2628;
wire n_3219;
wire n_3362;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_3510;
wire n_1389;
wire n_3393;
wire n_3172;
wire n_2155;
wire n_2659;
wire n_1139;
wire n_2836;
wire n_3688;
wire n_2439;
wire n_2864;
wire n_1312;
wire n_1717;
wire n_3604;
wire n_1812;
wire n_3651;
wire n_824;
wire n_2172;
wire n_2601;
wire n_3614;
wire n_892;
wire n_1880;
wire n_2365;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_3116;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_3176;
wire n_3629;
wire n_3666;
wire n_3372;
wire n_1623;
wire n_990;
wire n_3559;
wire n_1903;
wire n_867;
wire n_2147;
wire n_3479;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2888;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_2921;
wire n_3046;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_3021;
wire n_3257;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_3496;
wire n_3493;
wire n_2557;
wire n_2695;
wire n_2898;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_3567;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2954;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_2903;
wire n_974;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_3625;
wire n_2467;
wire n_3375;
wire n_2768;
wire n_1914;
wire n_965;
wire n_2253;
wire n_934;
wire n_2213;
wire n_3515;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_2924;
wire n_1209;
wire n_1563;
wire n_1020;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_3438;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_3187;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_3170;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_3147;
wire n_2287;
wire n_836;
wire n_2223;
wire n_3082;
wire n_1279;
wire n_3415;
wire n_3661;
wire n_2473;
wire n_3320;
wire n_2144;
wire n_2511;
wire n_3464;
wire n_3414;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_2919;
wire n_3210;
wire n_1483;
wire n_3108;
wire n_1363;
wire n_2681;
wire n_3397;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_3467;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_3031;
wire n_2262;
wire n_3179;
wire n_2565;
wire n_1237;
wire n_3262;
wire n_927;
wire n_1095;
wire n_2980;
wire n_1728;
wire n_2335;
wire n_3078;
wire n_706;
wire n_2120;
wire n_3239;
wire n_2631;
wire n_3215;
wire n_3311;
wire n_3516;
wire n_1401;
wire n_1419;
wire n_3138;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_3528;
wire n_1651;
wire n_3087;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_2677;
wire n_1826;
wire n_3171;
wire n_3577;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_3185;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_2996;
wire n_1592;
wire n_2812;
wire n_3660;
wire n_2662;
wire n_1259;
wire n_3300;
wire n_2801;
wire n_1177;
wire n_3104;
wire n_3074;
wire n_2655;
wire n_1231;
wire n_3246;
wire n_2132;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3589;
wire n_3623;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_3615;
wire n_3267;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_3054;
wire n_2811;
wire n_3019;
wire n_1795;
wire n_3200;
wire n_1384;
wire n_3642;
wire n_2237;
wire n_2146;
wire n_2983;
wire n_1868;
wire n_3276;
wire n_3601;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_3498;
wire n_3513;
wire n_3682;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_3377;
wire n_1518;
wire n_3323;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_3675;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_3466;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_3572;
wire n_2975;
wire n_3332;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_3374;
wire n_3471;
wire n_1484;
wire n_1901;
wire n_2055;
wire n_2998;
wire n_3465;
wire n_2027;
wire n_2932;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_3118;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_3039;
wire n_2195;
wire n_2194;
wire n_2937;
wire n_3508;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_3057;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1105;
wire n_3599;
wire n_3618;
wire n_3022;
wire n_703;
wire n_1349;
wire n_1709;
wire n_3318;
wire n_1061;
wire n_3385;
wire n_2102;
wire n_3477;
wire n_3286;
wire n_3370;
wire n_874;
wire n_2286;
wire n_3494;
wire n_2023;
wire n_1278;
wire n_707;
wire n_3443;
wire n_3401;
wire n_983;
wire n_3036;
wire n_2783;
wire n_2599;
wire n_727;
wire n_2075;
wire n_1726;
wire n_3263;
wire n_3569;
wire n_2523;
wire n_1945;
wire n_3542;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_1162;
wire n_2031;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_2118;
wire n_1740;
wire n_3222;
wire n_1602;
wire n_3139;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_3025;
wire n_3636;
wire n_3051;
wire n_3205;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_3653;
wire n_3035;
wire n_729;
wire n_887;
wire n_3403;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_1205;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2944;
wire n_2861;
wire n_2780;
wire n_3023;
wire n_1120;
wire n_3439;
wire n_1202;
wire n_2254;
wire n_3130;
wire n_3290;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_3602;
wire n_1402;
wire n_957;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_3418;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_3611;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_3338;
wire n_2962;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_3156;
wire n_2256;
wire n_1189;
wire n_3337;
wire n_1089;
wire n_3424;
wire n_3326;
wire n_3356;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_1502;
wire n_3044;
wire n_1523;
wire n_2190;
wire n_3501;
wire n_3492;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_3216;
wire n_3224;
wire n_3568;
wire n_1969;
wire n_2708;
wire n_735;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_2379;
wire n_3579;
wire n_3245;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_845;
wire n_888;
wire n_2894;
wire n_2300;
wire n_2949;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_3214;
wire n_3551;
wire n_1708;
wire n_3085;
wire n_3373;
wire n_1222;
wire n_2284;
wire n_3005;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_3364;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_1919;
wire n_710;
wire n_2994;
wire n_1791;
wire n_2508;
wire n_3186;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_3417;
wire n_2449;
wire n_890;
wire n_842;
wire n_3626;
wire n_1898;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_3180;
wire n_3648;
wire n_3423;
wire n_1975;
wire n_1373;
wire n_742;
wire n_1081;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_3671;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_3392;
wire n_1800;
wire n_982;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_2904;
wire n_3064;
wire n_3199;
wire n_1529;
wire n_3353;
wire n_1227;
wire n_3531;
wire n_2127;
wire n_2946;
wire n_3166;
wire n_3151;
wire n_3649;
wire n_3684;
wire n_3333;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_3065;
wire n_3016;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_3135;
wire n_3367;
wire n_3669;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_3024;
wire n_2772;
wire n_3564;
wire n_862;
wire n_1700;
wire n_2637;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_2893;
wire n_2959;
wire n_1532;
wire n_3277;
wire n_1171;
wire n_1030;
wire n_785;
wire n_3161;
wire n_3208;
wire n_2389;
wire n_1309;
wire n_3582;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2916;
wire n_2576;
wire n_3459;
wire n_3617;
wire n_704;
wire n_2958;
wire n_3365;
wire n_1060;
wire n_1714;
wire n_1044;
wire n_2696;
wire n_3340;
wire n_2140;
wire n_1748;
wire n_1301;
wire n_873;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_3400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_3486;
wire n_1527;
wire n_1513;
wire n_2581;
wire n_1783;
wire n_3656;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_3069;
wire n_2992;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_3197;
wire n_1993;
wire n_1545;
wire n_3586;
wire n_2629;
wire n_3369;
wire n_3256;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_3670;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_3302;
wire n_1605;
wire n_1078;
wire n_3060;
wire n_2486;
wire n_1897;
wire n_2984;
wire n_3646;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_3685;
wire n_811;
wire n_3097;
wire n_3507;
wire n_876;
wire n_791;
wire n_1191;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_3450;
wire n_2337;
wire n_2265;
wire n_2900;
wire n_797;
wire n_2026;
wire n_2912;
wire n_3524;
wire n_1786;
wire n_2627;
wire n_3173;
wire n_1327;
wire n_1475;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_3174;
wire n_3314;
wire n_2726;
wire n_2622;
wire n_3447;
wire n_2272;
wire n_3266;
wire n_1757;
wire n_3102;
wire n_1499;
wire n_854;
wire n_1318;
wire n_3452;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_2929;
wire n_3124;
wire n_3422;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_3411;
wire n_1526;
wire n_2991;
wire n_3463;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1873;
wire n_1137;
wire n_1258;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_2928;
wire n_943;
wire n_1118;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_3167;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_3110;
wire n_771;
wire n_1321;
wire n_3050;
wire n_3157;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_3142;
wire n_1984;
wire n_1350;
wire n_3453;
wire n_3129;
wire n_1556;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_3298;
wire n_3107;
wire n_3495;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_2700;
wire n_2606;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_2907;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_3543;
wire n_3640;
wire n_1776;
wire n_3448;
wire n_2936;
wire n_1154;
wire n_3609;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_2022;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2986;
wire n_2320;
wire n_3140;
wire n_979;
wire n_2329;
wire n_2570;
wire n_3017;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_2890;
wire n_2911;
wire n_3455;
wire n_807;
wire n_891;
wire n_3313;
wire n_885;
wire n_1659;
wire n_2354;
wire n_3591;
wire n_1864;
wire n_2760;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_1208;
wire n_3317;
wire n_3336;
wire n_1987;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_3635;
wire n_2352;
wire n_3541;
wire n_2502;
wire n_1256;
wire n_714;
wire n_3560;
wire n_3345;
wire n_2170;
wire n_3605;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_3566;
wire n_3421;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_3548;
wire n_2652;
wire n_1133;
wire n_3067;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_3236;
wire n_2222;
wire n_3468;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_3573;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_2943;
wire n_1426;
wire n_2250;
wire n_3319;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_3321;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_3291;
wire n_3654;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_3643;
wire n_2285;
wire n_3343;
wire n_3184;
wire n_3309;
wire n_2892;
wire n_1288;
wire n_1201;
wire n_2605;
wire n_2796;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2173;
wire n_2715;
wire n_3206;
wire n_3647;
wire n_1035;
wire n_3475;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_3134;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_2947;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_825;
wire n_1103;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_3098;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_3055;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_3341;
wire n_3600;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_3223;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_3386;
wire n_914;
wire n_1116;
wire n_3043;
wire n_3190;
wire n_1958;
wire n_2747;
wire n_3667;
wire n_3027;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_3462;
wire n_1197;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_2613;
wire n_3226;
wire n_1165;
wire n_3378;
wire n_2934;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_3444;
wire n_1128;
wire n_3141;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_3476;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3096;
wire n_2419;
wire n_1049;
wire n_3380;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_3238;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_3189;
wire n_3233;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_3175;
wire n_1440;
wire n_3289;
wire n_2666;
wire n_3322;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_2935;
wire n_715;
wire n_889;
wire n_3255;
wire n_1549;
wire n_1066;
wire n_2863;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2886;
wire n_2478;
wire n_911;
wire n_2658;
wire n_3509;
wire n_3587;
wire n_2608;
wire n_3620;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_1403;
wire n_1534;
wire n_1065;
wire n_1948;
wire n_3006;
wire n_2767;
wire n_810;
wire n_3381;
wire n_3376;
wire n_1290;
wire n_1959;
wire n_3497;
wire n_2396;
wire n_3243;
wire n_3368;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_3456;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_3117;
wire n_3595;
wire n_743;
wire n_1194;
wire n_2862;
wire n_1647;
wire n_1546;
wire n_3384;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_3490;
wire n_2459;
wire n_962;
wire n_941;
wire n_3396;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_3113;
wire n_3101;
wire n_1968;
wire n_918;
wire n_3307;
wire n_3662;
wire n_1885;
wire n_3288;
wire n_3251;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_3683;
wire n_3195;
wire n_3008;
wire n_1695;
wire n_3242;
wire n_2560;
wire n_1164;
wire n_3405;
wire n_2313;
wire n_3077;
wire n_1193;
wire n_3048;
wire n_3339;
wire n_1345;
wire n_3037;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_2963;
wire n_3532;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_3363;
wire n_3533;
wire n_1767;
wire n_1040;
wire n_3131;
wire n_1158;
wire n_3168;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_1749;
wire n_820;
wire n_1653;
wire n_872;
wire n_3409;
wire n_3522;
wire n_3583;
wire n_2882;
wire n_2303;
wire n_2669;
wire n_3540;
wire n_3241;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_3481;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_1814;
wire n_3689;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_2624;
wire n_3442;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_2938;
wire n_834;
wire n_3630;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_2803;
wire n_1756;
wire n_2887;
wire n_1606;
wire n_2189;
wire n_2648;
wire n_3305;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_3354;
wire n_1014;
wire n_724;
wire n_2204;
wire n_2931;
wire n_3433;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2977;
wire n_3106;
wire n_3597;
wire n_2199;
wire n_2881;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_3092;
wire n_3437;
wire n_2231;
wire n_2828;
wire n_1626;
wire n_3436;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_3553;
wire n_2305;
wire n_3645;
wire n_880;
wire n_793;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3304;
wire n_3574;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_3402;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_3247;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_2883;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_3406;
wire n_2951;
wire n_3664;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_3550;
wire n_2014;
wire n_975;
wire n_2974;
wire n_1645;
wire n_923;
wire n_1381;
wire n_1124;
wire n_2870;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_3686;
wire n_1326;
wire n_2889;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_3301;
wire n_981;
wire n_2910;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_2503;
wire n_2270;
wire n_3470;
wire n_3294;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_3610;
wire n_1204;
wire n_2865;
wire n_1554;
wire n_3279;
wire n_994;
wire n_2428;
wire n_2972;
wire n_2586;
wire n_2989;
wire n_1360;
wire n_973;
wire n_3178;
wire n_2858;
wire n_972;
wire n_3259;
wire n_2251;
wire n_2923;
wire n_3076;
wire n_2843;
wire n_3410;
wire n_856;
wire n_3100;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_3676;
wire n_1564;
wire n_2010;
wire n_3677;
wire n_1054;
wire n_1679;
wire n_3292;
wire n_3389;
wire n_2872;
wire n_2126;
wire n_3109;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_3125;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_3537;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_2941;
wire n_1411;
wire n_1359;
wire n_3079;
wire n_3638;
wire n_3269;
wire n_3536;
wire n_1721;
wire n_2564;
wire n_3558;
wire n_3576;
wire n_2591;
wire n_1445;
wire n_1317;
wire n_3034;
wire n_2050;
wire n_2197;
wire n_3502;
wire n_3248;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_3177;
wire n_3594;
wire n_1471;
wire n_2385;
wire n_3440;
wire n_2387;
wire n_1008;
wire n_3658;
wire n_3091;
wire n_1024;
wire n_830;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_3227;
wire n_3570;
wire n_3105;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_788;
wire n_908;
wire n_2639;
wire n_3521;
wire n_1036;
wire n_2169;
wire n_2985;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_3663;
wire n_2028;
wire n_1663;
wire n_919;
wire n_3114;
wire n_2901;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_3225;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_3621;
wire n_1458;
wire n_1630;
wire n_3473;
wire n_3644;
wire n_3047;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3163;
wire n_3680;
wire n_3431;
wire n_2176;
wire n_3565;
wire n_1412;
wire n_3355;
wire n_3059;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_3331;
wire n_1735;
wire n_1788;
wire n_940;
wire n_3520;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_3272;
wire n_3122;
wire n_3040;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_3360;
wire n_1930;
wire n_3687;
wire n_765;
wire n_1809;
wire n_2787;
wire n_3585;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_3211;
wire n_2395;
wire n_917;
wire n_2868;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_1170;
wire n_2724;
wire n_3575;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_3633;
wire n_857;
wire n_898;
wire n_3042;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_3278;
wire n_1462;
wire n_3328;
wire n_1937;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_3608;
wire n_1064;
wire n_900;
wire n_1446;
wire n_1282;
wire n_3004;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_3379;
wire n_3111;
wire n_761;
wire n_733;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_2997;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_3258;
wire n_2734;
wire n_2569;
wire n_758;
wire n_2252;
wire n_3598;
wire n_2111;
wire n_2420;
wire n_2948;
wire n_3099;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_816;
wire n_2897;
wire n_1322;
wire n_3273;
wire n_2583;
wire n_2918;
wire n_2987;
wire n_1473;
wire n_835;
wire n_3155;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_3316;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_3632;
wire n_2463;
wire n_3546;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2699;
wire n_2580;
wire n_1792;
wire n_3351;
wire n_2062;
wire n_3068;
wire n_1141;
wire n_3457;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_2973;
wire n_1459;
wire n_2153;
wire n_840;
wire n_2324;
wire n_1510;
wire n_3454;
wire n_3002;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_3146;
wire n_3394;
wire n_3038;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_3132;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_3581;
wire n_831;
wire n_3681;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3303;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_1902;
wire n_997;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_1643;
wire n_1320;
wire n_3188;
wire n_3001;
wire n_3232;
wire n_1113;
wire n_3218;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2990;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_3445;
wire n_1409;
wire n_1588;
wire n_1684;
wire n_1148;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_2290;
wire n_2933;
wire n_3253;
wire n_2856;
wire n_3235;
wire n_3387;
wire n_2088;
wire n_3265;
wire n_1275;
wire n_3103;
wire n_3018;
wire n_904;
wire n_2005;
wire n_3584;
wire n_2048;
wire n_1696;
wire n_3446;
wire n_3028;
wire n_1875;
wire n_1059;
wire n_3148;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_3285;
wire n_1039;
wire n_2246;
wire n_3616;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_2971;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1600;
wire n_1190;
wire n_1144;
wire n_3203;
wire n_838;
wire n_1558;
wire n_1941;
wire n_3628;
wire n_1316;
wire n_2519;
wire n_3637;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_1369;
wire n_2846;
wire n_3371;
wire n_1781;
wire n_709;
wire n_2917;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3143;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_3229;
wire n_3032;
wire n_1686;
wire n_1964;
wire n_3659;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_3461;
wire n_3366;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_1410;
wire n_939;
wire n_2297;
wire n_3094;
wire n_3441;
wire n_3020;
wire n_2964;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_2957;
wire n_865;
wire n_1273;
wire n_1983;
wire n_2982;
wire n_1041;
wire n_2451;
wire n_3312;
wire n_2115;
wire n_2913;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_3672;
wire n_922;
wire n_1004;
wire n_1810;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_1347;
wire n_2839;
wire n_3237;
wire n_860;
wire n_3555;
wire n_3072;
wire n_1043;
wire n_2961;
wire n_2869;
wire n_3534;
wire n_1923;
wire n_3655;
wire n_2955;
wire n_2670;
wire n_3631;
wire n_1764;
wire n_2674;
wire n_3556;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_3026;
wire n_2644;
wire n_902;
wire n_1031;
wire n_2979;
wire n_1723;
wire n_3674;
wire n_1638;
wire n_853;
wire n_3071;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_1946;
wire n_774;
wire n_933;
wire n_3244;
wire n_3499;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_3112;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_3296;
wire n_3196;
wire n_3593;
wire n_2673;
wire n_1591;
wire n_2585;
wire n_2995;
wire n_3361;
wire n_3293;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_3228;
wire n_3327;
wire n_2548;
wire n_3488;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_3149;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_3088;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_3590;
wire n_2058;
wire n_3231;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_2875;
wire n_1639;
wire n_3519;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_1000;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_2792;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_3398;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_3557;
wire n_3592;
wire n_2269;
wire n_2081;
wire n_1474;
wire n_937;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_3399;
wire n_3202;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_1232;
wire n_1211;
wire n_1368;
wire n_996;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2891;
wire n_2318;
wire n_1827;
wire n_3128;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1722;
wire n_1001;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_2880;
wire n_3075;
wire n_3030;
wire n_3505;
wire n_1339;
wire n_1644;
wire n_1002;
wire n_1051;
wire n_3547;
wire n_2551;
wire n_719;
wire n_1102;
wire n_2255;
wire n_1252;
wire n_2239;
wire n_1129;
wire n_3045;
wire n_1464;
wire n_1296;
wire n_3158;
wire n_773;
wire n_2798;
wire n_3221;
wire n_2316;
wire n_3217;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_3201;
wire n_3334;
wire n_2573;
wire n_2940;
wire n_3503;
wire n_3427;
wire n_2336;
wire n_1662;
wire n_3162;
wire n_1299;
wire n_1870;
wire n_3249;
wire n_3430;
wire n_3483;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2915;
wire n_3489;
wire n_3083;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_3213;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_3484;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2965;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2876;
wire n_2797;
wire n_3041;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_3080;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_3033;
wire n_1704;
wire n_893;
wire n_3525;
wire n_3308;
wire n_1582;
wire n_841;
wire n_2479;
wire n_3204;
wire n_886;
wire n_1981;
wire n_1069;
wire n_2824;
wire n_2037;
wire n_2953;
wire n_3428;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;

INVx1_ASAP7_75t_L g700 ( 
.A(n_304),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_413),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_52),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_380),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_597),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_28),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_539),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_281),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_358),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_503),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_657),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_620),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_456),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_637),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_653),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_689),
.Y(n_715)
);

CKINVDCx16_ASAP7_75t_R g716 ( 
.A(n_695),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_310),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_100),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_654),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_587),
.Y(n_720)
);

BUFx10_ASAP7_75t_L g721 ( 
.A(n_383),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_116),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_308),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_397),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_582),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_540),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_307),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_578),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_362),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_163),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_647),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_593),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_681),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_81),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_171),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_325),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_591),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_163),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_507),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_636),
.Y(n_740)
);

CKINVDCx16_ASAP7_75t_R g741 ( 
.A(n_592),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_678),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_506),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_214),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_186),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_440),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_398),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_698),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_696),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_299),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_435),
.Y(n_751)
);

BUFx2_ASAP7_75t_L g752 ( 
.A(n_687),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_353),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_317),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_91),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_660),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_659),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_55),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

CKINVDCx16_ASAP7_75t_R g760 ( 
.A(n_393),
.Y(n_760)
);

BUFx3_ASAP7_75t_L g761 ( 
.A(n_131),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_290),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_65),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_444),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_312),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_332),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_173),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_164),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_392),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_474),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_319),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_86),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_83),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_624),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_369),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_184),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_174),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_639),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_79),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_551),
.Y(n_780)
);

BUFx3_ASAP7_75t_L g781 ( 
.A(n_608),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_508),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_595),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_677),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_60),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_574),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_271),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_202),
.Y(n_788)
);

BUFx5_ASAP7_75t_L g789 ( 
.A(n_594),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_492),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_686),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_30),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_617),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_55),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_199),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_197),
.Y(n_796)
);

INVx1_ASAP7_75t_SL g797 ( 
.A(n_34),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_699),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_205),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_239),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_383),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_627),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_435),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_651),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_465),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_354),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_621),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_445),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_509),
.Y(n_809)
);

BUFx2_ASAP7_75t_L g810 ( 
.A(n_556),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_418),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_89),
.Y(n_812)
);

BUFx8_ASAP7_75t_SL g813 ( 
.A(n_641),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_454),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_478),
.Y(n_815)
);

INVx1_ASAP7_75t_SL g816 ( 
.A(n_557),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_19),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_175),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_135),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_614),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_622),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_607),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_643),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_7),
.Y(n_824)
);

CKINVDCx16_ASAP7_75t_R g825 ( 
.A(n_326),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_180),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_618),
.Y(n_827)
);

INVx2_ASAP7_75t_R g828 ( 
.A(n_250),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_609),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_664),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_605),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_509),
.Y(n_832)
);

BUFx10_ASAP7_75t_L g833 ( 
.A(n_575),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_272),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_488),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_191),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_255),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_288),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_119),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_652),
.Y(n_840)
);

CKINVDCx20_ASAP7_75t_R g841 ( 
.A(n_300),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_464),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_439),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_452),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_631),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_648),
.Y(n_846)
);

CKINVDCx20_ASAP7_75t_R g847 ( 
.A(n_417),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_172),
.Y(n_848)
);

CKINVDCx20_ASAP7_75t_R g849 ( 
.A(n_427),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_192),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_561),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_428),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_158),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_201),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_149),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_522),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_670),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_10),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_629),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_72),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_367),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_97),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_347),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_386),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_688),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_202),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_302),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_370),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_656),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_692),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_549),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_224),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_366),
.Y(n_873)
);

INVxp67_ASAP7_75t_L g874 ( 
.A(n_244),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_364),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_110),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_312),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_351),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_90),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_604),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_385),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_602),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_642),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_271),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_630),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_612),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_333),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_655),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_365),
.Y(n_889)
);

BUFx10_ASAP7_75t_L g890 ( 
.A(n_697),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_510),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_674),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_666),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_499),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_596),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_52),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_164),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_296),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_521),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_313),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_219),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_16),
.Y(n_902)
);

CKINVDCx20_ASAP7_75t_R g903 ( 
.A(n_531),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_662),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_159),
.Y(n_905)
);

CKINVDCx11_ASAP7_75t_R g906 ( 
.A(n_508),
.Y(n_906)
);

CKINVDCx20_ASAP7_75t_R g907 ( 
.A(n_451),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_570),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_667),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_471),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_168),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_682),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_385),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_320),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_264),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_84),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_303),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_638),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_183),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_487),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_10),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_690),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_419),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_443),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_467),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_366),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_599),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_489),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_542),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_193),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_298),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_468),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_534),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_103),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_573),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_684),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_548),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_356),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_436),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_126),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_632),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_13),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_669),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_184),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_396),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_691),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_22),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_113),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_514),
.Y(n_949)
);

INVx2_ASAP7_75t_SL g950 ( 
.A(n_276),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_320),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_255),
.Y(n_952)
);

INVx1_ASAP7_75t_SL g953 ( 
.A(n_186),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_215),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_672),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_409),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_245),
.Y(n_957)
);

CKINVDCx16_ASAP7_75t_R g958 ( 
.A(n_616),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_529),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_619),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_515),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_291),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_650),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_146),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_615),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_658),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_495),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_244),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_258),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_162),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_644),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_405),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_311),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_316),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_679),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_32),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_107),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_371),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_168),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_245),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_396),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_434),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_290),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_470),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_680),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_353),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_676),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_188),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_162),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_36),
.Y(n_990)
);

BUFx10_ASAP7_75t_L g991 ( 
.A(n_139),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_302),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_389),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_333),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_675),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_92),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_381),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_105),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_207),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_102),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_668),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_49),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_663),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_116),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_393),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_293),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_223),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_598),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_5),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_380),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_97),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_237),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_206),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_377),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_149),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_363),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_488),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_124),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_292),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_112),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_544),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_115),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_15),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_85),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_554),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_288),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_601),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_183),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_635),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_296),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_190),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_107),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_414),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_205),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_109),
.Y(n_1035)
);

BUFx3_ASAP7_75t_L g1036 ( 
.A(n_625),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_203),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_58),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_193),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_221),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_391),
.Y(n_1041)
);

INVx1_ASAP7_75t_SL g1042 ( 
.A(n_207),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_5),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_269),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_108),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_30),
.Y(n_1046)
);

INVx2_ASAP7_75t_SL g1047 ( 
.A(n_133),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_613),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_46),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_22),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_329),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_581),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_564),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_330),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_406),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_493),
.Y(n_1056)
);

BUFx5_ASAP7_75t_L g1057 ( 
.A(n_425),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_123),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_512),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_217),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_513),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_72),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_417),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_231),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_420),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_17),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_507),
.Y(n_1067)
);

INVxp33_ASAP7_75t_L g1068 ( 
.A(n_633),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_196),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_449),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_215),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_464),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_213),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_176),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_409),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_398),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_1),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_153),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_279),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_572),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_538),
.Y(n_1081)
);

INVx1_ASAP7_75t_SL g1082 ( 
.A(n_50),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_39),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_490),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_130),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_246),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_426),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_83),
.Y(n_1088)
);

CKINVDCx20_ASAP7_75t_R g1089 ( 
.A(n_217),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_44),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_73),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_155),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_3),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_175),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_423),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_673),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_480),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_571),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_44),
.Y(n_1099)
);

CKINVDCx16_ASAP7_75t_R g1100 ( 
.A(n_142),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_66),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_423),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_513),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_368),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_603),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_178),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_580),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_665),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_9),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_289),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_338),
.Y(n_1111)
);

CKINVDCx16_ASAP7_75t_R g1112 ( 
.A(n_555),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_27),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_210),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_73),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_98),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_306),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_64),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_405),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_355),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_541),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_470),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_293),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_661),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_94),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_685),
.Y(n_1126)
);

CKINVDCx20_ASAP7_75t_R g1127 ( 
.A(n_279),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_261),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_628),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_693),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_514),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_16),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_98),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_437),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_611),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_487),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_407),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_606),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_503),
.Y(n_1139)
);

CKINVDCx16_ASAP7_75t_R g1140 ( 
.A(n_345),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_154),
.Y(n_1141)
);

CKINVDCx14_ASAP7_75t_R g1142 ( 
.A(n_273),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_118),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_256),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_25),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_558),
.Y(n_1146)
);

INVx1_ASAP7_75t_SL g1147 ( 
.A(n_339),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_204),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_634),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_199),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_442),
.Y(n_1151)
);

INVx1_ASAP7_75t_SL g1152 ( 
.A(n_527),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_79),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_475),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_683),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_136),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_553),
.Y(n_1157)
);

INVx2_ASAP7_75t_SL g1158 ( 
.A(n_63),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_89),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_392),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_406),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_350),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_219),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_332),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_588),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_649),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_586),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_590),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_349),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_144),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_70),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_323),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_671),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_623),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_452),
.Y(n_1175)
);

BUFx2_ASAP7_75t_SL g1176 ( 
.A(n_147),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_54),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_324),
.Y(n_1178)
);

CKINVDCx20_ASAP7_75t_R g1179 ( 
.A(n_237),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_402),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_413),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_530),
.Y(n_1182)
);

INVx2_ASAP7_75t_SL g1183 ( 
.A(n_246),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_640),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_189),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_511),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_235),
.Y(n_1187)
);

BUFx5_ASAP7_75t_L g1188 ( 
.A(n_455),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_407),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_254),
.Y(n_1190)
);

INVx2_ASAP7_75t_SL g1191 ( 
.A(n_359),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_157),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_93),
.Y(n_1193)
);

CKINVDCx20_ASAP7_75t_R g1194 ( 
.A(n_447),
.Y(n_1194)
);

CKINVDCx20_ASAP7_75t_R g1195 ( 
.A(n_128),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_33),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_584),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_432),
.Y(n_1198)
);

CKINVDCx16_ASAP7_75t_R g1199 ( 
.A(n_600),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_646),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_610),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_694),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_626),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_11),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_70),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_425),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_569),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_467),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_378),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_395),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_63),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_537),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_645),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_270),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_781),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_761),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_761),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_776),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_776),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_770),
.Y(n_1220)
);

CKINVDCx16_ASAP7_75t_R g1221 ( 
.A(n_1142),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_803),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_803),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_809),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_906),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_809),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_834),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_837),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_752),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_837),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_852),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_852),
.Y(n_1232)
);

CKINVDCx20_ASAP7_75t_R g1233 ( 
.A(n_1142),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_902),
.Y(n_1234)
);

CKINVDCx20_ASAP7_75t_R g1235 ( 
.A(n_731),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_906),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_902),
.Y(n_1237)
);

CKINVDCx20_ASAP7_75t_R g1238 ( 
.A(n_731),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1007),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1007),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1134),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_770),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_810),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1163),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1163),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_770),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_770),
.Y(n_1248)
);

NOR2xp67_ASAP7_75t_L g1249 ( 
.A(n_911),
.B(n_0),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_770),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_770),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_770),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1057),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_813),
.Y(n_1254)
);

CKINVDCx16_ASAP7_75t_R g1255 ( 
.A(n_760),
.Y(n_1255)
);

INVxp33_ASAP7_75t_SL g1256 ( 
.A(n_824),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1057),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1057),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1057),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1057),
.Y(n_1260)
);

INVxp67_ASAP7_75t_SL g1261 ( 
.A(n_735),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1057),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_813),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_727),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1057),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1188),
.Y(n_1266)
);

INVx1_ASAP7_75t_SL g1267 ( 
.A(n_841),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1188),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_825),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1188),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1188),
.Y(n_1271)
);

INVxp33_ASAP7_75t_L g1272 ( 
.A(n_972),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1188),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1188),
.Y(n_1274)
);

HB1xp67_ASAP7_75t_L g1275 ( 
.A(n_1014),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_727),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1188),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_805),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1068),
.B(n_706),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_867),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_700),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_746),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1086),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_1009),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_701),
.Y(n_1285)
);

CKINVDCx16_ASAP7_75t_R g1286 ( 
.A(n_1100),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_705),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1140),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_707),
.Y(n_1289)
);

INVxp33_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_718),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_746),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_1127),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_723),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_724),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_729),
.Y(n_1296)
);

INVxp67_ASAP7_75t_L g1297 ( 
.A(n_735),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_747),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_755),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_768),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_784),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_784),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_769),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_771),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_798),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_775),
.Y(n_1306)
);

INVx2_ASAP7_75t_L g1307 ( 
.A(n_805),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_788),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_795),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_808),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_805),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_845),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_812),
.Y(n_1313)
);

BUFx3_ASAP7_75t_L g1314 ( 
.A(n_833),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_754),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_817),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_754),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_835),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_836),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_854),
.Y(n_1320)
);

INVxp33_ASAP7_75t_SL g1321 ( 
.A(n_1176),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_855),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_782),
.Y(n_1323)
);

INVxp67_ASAP7_75t_SL g1324 ( 
.A(n_782),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_833),
.Y(n_1325)
);

CKINVDCx16_ASAP7_75t_R g1326 ( 
.A(n_716),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_858),
.Y(n_1327)
);

CKINVDCx16_ASAP7_75t_R g1328 ( 
.A(n_741),
.Y(n_1328)
);

INVxp33_ASAP7_75t_L g1329 ( 
.A(n_799),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_861),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_866),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_833),
.Y(n_1332)
);

INVxp67_ASAP7_75t_SL g1333 ( 
.A(n_799),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_878),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_890),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_702),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_889),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_894),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_703),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_708),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_897),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_900),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_910),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_SL g1344 ( 
.A(n_890),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_913),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_915),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_890),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_923),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_939),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_709),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1247),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1248),
.Y(n_1352)
);

BUFx12f_ASAP7_75t_L g1353 ( 
.A(n_1254),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1215),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1278),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1307),
.Y(n_1356)
);

CKINVDCx20_ASAP7_75t_R g1357 ( 
.A(n_1235),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1311),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1279),
.B(n_958),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1344),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1312),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_1215),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1221),
.B(n_975),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1220),
.Y(n_1364)
);

INVx5_ASAP7_75t_L g1365 ( 
.A(n_1215),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1250),
.Y(n_1366)
);

BUFx6f_ASAP7_75t_L g1367 ( 
.A(n_1215),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1251),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1252),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_1243),
.Y(n_1370)
);

CKINVDCx16_ASAP7_75t_R g1371 ( 
.A(n_1326),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1258),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1279),
.B(n_1112),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1253),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1257),
.A2(n_783),
.B(n_719),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1259),
.Y(n_1377)
);

AND2x4_ASAP7_75t_L g1378 ( 
.A(n_1314),
.B(n_884),
.Y(n_1378)
);

BUFx6f_ASAP7_75t_L g1379 ( 
.A(n_1270),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_1273),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1260),
.Y(n_1381)
);

BUFx6f_ASAP7_75t_L g1382 ( 
.A(n_1262),
.Y(n_1382)
);

BUFx12f_ASAP7_75t_L g1383 ( 
.A(n_1263),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1225),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1329),
.B(n_1199),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1269),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1265),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1266),
.Y(n_1388)
);

OAI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1256),
.A2(n_847),
.B1(n_849),
.B2(n_796),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1271),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1274),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1216),
.Y(n_1392)
);

BUFx6f_ASAP7_75t_L g1393 ( 
.A(n_1277),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1217),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_L g1395 ( 
.A(n_1280),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1218),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1219),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1222),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1281),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1223),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1285),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1287),
.Y(n_1402)
);

INVx3_ASAP7_75t_L g1403 ( 
.A(n_1224),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1325),
.B(n_1068),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1226),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1289),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1228),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1291),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1238),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1332),
.B(n_711),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1335),
.B(n_714),
.Y(n_1411)
);

INVx4_ASAP7_75t_L g1412 ( 
.A(n_1344),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1230),
.Y(n_1413)
);

BUFx6f_ASAP7_75t_L g1414 ( 
.A(n_1294),
.Y(n_1414)
);

OA21x2_ASAP7_75t_L g1415 ( 
.A1(n_1295),
.A2(n_783),
.B(n_719),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1296),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1231),
.Y(n_1417)
);

BUFx6f_ASAP7_75t_L g1418 ( 
.A(n_1298),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1283),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1299),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1329),
.B(n_721),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1301),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1300),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1232),
.Y(n_1424)
);

BUFx6f_ASAP7_75t_L g1425 ( 
.A(n_1303),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1304),
.Y(n_1426)
);

AOI22x1_ASAP7_75t_SL g1427 ( 
.A1(n_1264),
.A2(n_847),
.B1(n_849),
.B2(n_796),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1306),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1234),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1347),
.B(n_721),
.Y(n_1430)
);

AND2x6_ASAP7_75t_L g1431 ( 
.A(n_1237),
.B(n_781),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1308),
.A2(n_1149),
.B(n_880),
.Y(n_1432)
);

CKINVDCx6p67_ASAP7_75t_R g1433 ( 
.A(n_1328),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1272),
.A2(n_857),
.B1(n_870),
.B2(n_798),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_1302),
.Y(n_1435)
);

BUFx6f_ASAP7_75t_L g1436 ( 
.A(n_1309),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1239),
.B(n_720),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1240),
.A2(n_733),
.B(n_726),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1310),
.A2(n_1149),
.B(n_880),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1313),
.A2(n_1168),
.B(n_1157),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1241),
.B(n_749),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1316),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1242),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1318),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1245),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1229),
.B(n_884),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1272),
.B(n_721),
.Y(n_1447)
);

BUFx2_ASAP7_75t_L g1448 ( 
.A(n_1284),
.Y(n_1448)
);

BUFx12f_ASAP7_75t_L g1449 ( 
.A(n_1236),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1246),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1319),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1320),
.Y(n_1452)
);

AOI22x1_ASAP7_75t_SL g1453 ( 
.A1(n_1264),
.A2(n_863),
.B1(n_879),
.B2(n_853),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1290),
.B(n_991),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1322),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1327),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1330),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1331),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1244),
.B(n_896),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1334),
.Y(n_1460)
);

BUFx12f_ASAP7_75t_L g1461 ( 
.A(n_1288),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1337),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1338),
.A2(n_807),
.B(n_759),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1336),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1339),
.Y(n_1465)
);

OA21x2_ASAP7_75t_L g1466 ( 
.A1(n_1341),
.A2(n_1168),
.B(n_1157),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1342),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1340),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1343),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1345),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_1305),
.Y(n_1471)
);

CKINVDCx5p33_ASAP7_75t_R g1472 ( 
.A(n_1267),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1346),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1362),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1396),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1472),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1362),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1397),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1405),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1351),
.B(n_1261),
.Y(n_1480)
);

INVxp67_ASAP7_75t_L g1481 ( 
.A(n_1385),
.Y(n_1481)
);

BUFx2_ASAP7_75t_L g1482 ( 
.A(n_1361),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1447),
.Y(n_1483)
);

AND2x6_ASAP7_75t_L g1484 ( 
.A(n_1421),
.B(n_856),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1354),
.Y(n_1485)
);

INVx3_ASAP7_75t_L g1486 ( 
.A(n_1362),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1351),
.B(n_1261),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1367),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1367),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1352),
.B(n_1366),
.Y(n_1490)
);

AOI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1359),
.A2(n_1374),
.B1(n_857),
.B2(n_882),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1407),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1413),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1367),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1352),
.B(n_1324),
.Y(n_1495)
);

AND2x4_ASAP7_75t_L g1496 ( 
.A(n_1430),
.B(n_1324),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1372),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1372),
.Y(n_1498)
);

BUFx6f_ASAP7_75t_L g1499 ( 
.A(n_1372),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1454),
.A2(n_882),
.B1(n_903),
.B2(n_870),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1417),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1379),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1424),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1378),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1463),
.A2(n_831),
.B(n_830),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1379),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1429),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1443),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_1401),
.B(n_856),
.Y(n_1509)
);

NOR2xp33_ASAP7_75t_L g1510 ( 
.A(n_1366),
.B(n_1321),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1379),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1380),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1380),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1380),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1445),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1378),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1382),
.B(n_1350),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1450),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1370),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1370),
.Y(n_1520)
);

AND2x4_ASAP7_75t_L g1521 ( 
.A(n_1446),
.B(n_1333),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1382),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1451),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1456),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1382),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1368),
.B(n_1333),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1390),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1390),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1390),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1368),
.B(n_1348),
.Y(n_1530)
);

INVxp33_ASAP7_75t_SL g1531 ( 
.A(n_1386),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1391),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1391),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1457),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1468),
.B(n_1290),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1391),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1393),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1393),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1393),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1355),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1356),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1358),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1369),
.B(n_1349),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1448),
.B(n_1255),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1401),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1402),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1414),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1404),
.B(n_1286),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1402),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1364),
.Y(n_1550)
);

NAND2xp33_ASAP7_75t_SL g1551 ( 
.A(n_1464),
.B(n_903),
.Y(n_1551)
);

BUFx6f_ASAP7_75t_L g1552 ( 
.A(n_1414),
.Y(n_1552)
);

OA21x2_ASAP7_75t_L g1553 ( 
.A1(n_1438),
.A2(n_885),
.B(n_846),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1406),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1465),
.B(n_1275),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1406),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1408),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1408),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1373),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1416),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1416),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1381),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1446),
.B(n_1297),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_SL g1564 ( 
.A(n_1369),
.B(n_893),
.Y(n_1564)
);

AND2x6_ASAP7_75t_L g1565 ( 
.A(n_1420),
.B(n_1473),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1420),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_R g1567 ( 
.A(n_1409),
.B(n_1233),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1444),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1414),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1418),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1444),
.Y(n_1571)
);

NAND2xp33_ASAP7_75t_R g1572 ( 
.A(n_1422),
.B(n_712),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1435),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1473),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1395),
.B(n_1275),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1371),
.B(n_1293),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1375),
.Y(n_1577)
);

BUFx8_ASAP7_75t_L g1578 ( 
.A(n_1384),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1375),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1377),
.B(n_912),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1377),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1387),
.B(n_929),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1387),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1388),
.Y(n_1584)
);

INVx3_ASAP7_75t_L g1585 ( 
.A(n_1418),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1388),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1399),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1461),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1418),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1425),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1425),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1425),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1426),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1423),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1426),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1426),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1459),
.B(n_1227),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1428),
.Y(n_1598)
);

NOR2xp33_ASAP7_75t_L g1599 ( 
.A(n_1410),
.B(n_1297),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1442),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1459),
.B(n_1227),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1353),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1469),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1455),
.B(n_1323),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1470),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1392),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1392),
.Y(n_1607)
);

INVx1_ASAP7_75t_SL g1608 ( 
.A(n_1576),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1521),
.B(n_1412),
.Y(n_1609)
);

INVx3_ASAP7_75t_L g1610 ( 
.A(n_1476),
.Y(n_1610)
);

INVxp67_ASAP7_75t_SL g1611 ( 
.A(n_1537),
.Y(n_1611)
);

BUFx10_ASAP7_75t_L g1612 ( 
.A(n_1573),
.Y(n_1612)
);

INVx5_ASAP7_75t_L g1613 ( 
.A(n_1565),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_SL g1614 ( 
.A(n_1481),
.B(n_1412),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1519),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1602),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1579),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1481),
.A2(n_904),
.B1(n_1105),
.B2(n_909),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1510),
.A2(n_1491),
.B1(n_1483),
.B2(n_1581),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1520),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1540),
.Y(n_1622)
);

BUFx6f_ASAP7_75t_L g1623 ( 
.A(n_1552),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1599),
.B(n_1431),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1599),
.B(n_1431),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1535),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1491),
.A2(n_828),
.B1(n_1431),
.B2(n_1389),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1544),
.Y(n_1628)
);

NOR3xp33_ASAP7_75t_SL g1629 ( 
.A(n_1572),
.B(n_722),
.C(n_717),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1531),
.B(n_1383),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1575),
.B(n_1471),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1583),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1584),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1510),
.B(n_1411),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1541),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1542),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1604),
.B(n_1431),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1482),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1496),
.B(n_1455),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1555),
.B(n_1434),
.Y(n_1640)
);

BUFx10_ASAP7_75t_L g1641 ( 
.A(n_1496),
.Y(n_1641)
);

CKINVDCx20_ASAP7_75t_R g1642 ( 
.A(n_1588),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1586),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1545),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1563),
.B(n_1449),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1563),
.B(n_1433),
.Y(n_1646)
);

INVx3_ASAP7_75t_L g1647 ( 
.A(n_1552),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1530),
.B(n_1462),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1483),
.B(n_1363),
.Y(n_1649)
);

AND2x6_ASAP7_75t_L g1650 ( 
.A(n_1546),
.B(n_1394),
.Y(n_1650)
);

AND2x6_ASAP7_75t_L g1651 ( 
.A(n_1549),
.B(n_1394),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1550),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1548),
.B(n_1436),
.C(n_1428),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1597),
.B(n_1360),
.Y(n_1654)
);

XNOR2xp5_ASAP7_75t_L g1655 ( 
.A(n_1500),
.B(n_1276),
.Y(n_1655)
);

AND2x6_ASAP7_75t_L g1656 ( 
.A(n_1554),
.B(n_1398),
.Y(n_1656)
);

AND2x6_ASAP7_75t_L g1657 ( 
.A(n_1556),
.B(n_1398),
.Y(n_1657)
);

NAND3xp33_ASAP7_75t_L g1658 ( 
.A(n_1551),
.B(n_1436),
.C(n_1428),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1601),
.Y(n_1659)
);

AO22x2_ASAP7_75t_L g1660 ( 
.A1(n_1500),
.A2(n_1453),
.B1(n_1427),
.B2(n_1282),
.Y(n_1660)
);

BUFx6f_ASAP7_75t_L g1661 ( 
.A(n_1552),
.Y(n_1661)
);

INVx4_ASAP7_75t_L g1662 ( 
.A(n_1565),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1557),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1572),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1558),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1551),
.A2(n_828),
.B1(n_1432),
.B2(n_1415),
.Y(n_1666)
);

NOR2x1p5_ASAP7_75t_L g1667 ( 
.A(n_1578),
.B(n_1462),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1521),
.B(n_1400),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1530),
.B(n_1543),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1560),
.Y(n_1670)
);

INVx4_ASAP7_75t_L g1671 ( 
.A(n_1565),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1559),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_1517),
.B(n_1357),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1517),
.B(n_1276),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_1504),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_L g1676 ( 
.A(n_1565),
.B(n_805),
.Y(n_1676)
);

INVx4_ASAP7_75t_L g1677 ( 
.A(n_1569),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1561),
.Y(n_1678)
);

NOR2xp33_ASAP7_75t_L g1679 ( 
.A(n_1504),
.B(n_1282),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1516),
.B(n_1400),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1484),
.A2(n_1415),
.B1(n_1439),
.B2(n_1432),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1516),
.B(n_1292),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1606),
.B(n_1292),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1484),
.A2(n_909),
.B1(n_1105),
.B2(n_904),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1566),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_SL g1686 ( 
.A(n_1569),
.B(n_1589),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1607),
.B(n_1315),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1568),
.Y(n_1688)
);

INVx4_ASAP7_75t_L g1689 ( 
.A(n_1569),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1571),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1543),
.B(n_1452),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_L g1692 ( 
.A(n_1480),
.B(n_1315),
.Y(n_1692)
);

INVx3_ASAP7_75t_L g1693 ( 
.A(n_1589),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1574),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1480),
.B(n_1452),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1567),
.Y(n_1696)
);

BUFx3_ASAP7_75t_L g1697 ( 
.A(n_1578),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1523),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_1562),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_SL g1700 ( 
.A(n_1589),
.B(n_1452),
.Y(n_1700)
);

INVx4_ASAP7_75t_L g1701 ( 
.A(n_1484),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1475),
.Y(n_1702)
);

INVx4_ASAP7_75t_L g1703 ( 
.A(n_1484),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1478),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1479),
.Y(n_1705)
);

NAND3xp33_ASAP7_75t_L g1706 ( 
.A(n_1487),
.B(n_1458),
.C(n_1436),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1492),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1487),
.B(n_1458),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1587),
.A2(n_1440),
.B1(n_1466),
.B2(n_1439),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1493),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1495),
.B(n_1460),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1490),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1495),
.B(n_1458),
.Y(n_1713)
);

INVx3_ASAP7_75t_L g1714 ( 
.A(n_1547),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1501),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1503),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1507),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1508),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1526),
.B(n_1317),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_SL g1721 ( 
.A(n_1547),
.B(n_1467),
.Y(n_1721)
);

INVx1_ASAP7_75t_SL g1722 ( 
.A(n_1585),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1594),
.B(n_1460),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1585),
.B(n_1598),
.Y(n_1724)
);

INVxp33_ASAP7_75t_L g1725 ( 
.A(n_1567),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1515),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1518),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_L g1728 ( 
.A(n_1598),
.B(n_1317),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1600),
.B(n_1467),
.Y(n_1729)
);

AND2x6_ASAP7_75t_L g1730 ( 
.A(n_1603),
.B(n_1403),
.Y(n_1730)
);

AND2x6_ASAP7_75t_L g1731 ( 
.A(n_1605),
.B(n_1403),
.Y(n_1731)
);

BUFx6f_ASAP7_75t_L g1732 ( 
.A(n_1497),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1485),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1524),
.B(n_1467),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1490),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1537),
.B(n_1200),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1534),
.B(n_1437),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1497),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1537),
.B(n_1200),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1580),
.Y(n_1740)
);

INVx5_ASAP7_75t_L g1741 ( 
.A(n_1509),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1509),
.Y(n_1742)
);

AND3x2_ASAP7_75t_L g1743 ( 
.A(n_1570),
.B(n_1453),
.C(n_1427),
.Y(n_1743)
);

AOI22xp33_ASAP7_75t_L g1744 ( 
.A1(n_1564),
.A2(n_1466),
.B1(n_1440),
.B2(n_1376),
.Y(n_1744)
);

INVx2_ASAP7_75t_SL g1745 ( 
.A(n_1590),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_R g1746 ( 
.A(n_1486),
.B(n_1419),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1591),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1592),
.B(n_1441),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1580),
.B(n_1323),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1593),
.Y(n_1750)
);

AND3x4_ASAP7_75t_L g1751 ( 
.A(n_1595),
.B(n_1249),
.C(n_863),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1497),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1596),
.B(n_942),
.Y(n_1753)
);

BUFx3_ASAP7_75t_L g1754 ( 
.A(n_1486),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1522),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1499),
.Y(n_1756)
);

AOI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1564),
.A2(n_1376),
.B1(n_879),
.B2(n_907),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1499),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1499),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1525),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1527),
.B(n_772),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1528),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1529),
.Y(n_1763)
);

AND2x6_ASAP7_75t_L g1764 ( 
.A(n_1532),
.B(n_1008),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1513),
.Y(n_1765)
);

INVx4_ASAP7_75t_SL g1766 ( 
.A(n_1509),
.Y(n_1766)
);

BUFx8_ASAP7_75t_SL g1767 ( 
.A(n_1474),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1669),
.B(n_1509),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_SL g1769 ( 
.A(n_1613),
.B(n_1513),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1712),
.B(n_1582),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1735),
.B(n_1582),
.Y(n_1771)
);

AOI22x1_ASAP7_75t_SL g1772 ( 
.A1(n_1642),
.A2(n_907),
.B1(n_934),
.B2(n_853),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1740),
.B(n_1648),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1617),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1622),
.Y(n_1775)
);

AOI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1620),
.A2(n_1649),
.B1(n_1720),
.B2(n_1692),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1749),
.B(n_1533),
.Y(n_1777)
);

AOI22xp33_ASAP7_75t_L g1778 ( 
.A1(n_1627),
.A2(n_957),
.B1(n_1010),
.B2(n_934),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1634),
.B(n_1536),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1640),
.B(n_787),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1618),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1664),
.B(n_1419),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1632),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1613),
.B(n_1513),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1635),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1613),
.B(n_1538),
.Y(n_1786)
);

AND2x6_ASAP7_75t_SL g1787 ( 
.A(n_1645),
.B(n_948),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_SL g1788 ( 
.A(n_1662),
.B(n_1539),
.Y(n_1788)
);

INVx4_ASAP7_75t_L g1789 ( 
.A(n_1767),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1619),
.A2(n_1010),
.B1(n_1017),
.B2(n_957),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1636),
.Y(n_1791)
);

AOI21xp5_ASAP7_75t_L g1792 ( 
.A1(n_1624),
.A2(n_1505),
.B(n_1502),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1639),
.B(n_1691),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_L g1794 ( 
.A(n_1650),
.B(n_1498),
.Y(n_1794)
);

NOR2xp67_ASAP7_75t_L g1795 ( 
.A(n_1610),
.B(n_1488),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1633),
.Y(n_1796)
);

INVx2_ASAP7_75t_SL g1797 ( 
.A(n_1638),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1695),
.B(n_1506),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1652),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1643),
.Y(n_1800)
);

NAND2xp33_ASAP7_75t_L g1801 ( 
.A(n_1650),
.B(n_1511),
.Y(n_1801)
);

OA21x2_ASAP7_75t_L g1802 ( 
.A1(n_1681),
.A2(n_1514),
.B(n_1512),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1713),
.B(n_1488),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1716),
.B(n_1489),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1644),
.B(n_1494),
.Y(n_1805)
);

INVxp67_ASAP7_75t_L g1806 ( 
.A(n_1626),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1663),
.B(n_1474),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1671),
.B(n_1474),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1626),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_SL g1810 ( 
.A(n_1609),
.B(n_1477),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1672),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1665),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1670),
.B(n_1477),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1609),
.B(n_1477),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1628),
.B(n_1017),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1699),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1684),
.A2(n_1032),
.B1(n_1043),
.B2(n_1019),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1631),
.B(n_1211),
.C(n_874),
.Y(n_1818)
);

AOI22xp33_ASAP7_75t_L g1819 ( 
.A1(n_1757),
.A2(n_1032),
.B1(n_1043),
.B2(n_1019),
.Y(n_1819)
);

OAI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1630),
.A2(n_1668),
.B1(n_1659),
.B2(n_1680),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1674),
.A2(n_1179),
.B1(n_1194),
.B2(n_1089),
.Y(n_1821)
);

BUFx5_ASAP7_75t_L g1822 ( 
.A(n_1650),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1678),
.B(n_797),
.Y(n_1823)
);

INVx8_ASAP7_75t_L g1824 ( 
.A(n_1645),
.Y(n_1824)
);

NAND3xp33_ASAP7_75t_L g1825 ( 
.A(n_1683),
.B(n_1179),
.C(n_1089),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1615),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1685),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1688),
.Y(n_1828)
);

OR2x6_ASAP7_75t_L g1829 ( 
.A(n_1616),
.B(n_753),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1687),
.B(n_1614),
.C(n_1673),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1690),
.Y(n_1831)
);

NOR3xp33_ASAP7_75t_L g1832 ( 
.A(n_1679),
.B(n_1682),
.C(n_1728),
.Y(n_1832)
);

OAI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1625),
.A2(n_1195),
.B1(n_1194),
.B2(n_734),
.Y(n_1833)
);

BUFx6f_ASAP7_75t_SL g1834 ( 
.A(n_1697),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1694),
.B(n_843),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1725),
.B(n_1675),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1723),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1646),
.B(n_1195),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1641),
.B(n_1365),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1616),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1729),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1722),
.B(n_1612),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1637),
.A2(n_736),
.B1(n_738),
.B2(n_730),
.Y(n_1843)
);

NAND2xp33_ASAP7_75t_L g1844 ( 
.A(n_1651),
.B(n_739),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1737),
.B(n_862),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1608),
.B(n_991),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1730),
.B(n_953),
.Y(n_1847)
);

NAND2x1_ASAP7_75t_L g1848 ( 
.A(n_1651),
.B(n_1553),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1730),
.B(n_1030),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_SL g1850 ( 
.A(n_1623),
.B(n_1365),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1730),
.B(n_1731),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1621),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1667),
.B(n_838),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1623),
.B(n_1365),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1736),
.B(n_1042),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_1654),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_1746),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1661),
.B(n_743),
.Y(n_1858)
);

A2O1A1Ixp33_ASAP7_75t_L g1859 ( 
.A1(n_1676),
.A2(n_943),
.B(n_960),
.C(n_937),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1696),
.Y(n_1860)
);

OAI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1701),
.A2(n_745),
.B1(n_750),
.B2(n_744),
.Y(n_1861)
);

NOR2xp33_ASAP7_75t_L g1862 ( 
.A(n_1739),
.B(n_1082),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1731),
.B(n_1147),
.Y(n_1863)
);

NOR2xp33_ASAP7_75t_L g1864 ( 
.A(n_1653),
.B(n_751),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1661),
.B(n_758),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1761),
.Y(n_1866)
);

OR2x6_ASAP7_75t_L g1867 ( 
.A(n_1660),
.B(n_1658),
.Y(n_1867)
);

INVx2_ASAP7_75t_SL g1868 ( 
.A(n_1698),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1766),
.B(n_949),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1731),
.B(n_896),
.Y(n_1870)
);

INVx2_ASAP7_75t_SL g1871 ( 
.A(n_1753),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1748),
.B(n_920),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_SL g1873 ( 
.A(n_1703),
.B(n_762),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1651),
.B(n_920),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1753),
.Y(n_1875)
);

CKINVDCx11_ASAP7_75t_R g1876 ( 
.A(n_1732),
.Y(n_1876)
);

INVxp67_ASAP7_75t_L g1877 ( 
.A(n_1655),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1702),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1733),
.B(n_763),
.Y(n_1879)
);

INVx2_ASAP7_75t_SL g1880 ( 
.A(n_1754),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1656),
.B(n_994),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1656),
.B(n_994),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1655),
.B(n_991),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1656),
.B(n_1070),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1660),
.B(n_1139),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_SL g1886 ( 
.A(n_1751),
.B(n_1139),
.Y(n_1886)
);

OAI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1741),
.A2(n_1037),
.B1(n_1047),
.B2(n_950),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1714),
.B(n_1206),
.C(n_1158),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1766),
.B(n_968),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1657),
.B(n_1070),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1741),
.B(n_764),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1704),
.B(n_765),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1705),
.B(n_766),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1707),
.Y(n_1894)
);

AND2x6_ASAP7_75t_SL g1895 ( 
.A(n_1724),
.B(n_970),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1710),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1657),
.B(n_1071),
.Y(n_1897)
);

AOI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1657),
.A2(n_1734),
.B1(n_1711),
.B2(n_1708),
.Y(n_1898)
);

AO22x2_ASAP7_75t_L g1899 ( 
.A1(n_1715),
.A2(n_1183),
.B1(n_1191),
.B2(n_1066),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1717),
.B(n_1718),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1719),
.B(n_1071),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1726),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1629),
.B(n_1139),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1727),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1666),
.B(n_1091),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1741),
.B(n_767),
.Y(n_1906)
);

OR2x2_ASAP7_75t_L g1907 ( 
.A(n_1747),
.B(n_1750),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1755),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1760),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1762),
.B(n_976),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_SL g1911 ( 
.A(n_1732),
.B(n_773),
.Y(n_1911)
);

INVx2_ASAP7_75t_L g1912 ( 
.A(n_1763),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1756),
.B(n_777),
.Y(n_1913)
);

INVx2_ASAP7_75t_SL g1914 ( 
.A(n_1756),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1745),
.B(n_1091),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1647),
.B(n_1170),
.Y(n_1916)
);

NAND2xp5_ASAP7_75t_L g1917 ( 
.A(n_1693),
.B(n_1170),
.Y(n_1917)
);

NAND2xp33_ASAP7_75t_L g1918 ( 
.A(n_1765),
.B(n_779),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1738),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1706),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1721),
.B(n_978),
.Y(n_1921)
);

AOI22xp33_ASAP7_75t_L g1922 ( 
.A1(n_1742),
.A2(n_993),
.B1(n_998),
.B2(n_988),
.Y(n_1922)
);

INVxp67_ASAP7_75t_SL g1923 ( 
.A(n_1765),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1752),
.B(n_785),
.Y(n_1924)
);

NAND2x1_ASAP7_75t_L g1925 ( 
.A(n_1677),
.B(n_1553),
.Y(n_1925)
);

AO22x2_ASAP7_75t_L g1926 ( 
.A1(n_1743),
.A2(n_1002),
.B1(n_1005),
.B2(n_1000),
.Y(n_1926)
);

NAND3xp33_ASAP7_75t_L g1927 ( 
.A(n_1689),
.B(n_832),
.C(n_819),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1742),
.A2(n_1018),
.B1(n_1024),
.B2(n_1006),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1758),
.B(n_790),
.Y(n_1929)
);

O2A1O1Ixp33_ASAP7_75t_L g1930 ( 
.A1(n_1700),
.A2(n_1033),
.B(n_1035),
.C(n_1028),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1764),
.A2(n_1039),
.B1(n_1040),
.B2(n_1038),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_SL g1932 ( 
.A(n_1759),
.B(n_792),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1611),
.B(n_1686),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1764),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_SL g1935 ( 
.A(n_1709),
.B(n_794),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1776),
.B(n_1773),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1836),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1876),
.Y(n_1938)
);

AO21x2_ASAP7_75t_L g1939 ( 
.A1(n_1935),
.A2(n_1744),
.B(n_987),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1857),
.B(n_1764),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1866),
.B(n_800),
.Y(n_1941)
);

CKINVDCx20_ASAP7_75t_R g1942 ( 
.A(n_1789),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_SL g1943 ( 
.A1(n_1886),
.A2(n_801),
.B1(n_811),
.B2(n_806),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1774),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1793),
.B(n_1204),
.Y(n_1945)
);

INVx3_ASAP7_75t_L g1946 ( 
.A(n_1824),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1845),
.B(n_1205),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1780),
.B(n_1209),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1777),
.B(n_1210),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1781),
.Y(n_1950)
);

BUFx6f_ASAP7_75t_L g1951 ( 
.A(n_1840),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1837),
.B(n_1841),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_L g1953 ( 
.A(n_1820),
.B(n_1806),
.Y(n_1953)
);

INVx1_ASAP7_75t_L g1954 ( 
.A(n_1783),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1796),
.B(n_814),
.Y(n_1955)
);

INVx3_ASAP7_75t_L g1956 ( 
.A(n_1824),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1800),
.B(n_818),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_1834),
.Y(n_1958)
);

XOR2xp5_ASAP7_75t_L g1959 ( 
.A(n_1772),
.B(n_826),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1812),
.B(n_839),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1827),
.B(n_842),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1809),
.B(n_844),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1828),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1831),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1797),
.Y(n_1965)
);

NAND3xp33_ASAP7_75t_SL g1966 ( 
.A(n_1832),
.B(n_860),
.C(n_848),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1838),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1770),
.B(n_864),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1771),
.B(n_868),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1789),
.B(n_1008),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1902),
.B(n_1190),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1878),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1856),
.Y(n_1973)
);

INVx5_ASAP7_75t_L g1974 ( 
.A(n_1853),
.Y(n_1974)
);

BUFx3_ASAP7_75t_L g1975 ( 
.A(n_1860),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1834),
.Y(n_1976)
);

OR2x6_ASAP7_75t_L g1977 ( 
.A(n_1853),
.B(n_1044),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1833),
.B(n_872),
.Y(n_1978)
);

INVx1_ASAP7_75t_SL g1979 ( 
.A(n_1829),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1894),
.Y(n_1980)
);

INVx2_ASAP7_75t_SL g1981 ( 
.A(n_1868),
.Y(n_1981)
);

INVx3_ASAP7_75t_L g1982 ( 
.A(n_1914),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1900),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1830),
.B(n_873),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1790),
.A2(n_876),
.B1(n_877),
.B2(n_875),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1896),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1871),
.B(n_881),
.Y(n_1987)
);

INVx1_ASAP7_75t_SL g1988 ( 
.A(n_1829),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1904),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1880),
.Y(n_1990)
);

OR2x6_ASAP7_75t_L g1991 ( 
.A(n_1875),
.B(n_1046),
.Y(n_1991)
);

BUFx3_ASAP7_75t_L g1992 ( 
.A(n_1782),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1817),
.B(n_887),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_L g1994 ( 
.A(n_1869),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1775),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1785),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1768),
.A2(n_1003),
.B(n_963),
.Y(n_1997)
);

OAI21xp33_ASAP7_75t_L g1998 ( 
.A1(n_1821),
.A2(n_898),
.B(n_891),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1908),
.Y(n_1999)
);

INVx2_ASAP7_75t_SL g2000 ( 
.A(n_1842),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1823),
.B(n_901),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1909),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1835),
.B(n_1187),
.Y(n_2003)
);

BUFx6f_ASAP7_75t_L g2004 ( 
.A(n_1869),
.Y(n_2004)
);

BUFx3_ASAP7_75t_L g2005 ( 
.A(n_1846),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1901),
.Y(n_2006)
);

NAND2x1p5_ASAP7_75t_L g2007 ( 
.A(n_1810),
.B(n_1036),
.Y(n_2007)
);

BUFx8_ASAP7_75t_L g2008 ( 
.A(n_1903),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1892),
.B(n_1189),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1889),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1877),
.B(n_905),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1795),
.B(n_1050),
.Y(n_2012)
);

BUFx2_ASAP7_75t_L g2013 ( 
.A(n_1889),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1923),
.B(n_1883),
.Y(n_2014)
);

AND2x4_ASAP7_75t_L g2015 ( 
.A(n_1839),
.B(n_1051),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1825),
.B(n_914),
.Y(n_2016)
);

AOI22xp33_ASAP7_75t_L g2017 ( 
.A1(n_1819),
.A2(n_917),
.B1(n_921),
.B2(n_916),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1907),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_SL g2019 ( 
.A(n_1822),
.B(n_924),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1791),
.Y(n_2020)
);

AOI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1778),
.A2(n_926),
.B1(n_928),
.B2(n_925),
.Y(n_2021)
);

INVx5_ASAP7_75t_L g2022 ( 
.A(n_1787),
.Y(n_2022)
);

AOI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1855),
.A2(n_931),
.B1(n_932),
.B2(n_930),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1799),
.Y(n_2024)
);

OR2x6_ASAP7_75t_L g2025 ( 
.A(n_1867),
.B(n_1054),
.Y(n_2025)
);

HB1xp67_ASAP7_75t_L g2026 ( 
.A(n_1910),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1814),
.B(n_1815),
.Y(n_2027)
);

NOR2xp33_ASAP7_75t_L g2028 ( 
.A(n_1847),
.B(n_938),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1919),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1893),
.B(n_1192),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1849),
.B(n_940),
.Y(n_2031)
);

BUFx3_ASAP7_75t_L g2032 ( 
.A(n_1826),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1811),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1816),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1874),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1862),
.B(n_944),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_SL g2037 ( 
.A(n_1822),
.B(n_945),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_1863),
.B(n_947),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1852),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1921),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1912),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1895),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1805),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1872),
.B(n_951),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1807),
.Y(n_2045)
);

BUFx8_ASAP7_75t_SL g2046 ( 
.A(n_1916),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1922),
.B(n_952),
.Y(n_2047)
);

BUFx8_ASAP7_75t_L g2048 ( 
.A(n_1885),
.Y(n_2048)
);

BUFx3_ASAP7_75t_L g2049 ( 
.A(n_1934),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1917),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1867),
.Y(n_2051)
);

BUFx3_ASAP7_75t_L g2052 ( 
.A(n_1813),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1779),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1928),
.B(n_954),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1822),
.B(n_956),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1822),
.B(n_961),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1924),
.B(n_962),
.Y(n_2057)
);

INVx5_ASAP7_75t_L g2058 ( 
.A(n_1822),
.Y(n_2058)
);

OAI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1792),
.A2(n_1803),
.B(n_1843),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_SL g2060 ( 
.A(n_1851),
.B(n_964),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_1818),
.B(n_967),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1879),
.B(n_969),
.Y(n_2062)
);

INVx3_ASAP7_75t_L g2063 ( 
.A(n_1926),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_1915),
.B(n_1186),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1864),
.B(n_973),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1870),
.B(n_974),
.Y(n_2066)
);

BUFx2_ASAP7_75t_L g2067 ( 
.A(n_1881),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_1861),
.B(n_977),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_1926),
.Y(n_2069)
);

CKINVDCx5p33_ASAP7_75t_R g2070 ( 
.A(n_1858),
.Y(n_2070)
);

INVx2_ASAP7_75t_SL g2071 ( 
.A(n_1865),
.Y(n_2071)
);

OR2x6_ASAP7_75t_L g2072 ( 
.A(n_1911),
.B(n_1059),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1899),
.Y(n_2073)
);

INVx5_ASAP7_75t_L g2074 ( 
.A(n_1794),
.Y(n_2074)
);

CKINVDCx5p33_ASAP7_75t_R g2075 ( 
.A(n_1913),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1882),
.Y(n_2076)
);

OR2x6_ASAP7_75t_L g2077 ( 
.A(n_1891),
.B(n_1067),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1887),
.B(n_979),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1898),
.B(n_980),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1884),
.Y(n_2080)
);

BUFx6f_ASAP7_75t_L g2081 ( 
.A(n_1850),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_1920),
.Y(n_2082)
);

AND2x4_ASAP7_75t_L g2083 ( 
.A(n_1888),
.B(n_1088),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1890),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1944),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_2010),
.B(n_1769),
.Y(n_2086)
);

AND2x4_ASAP7_75t_L g2087 ( 
.A(n_2013),
.B(n_1784),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1950),
.Y(n_2088)
);

BUFx3_ASAP7_75t_L g2089 ( 
.A(n_1951),
.Y(n_2089)
);

INVx2_ASAP7_75t_L g2090 ( 
.A(n_2041),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1936),
.B(n_1899),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2026),
.B(n_1931),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1937),
.B(n_1897),
.Y(n_2093)
);

HB1xp67_ASAP7_75t_L g2094 ( 
.A(n_2018),
.Y(n_2094)
);

BUFx4f_ASAP7_75t_L g2095 ( 
.A(n_1938),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_2035),
.Y(n_2096)
);

BUFx3_ASAP7_75t_L g2097 ( 
.A(n_1951),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1954),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2036),
.B(n_981),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1967),
.B(n_1918),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2040),
.B(n_1798),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1972),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1953),
.B(n_1930),
.Y(n_2103)
);

HB1xp67_ASAP7_75t_L g2104 ( 
.A(n_1973),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1980),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_1994),
.Y(n_2106)
);

NOR2xp33_ASAP7_75t_L g2107 ( 
.A(n_1992),
.B(n_1929),
.Y(n_2107)
);

INVx4_ASAP7_75t_L g2108 ( 
.A(n_1938),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1986),
.Y(n_2109)
);

AND3x1_ASAP7_75t_SL g2110 ( 
.A(n_1963),
.B(n_1092),
.C(n_1090),
.Y(n_2110)
);

BUFx6f_ASAP7_75t_L g2111 ( 
.A(n_1994),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2062),
.B(n_1932),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1952),
.B(n_1804),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_SL g2114 ( 
.A(n_1943),
.B(n_1859),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_1983),
.B(n_1844),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_SL g2116 ( 
.A(n_1958),
.B(n_1927),
.Y(n_2116)
);

INVx4_ASAP7_75t_L g2117 ( 
.A(n_1946),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2013),
.B(n_982),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1964),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_2043),
.B(n_1905),
.Y(n_2120)
);

CKINVDCx20_ASAP7_75t_R g2121 ( 
.A(n_1942),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_1956),
.Y(n_2122)
);

INVx4_ASAP7_75t_L g2123 ( 
.A(n_1990),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_2005),
.B(n_983),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1989),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1993),
.B(n_984),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_2059),
.A2(n_1801),
.B(n_1848),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1995),
.Y(n_2128)
);

BUFx6f_ASAP7_75t_L g2129 ( 
.A(n_2004),
.Y(n_2129)
);

AND2x2_ASAP7_75t_L g2130 ( 
.A(n_2014),
.B(n_986),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1996),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_2039),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_1990),
.Y(n_2133)
);

BUFx12f_ASAP7_75t_L g2134 ( 
.A(n_1970),
.Y(n_2134)
);

INVx2_ASAP7_75t_SL g2135 ( 
.A(n_1974),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_2004),
.B(n_2032),
.Y(n_2136)
);

NOR2xp33_ASAP7_75t_L g2137 ( 
.A(n_1966),
.B(n_1906),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1965),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2020),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1999),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_2002),
.Y(n_2141)
);

INVx4_ASAP7_75t_L g2142 ( 
.A(n_1976),
.Y(n_2142)
);

HB1xp67_ASAP7_75t_L g2143 ( 
.A(n_1973),
.Y(n_2143)
);

HB1xp67_ASAP7_75t_L g2144 ( 
.A(n_1991),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2053),
.B(n_989),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2082),
.B(n_992),
.Y(n_2146)
);

INVxp67_ASAP7_75t_L g2147 ( 
.A(n_1962),
.Y(n_2147)
);

AO22x1_ASAP7_75t_L g2148 ( 
.A1(n_2074),
.A2(n_1122),
.B1(n_1123),
.B2(n_1118),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2024),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_2081),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2016),
.A2(n_1802),
.B1(n_1788),
.B2(n_1873),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_SL g2152 ( 
.A(n_2074),
.B(n_1808),
.Y(n_2152)
);

NOR2xp33_ASAP7_75t_L g2153 ( 
.A(n_2068),
.B(n_1854),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1948),
.B(n_996),
.Y(n_2154)
);

BUFx2_ASAP7_75t_L g2155 ( 
.A(n_2046),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1945),
.B(n_997),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2028),
.B(n_2045),
.Y(n_2157)
);

BUFx2_ASAP7_75t_SL g2158 ( 
.A(n_1974),
.Y(n_2158)
);

NAND2xp5_ASAP7_75t_L g2159 ( 
.A(n_1991),
.B(n_999),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2061),
.B(n_1004),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_2009),
.B(n_1011),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2030),
.B(n_1012),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2033),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2073),
.B(n_1013),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2017),
.B(n_1015),
.Y(n_2165)
);

AOI22xp33_ASAP7_75t_L g2166 ( 
.A1(n_1998),
.A2(n_1802),
.B1(n_1933),
.B2(n_1786),
.Y(n_2166)
);

CKINVDCx6p67_ASAP7_75t_R g2167 ( 
.A(n_1974),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2034),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2029),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1947),
.B(n_1016),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_2050),
.B(n_1020),
.Y(n_2171)
);

NOR2xp67_ASAP7_75t_L g2172 ( 
.A(n_1981),
.B(n_516),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2006),
.Y(n_2173)
);

AND2x4_ASAP7_75t_L g2174 ( 
.A(n_1975),
.B(n_2051),
.Y(n_2174)
);

CKINVDCx16_ASAP7_75t_R g2175 ( 
.A(n_1940),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_2081),
.Y(n_2176)
);

OR2x6_ASAP7_75t_L g2177 ( 
.A(n_1977),
.B(n_1925),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_2052),
.Y(n_2178)
);

AOI22xp5_ASAP7_75t_L g2179 ( 
.A1(n_1979),
.A2(n_1022),
.B1(n_1026),
.B2(n_1023),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2084),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_1988),
.A2(n_1031),
.B1(n_1041),
.B2(n_1034),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2049),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2027),
.B(n_1045),
.Y(n_2183)
);

AND2x2_ASAP7_75t_L g2184 ( 
.A(n_2063),
.B(n_2069),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2067),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_2042),
.B(n_1049),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2042),
.B(n_1055),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2067),
.Y(n_2188)
);

CKINVDCx5p33_ASAP7_75t_R g2189 ( 
.A(n_2008),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1941),
.B(n_1056),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_2057),
.B(n_1058),
.Y(n_2191)
);

INVx2_ASAP7_75t_L g2192 ( 
.A(n_2076),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2080),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_2074),
.B(n_1212),
.Y(n_2194)
);

INVx3_ASAP7_75t_L g2195 ( 
.A(n_2058),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1955),
.Y(n_2196)
);

INVx2_ASAP7_75t_L g2197 ( 
.A(n_1982),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1957),
.Y(n_2198)
);

NAND2xp5_ASAP7_75t_L g2199 ( 
.A(n_1968),
.B(n_1969),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2001),
.B(n_1060),
.Y(n_2200)
);

BUFx12f_ASAP7_75t_L g2201 ( 
.A(n_1977),
.Y(n_2201)
);

AOI21xp5_ASAP7_75t_L g2202 ( 
.A1(n_1997),
.A2(n_1048),
.B(n_1021),
.Y(n_2202)
);

INVxp67_ASAP7_75t_SL g2203 ( 
.A(n_2066),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1960),
.Y(n_2204)
);

BUFx2_ASAP7_75t_L g2205 ( 
.A(n_2070),
.Y(n_2205)
);

NAND3xp33_ASAP7_75t_L g2206 ( 
.A(n_2065),
.B(n_1062),
.C(n_1061),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_2003),
.B(n_1063),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_SL g2208 ( 
.A(n_2000),
.B(n_2075),
.Y(n_2208)
);

AND2x2_ASAP7_75t_L g2209 ( 
.A(n_1985),
.B(n_1064),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1949),
.B(n_1065),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2011),
.B(n_1069),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_2048),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_2058),
.Y(n_2213)
);

AOI22xp33_ASAP7_75t_L g2214 ( 
.A1(n_2025),
.A2(n_1130),
.B1(n_1155),
.B2(n_1036),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1961),
.Y(n_2215)
);

BUFx3_ASAP7_75t_L g2216 ( 
.A(n_2071),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_SL g2217 ( 
.A(n_2058),
.B(n_1197),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2012),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1971),
.Y(n_2219)
);

CKINVDCx5p33_ASAP7_75t_R g2220 ( 
.A(n_2022),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2044),
.Y(n_2221)
);

NOR2xp33_ASAP7_75t_L g2222 ( 
.A(n_1984),
.B(n_1072),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_2023),
.B(n_1073),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2021),
.B(n_1074),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_2031),
.B(n_1075),
.Y(n_2225)
);

INVx2_ASAP7_75t_L g2226 ( 
.A(n_1939),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2038),
.B(n_1076),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_2064),
.B(n_1077),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_SL g2229 ( 
.A(n_2079),
.B(n_1052),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2077),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_SL g2231 ( 
.A1(n_1959),
.A2(n_1079),
.B1(n_1084),
.B2(n_1083),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2077),
.Y(n_2232)
);

AOI22x1_ASAP7_75t_L g2233 ( 
.A1(n_2007),
.A2(n_1087),
.B1(n_1093),
.B2(n_1085),
.Y(n_2233)
);

OAI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_1978),
.A2(n_1095),
.B1(n_1097),
.B2(n_1094),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2015),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2060),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1987),
.Y(n_2237)
);

BUFx6f_ASAP7_75t_L g2238 ( 
.A(n_2025),
.Y(n_2238)
);

CKINVDCx5p33_ASAP7_75t_R g2239 ( 
.A(n_2121),
.Y(n_2239)
);

NAND2x1_ASAP7_75t_L g2240 ( 
.A(n_2195),
.B(n_2072),
.Y(n_2240)
);

BUFx6f_ASAP7_75t_L g2241 ( 
.A(n_2089),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_2127),
.A2(n_2037),
.B(n_2019),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2125),
.Y(n_2243)
);

OAI21xp5_ASAP7_75t_L g2244 ( 
.A1(n_2126),
.A2(n_2222),
.B(n_2147),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_2102),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2157),
.B(n_2083),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2103),
.A2(n_2072),
.B1(n_2078),
.B2(n_2054),
.Y(n_2247)
);

OAI21x1_ASAP7_75t_L g2248 ( 
.A1(n_2226),
.A2(n_2056),
.B(n_2055),
.Y(n_2248)
);

INVx6_ASAP7_75t_L g2249 ( 
.A(n_2134),
.Y(n_2249)
);

NOR2x1_ASAP7_75t_SL g2250 ( 
.A(n_2177),
.B(n_2022),
.Y(n_2250)
);

OAI21x1_ASAP7_75t_L g2251 ( 
.A1(n_2195),
.A2(n_1096),
.B(n_1053),
.Y(n_2251)
);

AOI211x1_ASAP7_75t_L g2252 ( 
.A1(n_2209),
.A2(n_1214),
.B(n_1208),
.C(n_1132),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_2153),
.B(n_2022),
.Y(n_2253)
);

OAI21xp5_ASAP7_75t_L g2254 ( 
.A1(n_2199),
.A2(n_2047),
.B(n_1133),
.Y(n_2254)
);

OAI21x1_ASAP7_75t_L g2255 ( 
.A1(n_2166),
.A2(n_1184),
.B(n_1173),
.Y(n_2255)
);

OAI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2112),
.A2(n_1959),
.B1(n_1136),
.B2(n_1143),
.Y(n_2256)
);

AOI21xp5_ASAP7_75t_L g2257 ( 
.A1(n_2113),
.A2(n_1108),
.B(n_1107),
.Y(n_2257)
);

OAI21x1_ASAP7_75t_L g2258 ( 
.A1(n_2151),
.A2(n_1146),
.B(n_1135),
.Y(n_2258)
);

BUFx6f_ASAP7_75t_L g2259 ( 
.A(n_2097),
.Y(n_2259)
);

AOI21xp5_ASAP7_75t_L g2260 ( 
.A1(n_2120),
.A2(n_1174),
.B(n_1165),
.Y(n_2260)
);

AO31x2_ASAP7_75t_L g2261 ( 
.A1(n_2192),
.A2(n_1203),
.A3(n_1201),
.B(n_1145),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2094),
.B(n_1131),
.Y(n_2262)
);

AO21x1_ASAP7_75t_L g2263 ( 
.A1(n_2202),
.A2(n_1153),
.B(n_1150),
.Y(n_2263)
);

AOI21xp5_ASAP7_75t_L g2264 ( 
.A1(n_2152),
.A2(n_1182),
.B(n_1162),
.Y(n_2264)
);

OAI21x1_ASAP7_75t_L g2265 ( 
.A1(n_2173),
.A2(n_2088),
.B(n_2085),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2098),
.A2(n_1177),
.B(n_1154),
.Y(n_2266)
);

OAI22x1_ASAP7_75t_L g2267 ( 
.A1(n_2091),
.A2(n_1185),
.B1(n_1193),
.B2(n_1178),
.Y(n_2267)
);

OAI21x1_ASAP7_75t_L g2268 ( 
.A1(n_2119),
.A2(n_1198),
.B(n_1196),
.Y(n_2268)
);

AOI21x1_ASAP7_75t_L g2269 ( 
.A1(n_2148),
.A2(n_1155),
.B(n_1130),
.Y(n_2269)
);

BUFx12f_ASAP7_75t_L g2270 ( 
.A(n_2189),
.Y(n_2270)
);

BUFx4f_ASAP7_75t_SL g2271 ( 
.A(n_2201),
.Y(n_2271)
);

BUFx4_ASAP7_75t_SL g2272 ( 
.A(n_2212),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2115),
.A2(n_816),
.B(n_748),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2118),
.B(n_1099),
.Y(n_2274)
);

AOI21x1_ASAP7_75t_L g2275 ( 
.A1(n_2148),
.A2(n_789),
.B(n_815),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_2133),
.Y(n_2276)
);

OAI21x1_ASAP7_75t_L g2277 ( 
.A1(n_2140),
.A2(n_789),
.B(n_518),
.Y(n_2277)
);

OAI21xp5_ASAP7_75t_L g2278 ( 
.A1(n_2161),
.A2(n_1113),
.B(n_1101),
.Y(n_2278)
);

NOR2x1_ASAP7_75t_SL g2279 ( 
.A(n_2177),
.B(n_815),
.Y(n_2279)
);

OAI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2141),
.A2(n_789),
.B(n_519),
.Y(n_2280)
);

AOI21x1_ASAP7_75t_L g2281 ( 
.A1(n_2217),
.A2(n_789),
.B(n_815),
.Y(n_2281)
);

NOR2xp67_ASAP7_75t_SL g2282 ( 
.A(n_2175),
.B(n_815),
.Y(n_2282)
);

OAI21xp5_ASAP7_75t_L g2283 ( 
.A1(n_2162),
.A2(n_1172),
.B(n_1156),
.Y(n_2283)
);

NAND2x1p5_ASAP7_75t_L g2284 ( 
.A(n_2095),
.B(n_1152),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_L g2285 ( 
.A1(n_2203),
.A2(n_919),
.B(n_850),
.Y(n_2285)
);

OAI22x1_ASAP7_75t_L g2286 ( 
.A1(n_2232),
.A2(n_1103),
.B1(n_1104),
.B2(n_1102),
.Y(n_2286)
);

OAI21xp5_ASAP7_75t_L g2287 ( 
.A1(n_2191),
.A2(n_1141),
.B(n_1110),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_SL g2288 ( 
.A(n_2093),
.B(n_704),
.Y(n_2288)
);

OAI21xp5_ASAP7_75t_L g2289 ( 
.A1(n_2156),
.A2(n_2206),
.B(n_2190),
.Y(n_2289)
);

AOI21xp5_ASAP7_75t_L g2290 ( 
.A1(n_2213),
.A2(n_919),
.B(n_850),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2149),
.Y(n_2291)
);

NAND3xp33_ASAP7_75t_L g2292 ( 
.A(n_2114),
.B(n_1109),
.C(n_1106),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2213),
.A2(n_2221),
.B(n_2194),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2196),
.B(n_1111),
.Y(n_2294)
);

OAI21x1_ASAP7_75t_L g2295 ( 
.A1(n_2193),
.A2(n_789),
.B(n_520),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2198),
.B(n_1114),
.Y(n_2296)
);

INVx2_ASAP7_75t_L g2297 ( 
.A(n_2105),
.Y(n_2297)
);

INVx2_ASAP7_75t_SL g2298 ( 
.A(n_2136),
.Y(n_2298)
);

AOI21x1_ASAP7_75t_L g2299 ( 
.A1(n_2180),
.A2(n_789),
.B(n_850),
.Y(n_2299)
);

BUFx4f_ASAP7_75t_L g2300 ( 
.A(n_2167),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2163),
.Y(n_2301)
);

OAI21x1_ASAP7_75t_L g2302 ( 
.A1(n_2168),
.A2(n_789),
.B(n_523),
.Y(n_2302)
);

BUFx6f_ASAP7_75t_L g2303 ( 
.A(n_2106),
.Y(n_2303)
);

OAI21xp5_ASAP7_75t_L g2304 ( 
.A1(n_2200),
.A2(n_2207),
.B(n_2210),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2205),
.B(n_1115),
.Y(n_2305)
);

OAI21xp5_ASAP7_75t_L g2306 ( 
.A1(n_2170),
.A2(n_1175),
.B(n_1151),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_2204),
.B(n_1116),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2213),
.A2(n_919),
.B(n_850),
.Y(n_2308)
);

AOI21xp5_ASAP7_75t_SL g2309 ( 
.A1(n_2219),
.A2(n_990),
.B(n_919),
.Y(n_2309)
);

OAI22xp5_ASAP7_75t_L g2310 ( 
.A1(n_2137),
.A2(n_1119),
.B1(n_1120),
.B2(n_1117),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_2215),
.B(n_2150),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2139),
.Y(n_2312)
);

AO32x2_ASAP7_75t_L g2313 ( 
.A1(n_2234),
.A2(n_1125),
.A3(n_1148),
.B1(n_1137),
.B2(n_1128),
.Y(n_2313)
);

AO31x2_ASAP7_75t_L g2314 ( 
.A1(n_2128),
.A2(n_524),
.A3(n_525),
.B(n_517),
.Y(n_2314)
);

OAI21xp5_ASAP7_75t_L g2315 ( 
.A1(n_2154),
.A2(n_1169),
.B(n_1161),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2229),
.A2(n_1078),
.B(n_990),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2101),
.B(n_1160),
.Y(n_2317)
);

OAI21x1_ASAP7_75t_L g2318 ( 
.A1(n_2185),
.A2(n_528),
.B(n_526),
.Y(n_2318)
);

OAI21x1_ASAP7_75t_L g2319 ( 
.A1(n_2188),
.A2(n_533),
.B(n_532),
.Y(n_2319)
);

BUFx2_ASAP7_75t_L g2320 ( 
.A(n_2174),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2109),
.Y(n_2321)
);

AND2x6_ASAP7_75t_SL g2322 ( 
.A(n_2186),
.B(n_1164),
.Y(n_2322)
);

NOR2x1_ASAP7_75t_R g2323 ( 
.A(n_2108),
.B(n_1180),
.Y(n_2323)
);

OAI21xp5_ASAP7_75t_L g2324 ( 
.A1(n_2228),
.A2(n_2227),
.B(n_2225),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_L g2325 ( 
.A1(n_2224),
.A2(n_1181),
.B(n_713),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2090),
.Y(n_2326)
);

NAND3xp33_ASAP7_75t_L g2327 ( 
.A(n_2223),
.B(n_1078),
.C(n_990),
.Y(n_2327)
);

NAND3x1_ASAP7_75t_L g2328 ( 
.A(n_2107),
.B(n_0),
.C(n_1),
.Y(n_2328)
);

OAI21x1_ASAP7_75t_L g2329 ( 
.A1(n_2182),
.A2(n_536),
.B(n_535),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2092),
.B(n_990),
.Y(n_2330)
);

AO32x2_ASAP7_75t_L g2331 ( 
.A1(n_2135),
.A2(n_1171),
.A3(n_1144),
.B1(n_1078),
.B2(n_4),
.Y(n_2331)
);

INVx3_ASAP7_75t_L g2332 ( 
.A(n_2123),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2160),
.B(n_1078),
.Y(n_2333)
);

OA22x2_ASAP7_75t_L g2334 ( 
.A1(n_2230),
.A2(n_725),
.B1(n_728),
.B2(n_710),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2104),
.B(n_1144),
.Y(n_2335)
);

NAND3xp33_ASAP7_75t_L g2336 ( 
.A(n_2165),
.B(n_2233),
.C(n_2237),
.Y(n_2336)
);

OAI21x1_ASAP7_75t_L g2337 ( 
.A1(n_2236),
.A2(n_545),
.B(n_543),
.Y(n_2337)
);

AOI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2145),
.A2(n_1171),
.B(n_1144),
.Y(n_2338)
);

AO31x2_ASAP7_75t_L g2339 ( 
.A1(n_2131),
.A2(n_547),
.A3(n_550),
.B(n_546),
.Y(n_2339)
);

O2A1O1Ixp5_ASAP7_75t_L g2340 ( 
.A1(n_2208),
.A2(n_1171),
.B(n_1144),
.C(n_4),
.Y(n_2340)
);

AOI21xp5_ASAP7_75t_L g2341 ( 
.A1(n_2087),
.A2(n_1171),
.B(n_732),
.Y(n_2341)
);

AOI21xp5_ASAP7_75t_L g2342 ( 
.A1(n_2087),
.A2(n_2143),
.B(n_2171),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_2096),
.B(n_2),
.Y(n_2343)
);

AND2x2_ASAP7_75t_L g2344 ( 
.A(n_2099),
.B(n_2),
.Y(n_2344)
);

NOR2xp67_ASAP7_75t_SL g2345 ( 
.A(n_2158),
.B(n_1213),
.Y(n_2345)
);

AOI21xp5_ASAP7_75t_L g2346 ( 
.A1(n_2086),
.A2(n_737),
.B(n_715),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2164),
.B(n_3),
.Y(n_2347)
);

OAI21x1_ASAP7_75t_L g2348 ( 
.A1(n_2132),
.A2(n_559),
.B(n_552),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2169),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2144),
.B(n_6),
.Y(n_2350)
);

O2A1O1Ixp33_ASAP7_75t_L g2351 ( 
.A1(n_2211),
.A2(n_8),
.B(n_6),
.C(n_7),
.Y(n_2351)
);

OAI21x1_ASAP7_75t_L g2352 ( 
.A1(n_2184),
.A2(n_562),
.B(n_560),
.Y(n_2352)
);

CKINVDCx5p33_ASAP7_75t_R g2353 ( 
.A(n_2220),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2178),
.Y(n_2354)
);

NAND2xp33_ASAP7_75t_L g2355 ( 
.A(n_2150),
.B(n_2176),
.Y(n_2355)
);

INVxp67_ASAP7_75t_SL g2356 ( 
.A(n_2100),
.Y(n_2356)
);

OA22x2_ASAP7_75t_L g2357 ( 
.A1(n_2218),
.A2(n_742),
.B1(n_756),
.B2(n_740),
.Y(n_2357)
);

OAI21xp5_ASAP7_75t_L g2358 ( 
.A1(n_2159),
.A2(n_774),
.B(n_757),
.Y(n_2358)
);

AOI22x1_ASAP7_75t_L g2359 ( 
.A1(n_2117),
.A2(n_859),
.B1(n_895),
.B2(n_820),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2138),
.B(n_8),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2136),
.B(n_9),
.Y(n_2361)
);

OAI21xp5_ASAP7_75t_L g2362 ( 
.A1(n_2124),
.A2(n_786),
.B(n_778),
.Y(n_2362)
);

OAI21x1_ASAP7_75t_L g2363 ( 
.A1(n_2172),
.A2(n_565),
.B(n_563),
.Y(n_2363)
);

O2A1O1Ixp5_ASAP7_75t_L g2364 ( 
.A1(n_2142),
.A2(n_2086),
.B(n_2146),
.C(n_2197),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2150),
.Y(n_2365)
);

NOR4xp25_ASAP7_75t_L g2366 ( 
.A(n_2214),
.B(n_13),
.C(n_11),
.D(n_12),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2176),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_2238),
.B(n_2216),
.Y(n_2368)
);

OAI21xp5_ASAP7_75t_L g2369 ( 
.A1(n_2179),
.A2(n_791),
.B(n_780),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_2238),
.B(n_12),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2238),
.B(n_14),
.Y(n_2371)
);

AOI22xp33_ASAP7_75t_L g2372 ( 
.A1(n_2235),
.A2(n_802),
.B1(n_804),
.B2(n_793),
.Y(n_2372)
);

OAI21x1_ASAP7_75t_L g2373 ( 
.A1(n_2183),
.A2(n_567),
.B(n_566),
.Y(n_2373)
);

INVxp67_ASAP7_75t_SL g2374 ( 
.A(n_2106),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2176),
.Y(n_2375)
);

A2O1A1Ixp33_ASAP7_75t_L g2376 ( 
.A1(n_2231),
.A2(n_822),
.B(n_823),
.C(n_821),
.Y(n_2376)
);

OAI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2181),
.A2(n_829),
.B1(n_851),
.B2(n_840),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2130),
.B(n_2174),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2117),
.A2(n_865),
.B(n_827),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2123),
.B(n_2116),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_SL g2381 ( 
.A(n_2106),
.B(n_869),
.Y(n_2381)
);

OR2x2_ASAP7_75t_L g2382 ( 
.A(n_2111),
.B(n_14),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2291),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2245),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2301),
.Y(n_2385)
);

OAI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2244),
.A2(n_2187),
.B(n_2142),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2320),
.B(n_2108),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_L g2388 ( 
.A(n_2356),
.B(n_2111),
.Y(n_2388)
);

OR2x6_ASAP7_75t_L g2389 ( 
.A(n_2240),
.B(n_2380),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_2297),
.Y(n_2390)
);

AOI22xp33_ASAP7_75t_L g2391 ( 
.A1(n_2256),
.A2(n_2111),
.B1(n_2129),
.B2(n_2155),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2349),
.B(n_2129),
.Y(n_2392)
);

CKINVDCx5p33_ASAP7_75t_R g2393 ( 
.A(n_2272),
.Y(n_2393)
);

INVxp67_ASAP7_75t_SL g2394 ( 
.A(n_2265),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2241),
.Y(n_2395)
);

CKINVDCx20_ASAP7_75t_R g2396 ( 
.A(n_2239),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2335),
.Y(n_2397)
);

AOI21xp5_ASAP7_75t_L g2398 ( 
.A1(n_2242),
.A2(n_2129),
.B(n_2122),
.Y(n_2398)
);

INVx2_ASAP7_75t_SL g2399 ( 
.A(n_2241),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_2253),
.B(n_15),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2243),
.Y(n_2401)
);

CKINVDCx8_ASAP7_75t_R g2402 ( 
.A(n_2322),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2312),
.Y(n_2403)
);

OAI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2292),
.A2(n_2110),
.B1(n_933),
.B2(n_966),
.Y(n_2404)
);

AOI21xp33_ASAP7_75t_L g2405 ( 
.A1(n_2351),
.A2(n_935),
.B(n_886),
.Y(n_2405)
);

INVx5_ASAP7_75t_L g2406 ( 
.A(n_2303),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2321),
.Y(n_2407)
);

INVx3_ASAP7_75t_L g2408 ( 
.A(n_2259),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2326),
.Y(n_2409)
);

AND2x4_ASAP7_75t_L g2410 ( 
.A(n_2298),
.B(n_568),
.Y(n_2410)
);

AOI21xp5_ASAP7_75t_L g2411 ( 
.A1(n_2285),
.A2(n_883),
.B(n_871),
.Y(n_2411)
);

AOI21xp5_ASAP7_75t_L g2412 ( 
.A1(n_2338),
.A2(n_892),
.B(n_888),
.Y(n_2412)
);

OA21x2_ASAP7_75t_L g2413 ( 
.A1(n_2248),
.A2(n_908),
.B(n_899),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2354),
.Y(n_2414)
);

INVx4_ASAP7_75t_SL g2415 ( 
.A(n_2271),
.Y(n_2415)
);

BUFx2_ASAP7_75t_L g2416 ( 
.A(n_2374),
.Y(n_2416)
);

O2A1O1Ixp5_ASAP7_75t_SL g2417 ( 
.A1(n_2311),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2261),
.Y(n_2418)
);

AND2x4_ASAP7_75t_L g2419 ( 
.A(n_2276),
.B(n_576),
.Y(n_2419)
);

INVx4_ASAP7_75t_L g2420 ( 
.A(n_2300),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2342),
.B(n_18),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_2364),
.B(n_918),
.Y(n_2422)
);

AND2x2_ASAP7_75t_L g2423 ( 
.A(n_2347),
.B(n_20),
.Y(n_2423)
);

INVx4_ASAP7_75t_L g2424 ( 
.A(n_2353),
.Y(n_2424)
);

AND2x2_ASAP7_75t_L g2425 ( 
.A(n_2378),
.B(n_20),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2365),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_2293),
.B(n_922),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2250),
.B(n_577),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2246),
.B(n_2330),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2261),
.Y(n_2430)
);

INVx2_ASAP7_75t_L g2431 ( 
.A(n_2367),
.Y(n_2431)
);

AND2x4_ASAP7_75t_L g2432 ( 
.A(n_2375),
.B(n_579),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2343),
.B(n_21),
.Y(n_2433)
);

INVx5_ASAP7_75t_L g2434 ( 
.A(n_2303),
.Y(n_2434)
);

CKINVDCx5p33_ASAP7_75t_R g2435 ( 
.A(n_2270),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2261),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_2259),
.Y(n_2437)
);

CKINVDCx20_ASAP7_75t_R g2438 ( 
.A(n_2249),
.Y(n_2438)
);

OAI22xp5_ASAP7_75t_L g2439 ( 
.A1(n_2247),
.A2(n_1001),
.B1(n_1124),
.B2(n_941),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2344),
.B(n_21),
.Y(n_2440)
);

NOR2x1_ASAP7_75t_SL g2441 ( 
.A(n_2368),
.B(n_23),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2331),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2328),
.A2(n_1029),
.B1(n_1080),
.B2(n_955),
.Y(n_2443)
);

BUFx8_ASAP7_75t_L g2444 ( 
.A(n_2274),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2262),
.B(n_23),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2331),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_2304),
.B(n_2324),
.Y(n_2447)
);

INVx1_ASAP7_75t_SL g2448 ( 
.A(n_2249),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2331),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2333),
.B(n_24),
.Y(n_2450)
);

AND2x4_ASAP7_75t_L g2451 ( 
.A(n_2332),
.B(n_583),
.Y(n_2451)
);

INVx2_ASAP7_75t_L g2452 ( 
.A(n_2299),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_SL g2453 ( 
.A(n_2254),
.B(n_927),
.Y(n_2453)
);

OAI21x1_ASAP7_75t_SL g2454 ( 
.A1(n_2279),
.A2(n_26),
.B(n_25),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2309),
.A2(n_946),
.B(n_936),
.Y(n_2455)
);

BUFx12f_ASAP7_75t_L g2456 ( 
.A(n_2284),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2361),
.B(n_24),
.Y(n_2457)
);

INVx2_ASAP7_75t_SL g2458 ( 
.A(n_2382),
.Y(n_2458)
);

AOI21xp5_ASAP7_75t_L g2459 ( 
.A1(n_2257),
.A2(n_2260),
.B(n_2289),
.Y(n_2459)
);

NOR2xp67_ASAP7_75t_L g2460 ( 
.A(n_2336),
.B(n_26),
.Y(n_2460)
);

AOI22xp33_ASAP7_75t_L g2461 ( 
.A1(n_2267),
.A2(n_965),
.B1(n_971),
.B2(n_959),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2266),
.Y(n_2462)
);

A2O1A1Ixp33_ASAP7_75t_L g2463 ( 
.A1(n_2273),
.A2(n_995),
.B(n_1025),
.C(n_985),
.Y(n_2463)
);

BUFx6f_ASAP7_75t_L g2464 ( 
.A(n_2370),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_2360),
.B(n_27),
.Y(n_2465)
);

INVx1_ASAP7_75t_SL g2466 ( 
.A(n_2355),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_SL g2467 ( 
.A(n_2366),
.B(n_1027),
.Y(n_2467)
);

INVxp67_ASAP7_75t_SL g2468 ( 
.A(n_2263),
.Y(n_2468)
);

INVx3_ASAP7_75t_L g2469 ( 
.A(n_2334),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2314),
.Y(n_2470)
);

AND2x4_ASAP7_75t_L g2471 ( 
.A(n_2371),
.B(n_2350),
.Y(n_2471)
);

AND2x4_ASAP7_75t_L g2472 ( 
.A(n_2268),
.B(n_2352),
.Y(n_2472)
);

O2A1O1Ixp33_ASAP7_75t_L g2473 ( 
.A1(n_2310),
.A2(n_31),
.B(n_28),
.C(n_29),
.Y(n_2473)
);

INVx5_ASAP7_75t_L g2474 ( 
.A(n_2282),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2317),
.B(n_2252),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2305),
.B(n_29),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2314),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2357),
.B(n_31),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2381),
.Y(n_2479)
);

NOR2xp33_ASAP7_75t_L g2480 ( 
.A(n_2323),
.B(n_32),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2314),
.Y(n_2481)
);

OR2x2_ASAP7_75t_SL g2482 ( 
.A(n_2294),
.B(n_33),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2296),
.B(n_34),
.Y(n_2483)
);

AND2x4_ASAP7_75t_L g2484 ( 
.A(n_2251),
.B(n_585),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_2288),
.A2(n_1098),
.B(n_1081),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2339),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2339),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_2363),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2307),
.B(n_35),
.Y(n_2489)
);

NOR2xp67_ASAP7_75t_R g2490 ( 
.A(n_2474),
.B(n_2345),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2403),
.Y(n_2491)
);

AND2x2_ASAP7_75t_L g2492 ( 
.A(n_2416),
.B(n_2383),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_2447),
.B(n_2286),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2397),
.B(n_35),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_2385),
.B(n_2258),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2401),
.Y(n_2496)
);

CKINVDCx5p33_ASAP7_75t_R g2497 ( 
.A(n_2393),
.Y(n_2497)
);

BUFx6f_ASAP7_75t_L g2498 ( 
.A(n_2406),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_2407),
.Y(n_2499)
);

OR2x2_ASAP7_75t_L g2500 ( 
.A(n_2416),
.B(n_2327),
.Y(n_2500)
);

INVxp67_ASAP7_75t_SL g2501 ( 
.A(n_2394),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_2409),
.Y(n_2502)
);

AND2x4_ASAP7_75t_L g2503 ( 
.A(n_2389),
.B(n_2339),
.Y(n_2503)
);

AOI21xp5_ASAP7_75t_L g2504 ( 
.A1(n_2459),
.A2(n_2308),
.B(n_2290),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_2448),
.B(n_2376),
.Y(n_2505)
);

NOR2xp67_ASAP7_75t_L g2506 ( 
.A(n_2398),
.B(n_2275),
.Y(n_2506)
);

AOI21xp5_ASAP7_75t_L g2507 ( 
.A1(n_2422),
.A2(n_2340),
.B(n_2341),
.Y(n_2507)
);

NAND2xp5_ASAP7_75t_SL g2508 ( 
.A(n_2466),
.B(n_2358),
.Y(n_2508)
);

O2A1O1Ixp5_ASAP7_75t_L g2509 ( 
.A1(n_2467),
.A2(n_2325),
.B(n_2264),
.C(n_2283),
.Y(n_2509)
);

HB1xp67_ASAP7_75t_L g2510 ( 
.A(n_2392),
.Y(n_2510)
);

AOI21xp5_ASAP7_75t_L g2511 ( 
.A1(n_2427),
.A2(n_2280),
.B(n_2277),
.Y(n_2511)
);

A2O1A1Ixp33_ASAP7_75t_L g2512 ( 
.A1(n_2460),
.A2(n_2278),
.B(n_2287),
.C(n_2315),
.Y(n_2512)
);

AOI21xp33_ASAP7_75t_L g2513 ( 
.A1(n_2439),
.A2(n_2373),
.B(n_2329),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2431),
.Y(n_2514)
);

AND2x2_ASAP7_75t_L g2515 ( 
.A(n_2425),
.B(n_2313),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_2429),
.B(n_36),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2458),
.B(n_2255),
.Y(n_2517)
);

AND2x2_ASAP7_75t_L g2518 ( 
.A(n_2471),
.B(n_2313),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2414),
.Y(n_2519)
);

AND2x4_ASAP7_75t_L g2520 ( 
.A(n_2389),
.B(n_2295),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2426),
.Y(n_2521)
);

HB1xp67_ASAP7_75t_L g2522 ( 
.A(n_2388),
.Y(n_2522)
);

OA21x2_ASAP7_75t_L g2523 ( 
.A1(n_2477),
.A2(n_2302),
.B(n_2318),
.Y(n_2523)
);

AND2x2_ASAP7_75t_L g2524 ( 
.A(n_2387),
.B(n_2313),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_2444),
.B(n_37),
.Y(n_2525)
);

O2A1O1Ixp33_ASAP7_75t_L g2526 ( 
.A1(n_2453),
.A2(n_2306),
.B(n_2369),
.C(n_2377),
.Y(n_2526)
);

OA21x2_ASAP7_75t_L g2527 ( 
.A1(n_2481),
.A2(n_2319),
.B(n_2337),
.Y(n_2527)
);

OR2x6_ASAP7_75t_SL g2528 ( 
.A(n_2435),
.B(n_1121),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2384),
.Y(n_2529)
);

OR2x2_ASAP7_75t_L g2530 ( 
.A(n_2449),
.B(n_37),
.Y(n_2530)
);

AOI21xp5_ASAP7_75t_SL g2531 ( 
.A1(n_2421),
.A2(n_2428),
.B(n_2441),
.Y(n_2531)
);

A2O1A1Ixp33_ASAP7_75t_SL g2532 ( 
.A1(n_2400),
.A2(n_2473),
.B(n_2480),
.C(n_2476),
.Y(n_2532)
);

NAND2xp5_ASAP7_75t_L g2533 ( 
.A(n_2442),
.B(n_38),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_2423),
.B(n_38),
.Y(n_2534)
);

BUFx4_ASAP7_75t_R g2535 ( 
.A(n_2395),
.Y(n_2535)
);

INVx1_ASAP7_75t_L g2536 ( 
.A(n_2390),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2386),
.B(n_39),
.Y(n_2537)
);

NAND2x1p5_ASAP7_75t_L g2538 ( 
.A(n_2474),
.B(n_2269),
.Y(n_2538)
);

AOI21xp5_ASAP7_75t_L g2539 ( 
.A1(n_2472),
.A2(n_2362),
.B(n_2346),
.Y(n_2539)
);

NOR2xp67_ASAP7_75t_L g2540 ( 
.A(n_2486),
.B(n_2281),
.Y(n_2540)
);

AND2x2_ASAP7_75t_L g2541 ( 
.A(n_2440),
.B(n_40),
.Y(n_2541)
);

AND2x2_ASAP7_75t_L g2542 ( 
.A(n_2464),
.B(n_40),
.Y(n_2542)
);

INVx3_ASAP7_75t_L g2543 ( 
.A(n_2406),
.Y(n_2543)
);

OAI22xp5_ASAP7_75t_L g2544 ( 
.A1(n_2482),
.A2(n_2372),
.B1(n_2359),
.B2(n_2379),
.Y(n_2544)
);

INVx3_ASAP7_75t_L g2545 ( 
.A(n_2406),
.Y(n_2545)
);

NOR2xp67_ASAP7_75t_L g2546 ( 
.A(n_2487),
.B(n_2316),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_2446),
.B(n_41),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2418),
.Y(n_2548)
);

A2O1A1Ixp33_ASAP7_75t_L g2549 ( 
.A1(n_2443),
.A2(n_2348),
.B(n_1207),
.C(n_1129),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2450),
.B(n_41),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_R g2551 ( 
.A(n_2396),
.B(n_42),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2462),
.Y(n_2552)
);

A2O1A1Ixp33_ASAP7_75t_L g2553 ( 
.A1(n_2478),
.A2(n_1138),
.B(n_1166),
.C(n_1126),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2464),
.B(n_2433),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2408),
.B(n_42),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2430),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2437),
.B(n_2457),
.Y(n_2557)
);

NOR3xp33_ASAP7_75t_L g2558 ( 
.A(n_2465),
.B(n_1202),
.C(n_1167),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_2399),
.B(n_43),
.Y(n_2559)
);

AND2x2_ASAP7_75t_L g2560 ( 
.A(n_2424),
.B(n_2479),
.Y(n_2560)
);

AND2x2_ASAP7_75t_L g2561 ( 
.A(n_2434),
.B(n_43),
.Y(n_2561)
);

O2A1O1Ixp33_ASAP7_75t_L g2562 ( 
.A1(n_2445),
.A2(n_47),
.B(n_45),
.C(n_46),
.Y(n_2562)
);

CKINVDCx6p67_ASAP7_75t_R g2563 ( 
.A(n_2438),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2436),
.Y(n_2564)
);

NOR2xp67_ASAP7_75t_L g2565 ( 
.A(n_2470),
.B(n_45),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2452),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_2434),
.B(n_47),
.Y(n_2567)
);

O2A1O1Ixp5_ASAP7_75t_L g2568 ( 
.A1(n_2475),
.A2(n_58),
.B(n_67),
.C(n_48),
.Y(n_2568)
);

INVx1_ASAP7_75t_SL g2569 ( 
.A(n_2456),
.Y(n_2569)
);

AOI21xp5_ASAP7_75t_SL g2570 ( 
.A1(n_2468),
.A2(n_48),
.B(n_49),
.Y(n_2570)
);

O2A1O1Ixp5_ASAP7_75t_L g2571 ( 
.A1(n_2469),
.A2(n_61),
.B(n_71),
.C(n_50),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2564),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2548),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2499),
.Y(n_2574)
);

OAI21x1_ASAP7_75t_L g2575 ( 
.A1(n_2504),
.A2(n_2417),
.B(n_2413),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2492),
.B(n_2415),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2496),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_L g2578 ( 
.A1(n_2515),
.A2(n_2461),
.B1(n_2489),
.B2(n_2483),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2522),
.B(n_2415),
.Y(n_2579)
);

OA21x2_ASAP7_75t_L g2580 ( 
.A1(n_2501),
.A2(n_2454),
.B(n_2391),
.Y(n_2580)
);

HB1xp67_ASAP7_75t_L g2581 ( 
.A(n_2552),
.Y(n_2581)
);

AO21x2_ASAP7_75t_L g2582 ( 
.A1(n_2540),
.A2(n_2454),
.B(n_2405),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2556),
.Y(n_2583)
);

INVx1_ASAP7_75t_SL g2584 ( 
.A(n_2563),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2491),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2502),
.Y(n_2586)
);

CKINVDCx5p33_ASAP7_75t_R g2587 ( 
.A(n_2497),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2521),
.Y(n_2588)
);

OAI211xp5_ASAP7_75t_L g2589 ( 
.A1(n_2562),
.A2(n_2463),
.B(n_2402),
.C(n_2420),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2519),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2514),
.Y(n_2591)
);

OAI22xp5_ASAP7_75t_L g2592 ( 
.A1(n_2512),
.A2(n_2474),
.B1(n_2484),
.B2(n_2434),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2529),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2510),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2536),
.Y(n_2595)
);

OAI21x1_ASAP7_75t_L g2596 ( 
.A1(n_2511),
.A2(n_2417),
.B(n_2413),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2566),
.Y(n_2597)
);

BUFx2_ASAP7_75t_L g2598 ( 
.A(n_2543),
.Y(n_2598)
);

OAI21x1_ASAP7_75t_L g2599 ( 
.A1(n_2539),
.A2(n_2455),
.B(n_2412),
.Y(n_2599)
);

BUFx6f_ASAP7_75t_L g2600 ( 
.A(n_2498),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2495),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2523),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2557),
.B(n_2560),
.Y(n_2603)
);

NOR2xp33_ASAP7_75t_L g2604 ( 
.A(n_2493),
.B(n_2451),
.Y(n_2604)
);

BUFx2_ASAP7_75t_L g2605 ( 
.A(n_2543),
.Y(n_2605)
);

OAI21x1_ASAP7_75t_L g2606 ( 
.A1(n_2538),
.A2(n_2411),
.B(n_2404),
.Y(n_2606)
);

INVx2_ASAP7_75t_L g2607 ( 
.A(n_2523),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2500),
.Y(n_2608)
);

INVx1_ASAP7_75t_L g2609 ( 
.A(n_2530),
.Y(n_2609)
);

AOI221xp5_ASAP7_75t_L g2610 ( 
.A1(n_2570),
.A2(n_2485),
.B1(n_2419),
.B2(n_2432),
.C(n_2488),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_2533),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2547),
.Y(n_2612)
);

INVx3_ASAP7_75t_L g2613 ( 
.A(n_2545),
.Y(n_2613)
);

BUFx2_ASAP7_75t_L g2614 ( 
.A(n_2545),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2524),
.B(n_2488),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2518),
.B(n_2410),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2517),
.Y(n_2617)
);

BUFx2_ASAP7_75t_L g2618 ( 
.A(n_2498),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2498),
.Y(n_2619)
);

INVx2_ASAP7_75t_L g2620 ( 
.A(n_2527),
.Y(n_2620)
);

INVxp67_ASAP7_75t_L g2621 ( 
.A(n_2554),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2494),
.Y(n_2622)
);

AOI22xp33_ASAP7_75t_SL g2623 ( 
.A1(n_2551),
.A2(n_54),
.B1(n_51),
.B2(n_53),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2520),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2527),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2503),
.Y(n_2626)
);

BUFx12f_ASAP7_75t_L g2627 ( 
.A(n_2555),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2506),
.A2(n_51),
.B(n_53),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2506),
.Y(n_2629)
);

BUFx2_ASAP7_75t_L g2630 ( 
.A(n_2520),
.Y(n_2630)
);

BUFx3_ASAP7_75t_L g2631 ( 
.A(n_2542),
.Y(n_2631)
);

AND2x4_ASAP7_75t_L g2632 ( 
.A(n_2503),
.B(n_56),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2565),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2537),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2516),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2565),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2569),
.B(n_2534),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2559),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2568),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2546),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2546),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2561),
.Y(n_2642)
);

CKINVDCx9p33_ASAP7_75t_R g2643 ( 
.A(n_2535),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2567),
.Y(n_2644)
);

BUFx2_ASAP7_75t_L g2645 ( 
.A(n_2528),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2540),
.B(n_2508),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2550),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2571),
.Y(n_2648)
);

BUFx6f_ASAP7_75t_L g2649 ( 
.A(n_2490),
.Y(n_2649)
);

AND2x2_ASAP7_75t_L g2650 ( 
.A(n_2541),
.B(n_56),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2620),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2573),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2573),
.Y(n_2653)
);

AND2x4_ASAP7_75t_L g2654 ( 
.A(n_2646),
.B(n_2525),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2630),
.B(n_2505),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2583),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2603),
.B(n_2531),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2583),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2598),
.B(n_2605),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2608),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2614),
.B(n_2513),
.Y(n_2661)
);

AO31x2_ASAP7_75t_L g2662 ( 
.A1(n_2620),
.A2(n_2544),
.A3(n_2549),
.B(n_2507),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2625),
.Y(n_2663)
);

INVx3_ASAP7_75t_L g2664 ( 
.A(n_2646),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2624),
.B(n_2558),
.Y(n_2665)
);

BUFx2_ASAP7_75t_L g2666 ( 
.A(n_2643),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2625),
.Y(n_2667)
);

INVx3_ASAP7_75t_L g2668 ( 
.A(n_2624),
.Y(n_2668)
);

HB1xp67_ASAP7_75t_L g2669 ( 
.A(n_2581),
.Y(n_2669)
);

HB1xp67_ASAP7_75t_L g2670 ( 
.A(n_2581),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2615),
.B(n_2553),
.Y(n_2671)
);

OAI22xp33_ASAP7_75t_L g2672 ( 
.A1(n_2592),
.A2(n_2532),
.B1(n_2526),
.B2(n_2509),
.Y(n_2672)
);

INVxp67_ASAP7_75t_SL g2673 ( 
.A(n_2629),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2594),
.B(n_57),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2576),
.B(n_2579),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2602),
.Y(n_2676)
);

OAI22xp5_ASAP7_75t_L g2677 ( 
.A1(n_2578),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2578),
.A2(n_62),
.B1(n_59),
.B2(n_61),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2601),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2576),
.B(n_2613),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2613),
.B(n_62),
.Y(n_2681)
);

AOI22xp33_ASAP7_75t_L g2682 ( 
.A1(n_2648),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_2682)
);

INVx2_ASAP7_75t_L g2683 ( 
.A(n_2602),
.Y(n_2683)
);

AND2x4_ASAP7_75t_L g2684 ( 
.A(n_2617),
.B(n_67),
.Y(n_2684)
);

BUFx3_ASAP7_75t_L g2685 ( 
.A(n_2627),
.Y(n_2685)
);

NOR2x1p5_ASAP7_75t_L g2686 ( 
.A(n_2649),
.B(n_68),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2607),
.Y(n_2687)
);

AND2x4_ASAP7_75t_SL g2688 ( 
.A(n_2649),
.B(n_68),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2607),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2574),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_2634),
.B(n_69),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2634),
.B(n_69),
.Y(n_2692)
);

OR2x2_ASAP7_75t_L g2693 ( 
.A(n_2597),
.B(n_71),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2577),
.Y(n_2694)
);

AND2x4_ASAP7_75t_L g2695 ( 
.A(n_2632),
.B(n_74),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_2651),
.Y(n_2696)
);

AND2x2_ASAP7_75t_L g2697 ( 
.A(n_2664),
.B(n_2618),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_L g2698 ( 
.A(n_2669),
.B(n_2611),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2670),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2651),
.Y(n_2700)
);

OAI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2672),
.A2(n_2628),
.B(n_2623),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2666),
.Y(n_2702)
);

INVx5_ASAP7_75t_L g2703 ( 
.A(n_2681),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2690),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2663),
.Y(n_2705)
);

INVxp67_ASAP7_75t_L g2706 ( 
.A(n_2655),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2660),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2664),
.B(n_2612),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2664),
.B(n_2629),
.Y(n_2709)
);

AND2x2_ASAP7_75t_L g2710 ( 
.A(n_2657),
.B(n_2619),
.Y(n_2710)
);

AOI22xp33_ASAP7_75t_L g2711 ( 
.A1(n_2677),
.A2(n_2648),
.B1(n_2639),
.B2(n_2623),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2663),
.Y(n_2712)
);

AND2x2_ASAP7_75t_L g2713 ( 
.A(n_2657),
.B(n_2619),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2675),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2694),
.Y(n_2715)
);

BUFx3_ASAP7_75t_L g2716 ( 
.A(n_2685),
.Y(n_2716)
);

OR2x2_ASAP7_75t_L g2717 ( 
.A(n_2679),
.B(n_2609),
.Y(n_2717)
);

OR2x2_ASAP7_75t_L g2718 ( 
.A(n_2655),
.B(n_2622),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2652),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2659),
.B(n_2637),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2653),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2693),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2656),
.Y(n_2723)
);

AND2x2_ASAP7_75t_L g2724 ( 
.A(n_2659),
.B(n_2680),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2667),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2658),
.Y(n_2726)
);

INVx3_ASAP7_75t_L g2727 ( 
.A(n_2668),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2674),
.B(n_2635),
.Y(n_2728)
);

AND2x4_ASAP7_75t_L g2729 ( 
.A(n_2680),
.B(n_2640),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2661),
.B(n_2638),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2693),
.Y(n_2731)
);

AO31x2_ASAP7_75t_L g2732 ( 
.A1(n_2667),
.A2(n_2633),
.A3(n_2636),
.B(n_2635),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2703),
.B(n_2675),
.Y(n_2733)
);

INVx1_ASAP7_75t_L g2734 ( 
.A(n_2722),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2706),
.B(n_2674),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2732),
.Y(n_2736)
);

OR2x2_ASAP7_75t_L g2737 ( 
.A(n_2718),
.B(n_2647),
.Y(n_2737)
);

INVxp67_ASAP7_75t_SL g2738 ( 
.A(n_2702),
.Y(n_2738)
);

AOI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2701),
.A2(n_2678),
.B1(n_2639),
.B2(n_2671),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2704),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2707),
.Y(n_2741)
);

INVxp67_ASAP7_75t_L g2742 ( 
.A(n_2716),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2724),
.B(n_2661),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2732),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2731),
.Y(n_2745)
);

AND2x2_ASAP7_75t_L g2746 ( 
.A(n_2724),
.B(n_2668),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2732),
.Y(n_2747)
);

INVx2_ASAP7_75t_R g2748 ( 
.A(n_2703),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2715),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2732),
.Y(n_2750)
);

NOR2x1_ASAP7_75t_R g2751 ( 
.A(n_2716),
.B(n_2645),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2714),
.B(n_2668),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2708),
.B(n_2691),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2717),
.Y(n_2754)
);

AND2x2_ASAP7_75t_L g2755 ( 
.A(n_2703),
.B(n_2714),
.Y(n_2755)
);

HB1xp67_ASAP7_75t_L g2756 ( 
.A(n_2699),
.Y(n_2756)
);

AND2x2_ASAP7_75t_L g2757 ( 
.A(n_2703),
.B(n_2685),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2703),
.B(n_2654),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2698),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2708),
.B(n_2691),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2730),
.B(n_2684),
.Y(n_2761)
);

AOI222xp33_ASAP7_75t_L g2762 ( 
.A1(n_2711),
.A2(n_2682),
.B1(n_2686),
.B2(n_2654),
.C1(n_2671),
.C2(n_2589),
.Y(n_2762)
);

INVx1_ASAP7_75t_L g2763 ( 
.A(n_2728),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2710),
.B(n_2654),
.Y(n_2764)
);

INVx2_ASAP7_75t_L g2765 ( 
.A(n_2696),
.Y(n_2765)
);

AND2x4_ASAP7_75t_L g2766 ( 
.A(n_2710),
.B(n_2713),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2696),
.Y(n_2767)
);

HB1xp67_ASAP7_75t_L g2768 ( 
.A(n_2730),
.Y(n_2768)
);

INVx2_ASAP7_75t_L g2769 ( 
.A(n_2700),
.Y(n_2769)
);

AND2x2_ASAP7_75t_L g2770 ( 
.A(n_2697),
.B(n_2673),
.Y(n_2770)
);

OAI211xp5_ASAP7_75t_L g2771 ( 
.A1(n_2739),
.A2(n_2711),
.B(n_2589),
.C(n_2709),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2766),
.B(n_2720),
.Y(n_2772)
);

AOI22xp33_ASAP7_75t_L g2773 ( 
.A1(n_2739),
.A2(n_2695),
.B1(n_2610),
.B2(n_2628),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2736),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_L g2775 ( 
.A1(n_2762),
.A2(n_2695),
.B1(n_2580),
.B2(n_2650),
.Y(n_2775)
);

OAI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2766),
.A2(n_2720),
.B1(n_2713),
.B2(n_2695),
.Y(n_2776)
);

INVxp67_ASAP7_75t_SL g2777 ( 
.A(n_2751),
.Y(n_2777)
);

HB1xp67_ASAP7_75t_L g2778 ( 
.A(n_2756),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2742),
.B(n_2584),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2740),
.Y(n_2780)
);

INVx3_ASAP7_75t_L g2781 ( 
.A(n_2766),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2741),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2736),
.Y(n_2783)
);

OAI211xp5_ASAP7_75t_L g2784 ( 
.A1(n_2738),
.A2(n_2709),
.B(n_2681),
.C(n_2727),
.Y(n_2784)
);

HB1xp67_ASAP7_75t_L g2785 ( 
.A(n_2756),
.Y(n_2785)
);

INVx2_ASAP7_75t_SL g2786 ( 
.A(n_2764),
.Y(n_2786)
);

BUFx3_ASAP7_75t_L g2787 ( 
.A(n_2757),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2749),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2744),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_2744),
.Y(n_2790)
);

OAI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2758),
.A2(n_2755),
.B(n_2768),
.Y(n_2791)
);

INVx2_ASAP7_75t_SL g2792 ( 
.A(n_2764),
.Y(n_2792)
);

AOI21x1_ASAP7_75t_L g2793 ( 
.A1(n_2734),
.A2(n_2733),
.B(n_2770),
.Y(n_2793)
);

A2O1A1Ixp33_ASAP7_75t_SL g2794 ( 
.A1(n_2759),
.A2(n_2727),
.B(n_2697),
.C(n_2665),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2745),
.Y(n_2795)
);

AO21x2_ASAP7_75t_L g2796 ( 
.A1(n_2747),
.A2(n_2721),
.B(n_2719),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2747),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2737),
.Y(n_2798)
);

BUFx2_ASAP7_75t_L g2799 ( 
.A(n_2764),
.Y(n_2799)
);

AND2x2_ASAP7_75t_L g2800 ( 
.A(n_2768),
.B(n_2729),
.Y(n_2800)
);

AOI22xp33_ASAP7_75t_L g2801 ( 
.A1(n_2735),
.A2(n_2580),
.B1(n_2604),
.B2(n_2684),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2754),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2750),
.Y(n_2803)
);

BUFx2_ASAP7_75t_L g2804 ( 
.A(n_2761),
.Y(n_2804)
);

AOI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2763),
.A2(n_2632),
.B1(n_2665),
.B2(n_2604),
.Y(n_2805)
);

OAI221xp5_ASAP7_75t_SL g2806 ( 
.A1(n_2743),
.A2(n_2753),
.B1(n_2760),
.B2(n_2770),
.C(n_2750),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2781),
.Y(n_2807)
);

BUFx3_ASAP7_75t_L g2808 ( 
.A(n_2787),
.Y(n_2808)
);

AND2x2_ASAP7_75t_L g2809 ( 
.A(n_2772),
.B(n_2743),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2778),
.B(n_2723),
.Y(n_2810)
);

OR2x2_ASAP7_75t_L g2811 ( 
.A(n_2798),
.B(n_2748),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2785),
.B(n_2726),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2781),
.B(n_2748),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2780),
.Y(n_2814)
);

OR2x2_ASAP7_75t_L g2815 ( 
.A(n_2802),
.B(n_2746),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2782),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2788),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2781),
.Y(n_2818)
);

INVxp67_ASAP7_75t_L g2819 ( 
.A(n_2779),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2799),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2787),
.Y(n_2821)
);

AND2x2_ASAP7_75t_L g2822 ( 
.A(n_2777),
.B(n_2800),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2786),
.B(n_2746),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2795),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2804),
.Y(n_2825)
);

INVx2_ASAP7_75t_L g2826 ( 
.A(n_2786),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2792),
.B(n_2752),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2771),
.B(n_2775),
.Y(n_2828)
);

AND3x2_ASAP7_75t_L g2829 ( 
.A(n_2779),
.B(n_2692),
.C(n_2684),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_2792),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2775),
.B(n_2590),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2791),
.B(n_2752),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2774),
.Y(n_2833)
);

NAND2x1_ASAP7_75t_L g2834 ( 
.A(n_2776),
.B(n_2727),
.Y(n_2834)
);

NOR2xp67_ASAP7_75t_L g2835 ( 
.A(n_2784),
.B(n_2793),
.Y(n_2835)
);

INVx2_ASAP7_75t_L g2836 ( 
.A(n_2796),
.Y(n_2836)
);

BUFx3_ASAP7_75t_L g2837 ( 
.A(n_2805),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2796),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2801),
.B(n_2729),
.Y(n_2839)
);

OR2x2_ASAP7_75t_L g2840 ( 
.A(n_2806),
.B(n_2729),
.Y(n_2840)
);

INVx1_ASAP7_75t_SL g2841 ( 
.A(n_2803),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2801),
.B(n_2587),
.Y(n_2842)
);

OR2x2_ASAP7_75t_L g2843 ( 
.A(n_2794),
.B(n_2662),
.Y(n_2843)
);

AND2x4_ASAP7_75t_L g2844 ( 
.A(n_2773),
.B(n_2688),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_2794),
.B(n_2765),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2773),
.B(n_2765),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2774),
.Y(n_2847)
);

AND2x2_ASAP7_75t_L g2848 ( 
.A(n_2783),
.B(n_2692),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2783),
.B(n_2767),
.Y(n_2849)
);

OR2x2_ASAP7_75t_L g2850 ( 
.A(n_2789),
.B(n_2662),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2789),
.B(n_2767),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2803),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2790),
.Y(n_2853)
);

INVx2_ASAP7_75t_L g2854 ( 
.A(n_2808),
.Y(n_2854)
);

NAND2xp5_ASAP7_75t_L g2855 ( 
.A(n_2819),
.B(n_2809),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2810),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2810),
.Y(n_2857)
);

INVxp67_ASAP7_75t_L g2858 ( 
.A(n_2822),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2812),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2813),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2812),
.Y(n_2861)
);

AND2x4_ASAP7_75t_L g2862 ( 
.A(n_2821),
.B(n_2643),
.Y(n_2862)
);

NOR2x1_ASAP7_75t_L g2863 ( 
.A(n_2821),
.B(n_2790),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2819),
.B(n_2797),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2823),
.B(n_2627),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2838),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2825),
.B(n_2797),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2841),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2820),
.B(n_2688),
.Y(n_2869)
);

INVx1_ASAP7_75t_L g2870 ( 
.A(n_2841),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2836),
.Y(n_2871)
);

NOR3xp33_ASAP7_75t_L g2872 ( 
.A(n_2828),
.B(n_2769),
.C(n_2599),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2829),
.B(n_2662),
.Y(n_2873)
);

AOI211xp5_ASAP7_75t_L g2874 ( 
.A1(n_2835),
.A2(n_2649),
.B(n_2596),
.C(n_2769),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2833),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2847),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2852),
.Y(n_2877)
);

AND2x2_ASAP7_75t_L g2878 ( 
.A(n_2827),
.B(n_2631),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2826),
.Y(n_2879)
);

INVx3_ASAP7_75t_L g2880 ( 
.A(n_2834),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2829),
.B(n_2662),
.Y(n_2881)
);

INVx2_ASAP7_75t_SL g2882 ( 
.A(n_2830),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2853),
.Y(n_2883)
);

OR2x2_ASAP7_75t_L g2884 ( 
.A(n_2815),
.B(n_2662),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2807),
.B(n_2676),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2818),
.B(n_2676),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2828),
.B(n_2683),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_SL g2888 ( 
.A(n_2844),
.B(n_2649),
.Y(n_2888)
);

BUFx2_ASAP7_75t_L g2889 ( 
.A(n_2832),
.Y(n_2889)
);

AND2x2_ASAP7_75t_L g2890 ( 
.A(n_2842),
.B(n_2631),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2848),
.B(n_2683),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2840),
.B(n_2642),
.Y(n_2892)
);

AND2x2_ASAP7_75t_L g2893 ( 
.A(n_2839),
.B(n_2644),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2814),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2816),
.Y(n_2895)
);

INVx1_ASAP7_75t_L g2896 ( 
.A(n_2817),
.Y(n_2896)
);

OR2x2_ASAP7_75t_L g2897 ( 
.A(n_2831),
.B(n_2687),
.Y(n_2897)
);

AOI22xp5_ASAP7_75t_L g2898 ( 
.A1(n_2844),
.A2(n_2689),
.B1(n_2687),
.B2(n_2700),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2824),
.B(n_2689),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2811),
.Y(n_2900)
);

AND2x4_ASAP7_75t_L g2901 ( 
.A(n_2837),
.B(n_2705),
.Y(n_2901)
);

AND2x2_ASAP7_75t_L g2902 ( 
.A(n_2845),
.B(n_2621),
.Y(n_2902)
);

INVxp67_ASAP7_75t_SL g2903 ( 
.A(n_2845),
.Y(n_2903)
);

CKINVDCx16_ASAP7_75t_R g2904 ( 
.A(n_2846),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2849),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2831),
.B(n_2846),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_L g2907 ( 
.A(n_2843),
.B(n_2621),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2851),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2849),
.B(n_2616),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2851),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2850),
.B(n_2600),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2810),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2810),
.Y(n_2913)
);

OR2x2_ASAP7_75t_L g2914 ( 
.A(n_2825),
.B(n_2705),
.Y(n_2914)
);

OR2x2_ASAP7_75t_L g2915 ( 
.A(n_2825),
.B(n_2712),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2810),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2810),
.Y(n_2917)
);

AND2x2_ASAP7_75t_L g2918 ( 
.A(n_2809),
.B(n_2600),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2819),
.B(n_2712),
.Y(n_2919)
);

INVx4_ASAP7_75t_L g2920 ( 
.A(n_2808),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2819),
.B(n_2725),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2862),
.B(n_2725),
.Y(n_2922)
);

NOR2x1p5_ASAP7_75t_SL g2923 ( 
.A(n_2900),
.B(n_2641),
.Y(n_2923)
);

OAI221xp5_ASAP7_75t_L g2924 ( 
.A1(n_2903),
.A2(n_2580),
.B1(n_2591),
.B2(n_2595),
.C(n_2586),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2871),
.Y(n_2925)
);

BUFx2_ASAP7_75t_L g2926 ( 
.A(n_2862),
.Y(n_2926)
);

NAND2xp33_ASAP7_75t_R g2927 ( 
.A(n_2906),
.B(n_74),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2889),
.B(n_2600),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2868),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2904),
.B(n_2582),
.Y(n_2930)
);

OR2x2_ASAP7_75t_L g2931 ( 
.A(n_2855),
.B(n_75),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2870),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2879),
.Y(n_2933)
);

INVx2_ASAP7_75t_L g2934 ( 
.A(n_2920),
.Y(n_2934)
);

OR2x2_ASAP7_75t_L g2935 ( 
.A(n_2858),
.B(n_75),
.Y(n_2935)
);

BUFx2_ASAP7_75t_L g2936 ( 
.A(n_2920),
.Y(n_2936)
);

CKINVDCx5p33_ASAP7_75t_R g2937 ( 
.A(n_2854),
.Y(n_2937)
);

NAND2xp33_ASAP7_75t_R g2938 ( 
.A(n_2880),
.B(n_76),
.Y(n_2938)
);

AND2x2_ASAP7_75t_L g2939 ( 
.A(n_2878),
.B(n_2600),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2882),
.B(n_2582),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2864),
.Y(n_2941)
);

NOR3xp33_ASAP7_75t_L g2942 ( 
.A(n_2887),
.B(n_2606),
.C(n_2575),
.Y(n_2942)
);

INVx2_ASAP7_75t_SL g2943 ( 
.A(n_2865),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2909),
.B(n_76),
.Y(n_2944)
);

INVx2_ASAP7_75t_L g2945 ( 
.A(n_2869),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_R g2946 ( 
.A(n_2856),
.B(n_2857),
.Y(n_2946)
);

AOI21xp5_ASAP7_75t_L g2947 ( 
.A1(n_2874),
.A2(n_2626),
.B(n_2593),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2866),
.Y(n_2948)
);

AND2x4_ASAP7_75t_L g2949 ( 
.A(n_2863),
.B(n_2626),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2859),
.B(n_77),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2861),
.B(n_77),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2912),
.B(n_78),
.Y(n_2952)
);

NAND2xp33_ASAP7_75t_SL g2953 ( 
.A(n_2880),
.B(n_78),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2860),
.B(n_80),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2867),
.Y(n_2955)
);

OR2x2_ASAP7_75t_L g2956 ( 
.A(n_2914),
.B(n_80),
.Y(n_2956)
);

OR2x2_ASAP7_75t_L g2957 ( 
.A(n_2915),
.B(n_2913),
.Y(n_2957)
);

AND2x2_ASAP7_75t_L g2958 ( 
.A(n_2890),
.B(n_81),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2869),
.Y(n_2959)
);

NOR2xp67_ASAP7_75t_L g2960 ( 
.A(n_2905),
.B(n_82),
.Y(n_2960)
);

INVx1_ASAP7_75t_SL g2961 ( 
.A(n_2888),
.Y(n_2961)
);

INVx1_ASAP7_75t_SL g2962 ( 
.A(n_2902),
.Y(n_2962)
);

AOI31xp33_ASAP7_75t_L g2963 ( 
.A1(n_2916),
.A2(n_85),
.A3(n_82),
.B(n_84),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_2917),
.B(n_86),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2919),
.Y(n_2965)
);

AND2x4_ASAP7_75t_L g2966 ( 
.A(n_2875),
.B(n_2588),
.Y(n_2966)
);

BUFx12f_ASAP7_75t_L g2967 ( 
.A(n_2918),
.Y(n_2967)
);

AND2x4_ASAP7_75t_L g2968 ( 
.A(n_2876),
.B(n_2588),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2901),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2908),
.B(n_87),
.Y(n_2970)
);

OR2x6_ASAP7_75t_L g2971 ( 
.A(n_2877),
.B(n_2593),
.Y(n_2971)
);

INVxp67_ASAP7_75t_L g2972 ( 
.A(n_2921),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2910),
.Y(n_2973)
);

NAND2xp33_ASAP7_75t_R g2974 ( 
.A(n_2873),
.B(n_87),
.Y(n_2974)
);

NAND2xp33_ASAP7_75t_SL g2975 ( 
.A(n_2894),
.B(n_2895),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2901),
.Y(n_2976)
);

INVxp67_ASAP7_75t_L g2977 ( 
.A(n_2896),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2883),
.Y(n_2978)
);

AND2x2_ASAP7_75t_L g2979 ( 
.A(n_2892),
.B(n_88),
.Y(n_2979)
);

INVx2_ASAP7_75t_L g2980 ( 
.A(n_2911),
.Y(n_2980)
);

HB1xp67_ASAP7_75t_L g2981 ( 
.A(n_2907),
.Y(n_2981)
);

INVx5_ASAP7_75t_L g2982 ( 
.A(n_2893),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2872),
.B(n_88),
.Y(n_2983)
);

INVx1_ASAP7_75t_SL g2984 ( 
.A(n_2884),
.Y(n_2984)
);

NAND3xp33_ASAP7_75t_L g2985 ( 
.A(n_2881),
.B(n_90),
.C(n_91),
.Y(n_2985)
);

AOI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2897),
.A2(n_2585),
.B1(n_2572),
.B2(n_94),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2899),
.B(n_92),
.Y(n_2987)
);

NOR2x1_ASAP7_75t_L g2988 ( 
.A(n_2885),
.B(n_93),
.Y(n_2988)
);

OR2x2_ASAP7_75t_L g2989 ( 
.A(n_2886),
.B(n_95),
.Y(n_2989)
);

NOR2xp33_ASAP7_75t_L g2990 ( 
.A(n_2891),
.B(n_2898),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2862),
.Y(n_2991)
);

NOR2x1p5_ASAP7_75t_L g2992 ( 
.A(n_2920),
.B(n_95),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2920),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2871),
.Y(n_2994)
);

AND2x2_ASAP7_75t_L g2995 ( 
.A(n_2862),
.B(n_96),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2871),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2862),
.B(n_96),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2871),
.Y(n_2998)
);

NAND4xp25_ASAP7_75t_L g2999 ( 
.A(n_2889),
.B(n_101),
.C(n_99),
.D(n_100),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2871),
.Y(n_3000)
);

OAI31xp33_ASAP7_75t_L g3001 ( 
.A1(n_2906),
.A2(n_2572),
.A3(n_2585),
.B(n_102),
.Y(n_3001)
);

NAND2xp33_ASAP7_75t_SL g3002 ( 
.A(n_2920),
.B(n_99),
.Y(n_3002)
);

OR2x2_ASAP7_75t_L g3003 ( 
.A(n_2855),
.B(n_101),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2904),
.B(n_103),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2871),
.Y(n_3005)
);

OR2x2_ASAP7_75t_L g3006 ( 
.A(n_2855),
.B(n_104),
.Y(n_3006)
);

INVx2_ASAP7_75t_SL g3007 ( 
.A(n_2862),
.Y(n_3007)
);

INVxp67_ASAP7_75t_SL g3008 ( 
.A(n_2858),
.Y(n_3008)
);

NOR2xp33_ASAP7_75t_L g3009 ( 
.A(n_2920),
.B(n_104),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2871),
.Y(n_3010)
);

NAND3xp33_ASAP7_75t_L g3011 ( 
.A(n_2904),
.B(n_105),
.C(n_106),
.Y(n_3011)
);

AND2x2_ASAP7_75t_L g3012 ( 
.A(n_2862),
.B(n_106),
.Y(n_3012)
);

OR2x4_ASAP7_75t_L g3013 ( 
.A(n_2855),
.B(n_108),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_3004),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2926),
.B(n_109),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2992),
.Y(n_3016)
);

OR2x2_ASAP7_75t_L g3017 ( 
.A(n_2962),
.B(n_110),
.Y(n_3017)
);

AOI221xp5_ASAP7_75t_L g3018 ( 
.A1(n_2983),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.C(n_114),
.Y(n_3018)
);

BUFx2_ASAP7_75t_L g3019 ( 
.A(n_2967),
.Y(n_3019)
);

OR2x2_ASAP7_75t_L g3020 ( 
.A(n_2933),
.B(n_111),
.Y(n_3020)
);

INVx2_ASAP7_75t_L g3021 ( 
.A(n_2936),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2956),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_3008),
.Y(n_3023)
);

HB1xp67_ASAP7_75t_L g3024 ( 
.A(n_2938),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2931),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_3003),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_3006),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2963),
.B(n_114),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_L g3029 ( 
.A(n_2979),
.B(n_115),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_2955),
.B(n_2957),
.Y(n_3030)
);

INVxp67_ASAP7_75t_L g3031 ( 
.A(n_2927),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2954),
.B(n_117),
.Y(n_3032)
);

INVx2_ASAP7_75t_L g3033 ( 
.A(n_2982),
.Y(n_3033)
);

NOR3xp33_ASAP7_75t_L g3034 ( 
.A(n_3011),
.B(n_2985),
.C(n_2953),
.Y(n_3034)
);

AND2x2_ASAP7_75t_L g3035 ( 
.A(n_2991),
.B(n_117),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2958),
.B(n_118),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2935),
.Y(n_3037)
);

INVx2_ASAP7_75t_SL g3038 ( 
.A(n_2982),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2944),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2989),
.Y(n_3040)
);

INVx2_ASAP7_75t_SL g3041 ( 
.A(n_2982),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_3009),
.B(n_119),
.Y(n_3042)
);

OR2x2_ASAP7_75t_L g3043 ( 
.A(n_2929),
.B(n_120),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2970),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_3007),
.B(n_120),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2928),
.B(n_121),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2950),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2951),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_2952),
.Y(n_3049)
);

INVx2_ASAP7_75t_L g3050 ( 
.A(n_2937),
.Y(n_3050)
);

OR2x2_ASAP7_75t_L g3051 ( 
.A(n_2932),
.B(n_121),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2995),
.B(n_122),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2987),
.Y(n_3053)
);

OR2x2_ASAP7_75t_L g3054 ( 
.A(n_2941),
.B(n_122),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2981),
.Y(n_3055)
);

OR2x2_ASAP7_75t_L g3056 ( 
.A(n_2934),
.B(n_123),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_2993),
.B(n_124),
.Y(n_3057)
);

INVx3_ASAP7_75t_L g3058 ( 
.A(n_2945),
.Y(n_3058)
);

INVx1_ASAP7_75t_L g3059 ( 
.A(n_3013),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2997),
.B(n_125),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2988),
.Y(n_3061)
);

INVx3_ASAP7_75t_L g3062 ( 
.A(n_2959),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2969),
.Y(n_3063)
);

AOI22xp33_ASAP7_75t_L g3064 ( 
.A1(n_2942),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_3012),
.B(n_127),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2976),
.Y(n_3066)
);

NOR2xp33_ASAP7_75t_L g3067 ( 
.A(n_2999),
.B(n_128),
.Y(n_3067)
);

INVx2_ASAP7_75t_SL g3068 ( 
.A(n_2922),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2948),
.Y(n_3069)
);

AND2x2_ASAP7_75t_L g3070 ( 
.A(n_2961),
.B(n_2943),
.Y(n_3070)
);

INVx2_ASAP7_75t_L g3071 ( 
.A(n_2949),
.Y(n_3071)
);

NOR2xp33_ASAP7_75t_L g3072 ( 
.A(n_3002),
.B(n_129),
.Y(n_3072)
);

INVx1_ASAP7_75t_L g3073 ( 
.A(n_2960),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2925),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_2946),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2964),
.B(n_129),
.Y(n_3076)
);

BUFx2_ASAP7_75t_L g3077 ( 
.A(n_2975),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2994),
.Y(n_3078)
);

OR2x2_ASAP7_75t_L g3079 ( 
.A(n_2965),
.B(n_130),
.Y(n_3079)
);

NAND2xp33_ASAP7_75t_L g3080 ( 
.A(n_2980),
.B(n_2939),
.Y(n_3080)
);

OR2x2_ASAP7_75t_L g3081 ( 
.A(n_2977),
.B(n_131),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2996),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2984),
.B(n_132),
.Y(n_3083)
);

AND2x2_ASAP7_75t_L g3084 ( 
.A(n_2973),
.B(n_132),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2978),
.B(n_133),
.Y(n_3085)
);

INVx1_ASAP7_75t_L g3086 ( 
.A(n_2998),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2972),
.B(n_134),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_3000),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2990),
.B(n_134),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_3005),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3010),
.B(n_135),
.Y(n_3091)
);

A2O1A1Ixp33_ASAP7_75t_L g3092 ( 
.A1(n_2923),
.A2(n_138),
.B(n_136),
.C(n_137),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2966),
.B(n_137),
.Y(n_3093)
);

INVx1_ASAP7_75t_SL g3094 ( 
.A(n_2930),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2966),
.B(n_138),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2968),
.B(n_139),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2968),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2971),
.Y(n_3098)
);

INVxp67_ASAP7_75t_L g3099 ( 
.A(n_2974),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_2949),
.B(n_2971),
.Y(n_3100)
);

INVx1_ASAP7_75t_SL g3101 ( 
.A(n_2940),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_3001),
.B(n_2986),
.Y(n_3102)
);

AND2x2_ASAP7_75t_SL g3103 ( 
.A(n_2924),
.B(n_140),
.Y(n_3103)
);

NAND2x1p5_ASAP7_75t_L g3104 ( 
.A(n_2947),
.B(n_140),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2992),
.Y(n_3105)
);

A2O1A1Ixp33_ASAP7_75t_L g3106 ( 
.A1(n_2983),
.A2(n_143),
.B(n_141),
.C(n_142),
.Y(n_3106)
);

NOR2xp33_ASAP7_75t_L g3107 ( 
.A(n_3013),
.B(n_141),
.Y(n_3107)
);

OR2x2_ASAP7_75t_L g3108 ( 
.A(n_2962),
.B(n_143),
.Y(n_3108)
);

NOR3xp33_ASAP7_75t_L g3109 ( 
.A(n_3004),
.B(n_144),
.C(n_145),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2926),
.B(n_145),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2992),
.Y(n_3111)
);

INVxp67_ASAP7_75t_SL g3112 ( 
.A(n_2938),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_3004),
.Y(n_3113)
);

NAND2xp5_ASAP7_75t_L g3114 ( 
.A(n_2963),
.B(n_146),
.Y(n_3114)
);

INVx1_ASAP7_75t_SL g3115 ( 
.A(n_2953),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2963),
.B(n_147),
.Y(n_3116)
);

NOR2xp33_ASAP7_75t_L g3117 ( 
.A(n_3013),
.B(n_148),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2926),
.B(n_148),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_3004),
.Y(n_3119)
);

NOR2xp33_ASAP7_75t_L g3120 ( 
.A(n_3013),
.B(n_150),
.Y(n_3120)
);

NAND2x1p5_ASAP7_75t_L g3121 ( 
.A(n_2936),
.B(n_150),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_3004),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_3004),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2926),
.B(n_151),
.Y(n_3124)
);

INVxp67_ASAP7_75t_L g3125 ( 
.A(n_2938),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2963),
.B(n_151),
.Y(n_3126)
);

AOI21xp33_ASAP7_75t_L g3127 ( 
.A1(n_2927),
.A2(n_152),
.B(n_153),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2963),
.B(n_152),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2963),
.B(n_154),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2963),
.B(n_155),
.Y(n_3130)
);

OAI21xp33_ASAP7_75t_L g3131 ( 
.A1(n_3007),
.A2(n_156),
.B(n_157),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2963),
.B(n_156),
.Y(n_3132)
);

AND2x2_ASAP7_75t_L g3133 ( 
.A(n_2926),
.B(n_158),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_3004),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2926),
.B(n_159),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2963),
.B(n_160),
.Y(n_3136)
);

INVx1_ASAP7_75t_L g3137 ( 
.A(n_3004),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2963),
.B(n_160),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2926),
.B(n_161),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2926),
.B(n_161),
.Y(n_3140)
);

NOR2xp33_ASAP7_75t_L g3141 ( 
.A(n_3013),
.B(n_165),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2963),
.B(n_165),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2963),
.B(n_166),
.Y(n_3143)
);

HB1xp67_ASAP7_75t_L g3144 ( 
.A(n_2992),
.Y(n_3144)
);

OR2x2_ASAP7_75t_L g3145 ( 
.A(n_2962),
.B(n_166),
.Y(n_3145)
);

INVx1_ASAP7_75t_L g3146 ( 
.A(n_3004),
.Y(n_3146)
);

AND2x2_ASAP7_75t_L g3147 ( 
.A(n_2926),
.B(n_167),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2992),
.Y(n_3148)
);

NOR2xp67_ASAP7_75t_L g3149 ( 
.A(n_2982),
.B(n_167),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2963),
.B(n_169),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2926),
.B(n_169),
.Y(n_3151)
);

INVx1_ASAP7_75t_L g3152 ( 
.A(n_3004),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_3004),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2992),
.Y(n_3154)
);

AND2x2_ASAP7_75t_L g3155 ( 
.A(n_2926),
.B(n_170),
.Y(n_3155)
);

OR2x2_ASAP7_75t_L g3156 ( 
.A(n_2962),
.B(n_170),
.Y(n_3156)
);

NAND2xp5_ASAP7_75t_L g3157 ( 
.A(n_2963),
.B(n_171),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_L g3158 ( 
.A(n_2963),
.B(n_172),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2963),
.B(n_173),
.Y(n_3159)
);

HB1xp67_ASAP7_75t_L g3160 ( 
.A(n_2992),
.Y(n_3160)
);

NAND4xp25_ASAP7_75t_SL g3161 ( 
.A(n_2961),
.B(n_177),
.C(n_174),
.D(n_176),
.Y(n_3161)
);

AND2x2_ASAP7_75t_L g3162 ( 
.A(n_2926),
.B(n_177),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2926),
.B(n_178),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_3004),
.Y(n_3164)
);

NAND2x1p5_ASAP7_75t_L g3165 ( 
.A(n_2936),
.B(n_179),
.Y(n_3165)
);

OR2x2_ASAP7_75t_L g3166 ( 
.A(n_2962),
.B(n_179),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3004),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_L g3168 ( 
.A(n_3013),
.B(n_180),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_3077),
.A2(n_181),
.B(n_182),
.Y(n_3169)
);

OAI221xp5_ASAP7_75t_L g3170 ( 
.A1(n_3064),
.A2(n_185),
.B1(n_181),
.B2(n_182),
.C(n_187),
.Y(n_3170)
);

NOR3xp33_ASAP7_75t_L g3171 ( 
.A(n_3125),
.B(n_185),
.C(n_187),
.Y(n_3171)
);

OAI21xp5_ASAP7_75t_L g3172 ( 
.A1(n_3099),
.A2(n_188),
.B(n_189),
.Y(n_3172)
);

OAI22xp33_ASAP7_75t_L g3173 ( 
.A1(n_3115),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_3121),
.Y(n_3174)
);

INVx1_ASAP7_75t_SL g3175 ( 
.A(n_3070),
.Y(n_3175)
);

NAND3xp33_ASAP7_75t_L g3176 ( 
.A(n_3075),
.B(n_3024),
.C(n_3059),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_3028),
.A2(n_194),
.B(n_195),
.Y(n_3177)
);

OR2x2_ASAP7_75t_L g3178 ( 
.A(n_3030),
.B(n_194),
.Y(n_3178)
);

AOI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_3112),
.A2(n_3031),
.B1(n_3105),
.B2(n_3016),
.Y(n_3179)
);

OAI33xp33_ASAP7_75t_L g3180 ( 
.A1(n_3063),
.A2(n_197),
.A3(n_200),
.B1(n_195),
.B2(n_196),
.B3(n_198),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_3058),
.Y(n_3181)
);

AOI221xp5_ASAP7_75t_L g3182 ( 
.A1(n_3061),
.A2(n_201),
.B1(n_198),
.B2(n_200),
.C(n_203),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3058),
.Y(n_3183)
);

AOI322xp5_ASAP7_75t_L g3184 ( 
.A1(n_3034),
.A2(n_211),
.A3(n_210),
.B1(n_208),
.B2(n_204),
.C1(n_206),
.C2(n_209),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3149),
.B(n_208),
.Y(n_3185)
);

NOR2xp33_ASAP7_75t_L g3186 ( 
.A(n_3019),
.B(n_3050),
.Y(n_3186)
);

OAI21xp5_ASAP7_75t_L g3187 ( 
.A1(n_3106),
.A2(n_209),
.B(n_211),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3062),
.B(n_212),
.Y(n_3188)
);

AOI221xp5_ASAP7_75t_L g3189 ( 
.A1(n_3094),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.C(n_216),
.Y(n_3189)
);

XNOR2x1_ASAP7_75t_L g3190 ( 
.A(n_3111),
.B(n_216),
.Y(n_3190)
);

AOI221xp5_ASAP7_75t_L g3191 ( 
.A1(n_3014),
.A2(n_3167),
.B1(n_3164),
.B2(n_3127),
.C(n_3160),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_3062),
.B(n_218),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3015),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_3110),
.B(n_218),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3118),
.Y(n_3195)
);

NAND2xp33_ASAP7_75t_SL g3196 ( 
.A(n_3068),
.B(n_220),
.Y(n_3196)
);

A2O1A1Ixp33_ASAP7_75t_L g3197 ( 
.A1(n_3072),
.A2(n_222),
.B(n_220),
.C(n_221),
.Y(n_3197)
);

BUFx2_ASAP7_75t_L g3198 ( 
.A(n_3165),
.Y(n_3198)
);

AOI222xp33_ASAP7_75t_L g3199 ( 
.A1(n_3103),
.A2(n_224),
.B1(n_226),
.B2(n_222),
.C1(n_223),
.C2(n_225),
.Y(n_3199)
);

AOI21xp5_ASAP7_75t_L g3200 ( 
.A1(n_3114),
.A2(n_225),
.B(n_226),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3124),
.B(n_227),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3133),
.Y(n_3202)
);

NOR2xp33_ASAP7_75t_R g3203 ( 
.A(n_3055),
.B(n_227),
.Y(n_3203)
);

AO32x1_ASAP7_75t_L g3204 ( 
.A1(n_3038),
.A2(n_230),
.A3(n_228),
.B1(n_229),
.B2(n_231),
.Y(n_3204)
);

AOI22xp5_ASAP7_75t_L g3205 ( 
.A1(n_3148),
.A2(n_3154),
.B1(n_3164),
.B2(n_3014),
.Y(n_3205)
);

OAI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3023),
.A2(n_3144),
.B1(n_3041),
.B2(n_3108),
.Y(n_3206)
);

NOR2xp67_ASAP7_75t_L g3207 ( 
.A(n_3161),
.B(n_228),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3135),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3139),
.B(n_229),
.Y(n_3209)
);

OA211x2_ASAP7_75t_L g3210 ( 
.A1(n_3131),
.A2(n_233),
.B(n_230),
.C(n_232),
.Y(n_3210)
);

AOI21xp33_ASAP7_75t_L g3211 ( 
.A1(n_3073),
.A2(n_3026),
.B(n_3025),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3140),
.B(n_232),
.Y(n_3212)
);

INVx2_ASAP7_75t_SL g3213 ( 
.A(n_3147),
.Y(n_3213)
);

OAI21xp33_ASAP7_75t_L g3214 ( 
.A1(n_3080),
.A2(n_233),
.B(n_234),
.Y(n_3214)
);

OAI222xp33_ASAP7_75t_L g3215 ( 
.A1(n_3104),
.A2(n_236),
.B1(n_239),
.B2(n_234),
.C1(n_235),
.C2(n_238),
.Y(n_3215)
);

INVxp67_ASAP7_75t_L g3216 ( 
.A(n_3151),
.Y(n_3216)
);

INVx1_ASAP7_75t_SL g3217 ( 
.A(n_3155),
.Y(n_3217)
);

AOI22xp5_ASAP7_75t_L g3218 ( 
.A1(n_3167),
.A2(n_240),
.B1(n_236),
.B2(n_238),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_3162),
.Y(n_3219)
);

AOI211xp5_ASAP7_75t_L g3220 ( 
.A1(n_3113),
.A2(n_242),
.B(n_240),
.C(n_241),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_3163),
.Y(n_3221)
);

OAI22xp5_ASAP7_75t_L g3222 ( 
.A1(n_3017),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_3222)
);

AOI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_3119),
.A2(n_248),
.B1(n_243),
.B2(n_247),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3107),
.B(n_247),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3145),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_SL g3226 ( 
.A(n_3021),
.B(n_248),
.Y(n_3226)
);

NOR4xp25_ASAP7_75t_L g3227 ( 
.A(n_3066),
.B(n_251),
.C(n_249),
.D(n_250),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3156),
.Y(n_3228)
);

OAI221xp5_ASAP7_75t_L g3229 ( 
.A1(n_3092),
.A2(n_252),
.B1(n_249),
.B2(n_251),
.C(n_253),
.Y(n_3229)
);

OAI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_3166),
.A2(n_254),
.B1(n_252),
.B2(n_253),
.Y(n_3230)
);

AOI22xp5_ASAP7_75t_L g3231 ( 
.A1(n_3122),
.A2(n_258),
.B1(n_256),
.B2(n_257),
.Y(n_3231)
);

NAND2xp5_ASAP7_75t_L g3232 ( 
.A(n_3117),
.B(n_257),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_3120),
.B(n_259),
.Y(n_3233)
);

AOI22xp5_ASAP7_75t_L g3234 ( 
.A1(n_3123),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_3234)
);

INVx2_ASAP7_75t_L g3235 ( 
.A(n_3052),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3141),
.B(n_260),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3054),
.Y(n_3237)
);

AOI21xp5_ASAP7_75t_L g3238 ( 
.A1(n_3116),
.A2(n_262),
.B(n_263),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3091),
.Y(n_3239)
);

AND2x2_ASAP7_75t_L g3240 ( 
.A(n_3046),
.B(n_3045),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_3060),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_3065),
.Y(n_3242)
);

INVxp67_ASAP7_75t_SL g3243 ( 
.A(n_3126),
.Y(n_3243)
);

AOI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3134),
.A2(n_264),
.B1(n_262),
.B2(n_263),
.Y(n_3244)
);

OAI21xp5_ASAP7_75t_SL g3245 ( 
.A1(n_3033),
.A2(n_265),
.B(n_266),
.Y(n_3245)
);

NOR2xp67_ASAP7_75t_L g3246 ( 
.A(n_3020),
.B(n_265),
.Y(n_3246)
);

AOI222xp33_ASAP7_75t_L g3247 ( 
.A1(n_3101),
.A2(n_268),
.B1(n_270),
.B2(n_266),
.C1(n_267),
.C2(n_269),
.Y(n_3247)
);

NAND2x1_ASAP7_75t_L g3248 ( 
.A(n_3035),
.B(n_267),
.Y(n_3248)
);

AOI22xp5_ASAP7_75t_L g3249 ( 
.A1(n_3137),
.A2(n_273),
.B1(n_268),
.B2(n_272),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_SL g3250 ( 
.A(n_3071),
.B(n_274),
.Y(n_3250)
);

AOI221xp5_ASAP7_75t_L g3251 ( 
.A1(n_3146),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.C(n_277),
.Y(n_3251)
);

OAI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_3083),
.A2(n_275),
.B(n_277),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_3084),
.Y(n_3253)
);

OAI31xp33_ASAP7_75t_L g3254 ( 
.A1(n_3089),
.A2(n_281),
.A3(n_278),
.B(n_280),
.Y(n_3254)
);

AOI311xp33_ASAP7_75t_L g3255 ( 
.A1(n_3069),
.A2(n_282),
.A3(n_278),
.B(n_280),
.C(n_283),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3029),
.Y(n_3256)
);

INVxp67_ASAP7_75t_L g3257 ( 
.A(n_3168),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3085),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_3079),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3036),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3043),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3051),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3128),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3129),
.Y(n_3264)
);

AOI22xp5_ASAP7_75t_L g3265 ( 
.A1(n_3152),
.A2(n_284),
.B1(n_282),
.B2(n_283),
.Y(n_3265)
);

NOR3xp33_ASAP7_75t_L g3266 ( 
.A(n_3153),
.B(n_284),
.C(n_285),
.Y(n_3266)
);

OAI322xp33_ASAP7_75t_L g3267 ( 
.A1(n_3074),
.A2(n_285),
.A3(n_286),
.B1(n_287),
.B2(n_289),
.C1(n_291),
.C2(n_292),
.Y(n_3267)
);

NOR4xp25_ASAP7_75t_L g3268 ( 
.A(n_3037),
.B(n_294),
.C(n_286),
.D(n_287),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3027),
.B(n_294),
.Y(n_3269)
);

NAND2xp5_ASAP7_75t_L g3270 ( 
.A(n_3095),
.B(n_295),
.Y(n_3270)
);

AOI21xp33_ASAP7_75t_L g3271 ( 
.A1(n_3040),
.A2(n_295),
.B(n_297),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3130),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3078),
.B(n_297),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3132),
.Y(n_3274)
);

NOR2xp67_ASAP7_75t_L g3275 ( 
.A(n_3081),
.B(n_298),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3136),
.Y(n_3276)
);

INVx1_ASAP7_75t_SL g3277 ( 
.A(n_3138),
.Y(n_3277)
);

INVxp67_ASAP7_75t_L g3278 ( 
.A(n_3142),
.Y(n_3278)
);

AOI22xp33_ASAP7_75t_L g3279 ( 
.A1(n_3022),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_3279)
);

INVxp67_ASAP7_75t_L g3280 ( 
.A(n_3143),
.Y(n_3280)
);

OAI222xp33_ASAP7_75t_L g3281 ( 
.A1(n_3102),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.C1(n_305),
.C2(n_306),
.Y(n_3281)
);

INVxp67_ASAP7_75t_L g3282 ( 
.A(n_3150),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_3157),
.Y(n_3283)
);

INVxp33_ASAP7_75t_SL g3284 ( 
.A(n_3067),
.Y(n_3284)
);

NOR2x1_ASAP7_75t_L g3285 ( 
.A(n_3158),
.B(n_305),
.Y(n_3285)
);

AOI321xp33_ASAP7_75t_L g3286 ( 
.A1(n_3100),
.A2(n_3098),
.A3(n_3097),
.B1(n_3090),
.B2(n_3086),
.C(n_3088),
.Y(n_3286)
);

OAI211xp5_ASAP7_75t_L g3287 ( 
.A1(n_3082),
.A2(n_3047),
.B(n_3048),
.C(n_3044),
.Y(n_3287)
);

NAND2xp33_ASAP7_75t_SL g3288 ( 
.A(n_3159),
.B(n_307),
.Y(n_3288)
);

INVx2_ASAP7_75t_SL g3289 ( 
.A(n_3056),
.Y(n_3289)
);

NOR3xp33_ASAP7_75t_SL g3290 ( 
.A(n_3049),
.B(n_308),
.C(n_309),
.Y(n_3290)
);

AOI21xp33_ASAP7_75t_L g3291 ( 
.A1(n_3039),
.A2(n_3053),
.B(n_3098),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3204),
.Y(n_3292)
);

AOI21xp33_ASAP7_75t_SL g3293 ( 
.A1(n_3213),
.A2(n_3057),
.B(n_3087),
.Y(n_3293)
);

OAI21xp33_ASAP7_75t_L g3294 ( 
.A1(n_3179),
.A2(n_3076),
.B(n_3042),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3204),
.Y(n_3295)
);

AND2x2_ASAP7_75t_L g3296 ( 
.A(n_3175),
.B(n_3109),
.Y(n_3296)
);

NAND4xp25_ASAP7_75t_L g3297 ( 
.A(n_3286),
.B(n_3018),
.C(n_3096),
.D(n_3093),
.Y(n_3297)
);

AND2x2_ASAP7_75t_L g3298 ( 
.A(n_3198),
.B(n_3032),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_3240),
.B(n_309),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3204),
.Y(n_3300)
);

OAI221xp5_ASAP7_75t_L g3301 ( 
.A1(n_3243),
.A2(n_313),
.B1(n_310),
.B2(n_311),
.C(n_314),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3178),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_L g3303 ( 
.A1(n_3263),
.A2(n_316),
.B1(n_314),
.B2(n_315),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3181),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3268),
.B(n_3227),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3183),
.Y(n_3306)
);

AND2x2_ASAP7_75t_SL g3307 ( 
.A(n_3186),
.B(n_315),
.Y(n_3307)
);

AND2x2_ASAP7_75t_L g3308 ( 
.A(n_3174),
.B(n_317),
.Y(n_3308)
);

INVx1_ASAP7_75t_L g3309 ( 
.A(n_3185),
.Y(n_3309)
);

INVx2_ASAP7_75t_L g3310 ( 
.A(n_3248),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_3207),
.B(n_318),
.Y(n_3311)
);

INVx1_ASAP7_75t_L g3312 ( 
.A(n_3194),
.Y(n_3312)
);

INVx2_ASAP7_75t_SL g3313 ( 
.A(n_3273),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3190),
.Y(n_3314)
);

INVx2_ASAP7_75t_L g3315 ( 
.A(n_3235),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3206),
.B(n_3217),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3201),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3241),
.B(n_318),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_3242),
.B(n_319),
.Y(n_3319)
);

OR2x2_ASAP7_75t_L g3320 ( 
.A(n_3176),
.B(n_321),
.Y(n_3320)
);

AND2x2_ASAP7_75t_L g3321 ( 
.A(n_3255),
.B(n_3264),
.Y(n_3321)
);

NAND2xp5_ASAP7_75t_L g3322 ( 
.A(n_3289),
.B(n_3290),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3193),
.B(n_321),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_L g3324 ( 
.A(n_3195),
.B(n_322),
.Y(n_3324)
);

AND2x2_ASAP7_75t_L g3325 ( 
.A(n_3272),
.B(n_322),
.Y(n_3325)
);

INVx2_ASAP7_75t_SL g3326 ( 
.A(n_3226),
.Y(n_3326)
);

OR2x2_ASAP7_75t_L g3327 ( 
.A(n_3202),
.B(n_323),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3208),
.B(n_324),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3219),
.B(n_325),
.Y(n_3329)
);

NOR2xp33_ASAP7_75t_L g3330 ( 
.A(n_3180),
.B(n_326),
.Y(n_3330)
);

INVx1_ASAP7_75t_SL g3331 ( 
.A(n_3196),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3209),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3212),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3188),
.Y(n_3334)
);

NAND2xp33_ASAP7_75t_R g3335 ( 
.A(n_3203),
.B(n_327),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_L g3336 ( 
.A(n_3221),
.B(n_327),
.Y(n_3336)
);

OAI21xp5_ASAP7_75t_SL g3337 ( 
.A1(n_3211),
.A2(n_328),
.B(n_329),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_3191),
.B(n_328),
.Y(n_3338)
);

OR2x2_ASAP7_75t_L g3339 ( 
.A(n_3192),
.B(n_330),
.Y(n_3339)
);

INVx1_ASAP7_75t_SL g3340 ( 
.A(n_3288),
.Y(n_3340)
);

AND2x2_ASAP7_75t_L g3341 ( 
.A(n_3274),
.B(n_331),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3285),
.Y(n_3342)
);

NAND2x1_ASAP7_75t_SL g3343 ( 
.A(n_3205),
.B(n_331),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_3276),
.B(n_334),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_3246),
.Y(n_3345)
);

INVxp67_ASAP7_75t_L g3346 ( 
.A(n_3275),
.Y(n_3346)
);

INVxp33_ASAP7_75t_L g3347 ( 
.A(n_3171),
.Y(n_3347)
);

OAI22xp33_ASAP7_75t_L g3348 ( 
.A1(n_3277),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_3210),
.Y(n_3349)
);

AND2x2_ASAP7_75t_L g3350 ( 
.A(n_3283),
.B(n_335),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_3216),
.B(n_336),
.Y(n_3351)
);

OR2x2_ASAP7_75t_L g3352 ( 
.A(n_3269),
.B(n_337),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3245),
.B(n_3239),
.Y(n_3353)
);

INVx2_ASAP7_75t_SL g3354 ( 
.A(n_3253),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3258),
.B(n_3225),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3228),
.Y(n_3356)
);

OAI21xp5_ASAP7_75t_SL g3357 ( 
.A1(n_3287),
.A2(n_337),
.B(n_338),
.Y(n_3357)
);

AND2x2_ASAP7_75t_L g3358 ( 
.A(n_3172),
.B(n_339),
.Y(n_3358)
);

INVx2_ASAP7_75t_SL g3359 ( 
.A(n_3270),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3237),
.B(n_340),
.Y(n_3360)
);

OR2x2_ASAP7_75t_L g3361 ( 
.A(n_3278),
.B(n_340),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3259),
.B(n_341),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3261),
.Y(n_3363)
);

NOR2x1_ASAP7_75t_L g3364 ( 
.A(n_3173),
.B(n_341),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3262),
.Y(n_3365)
);

INVx1_ASAP7_75t_L g3366 ( 
.A(n_3256),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3260),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3267),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3247),
.B(n_342),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_SL g3370 ( 
.A(n_3169),
.B(n_342),
.Y(n_3370)
);

AND2x2_ASAP7_75t_SL g3371 ( 
.A(n_3266),
.B(n_343),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3224),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3280),
.B(n_343),
.Y(n_3373)
);

INVx3_ASAP7_75t_L g3374 ( 
.A(n_3232),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3233),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_3236),
.Y(n_3376)
);

OAI21xp5_ASAP7_75t_L g3377 ( 
.A1(n_3177),
.A2(n_344),
.B(n_345),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3200),
.B(n_344),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_3222),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3282),
.B(n_346),
.Y(n_3380)
);

AND2x2_ASAP7_75t_L g3381 ( 
.A(n_3214),
.B(n_346),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_3189),
.B(n_347),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3238),
.B(n_348),
.Y(n_3383)
);

AND2x2_ASAP7_75t_L g3384 ( 
.A(n_3252),
.B(n_348),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3230),
.Y(n_3385)
);

CKINVDCx14_ASAP7_75t_R g3386 ( 
.A(n_3223),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3218),
.Y(n_3387)
);

NAND2xp5_ASAP7_75t_L g3388 ( 
.A(n_3254),
.B(n_349),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3220),
.B(n_350),
.Y(n_3389)
);

NAND2xp5_ASAP7_75t_L g3390 ( 
.A(n_3184),
.B(n_351),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3231),
.Y(n_3391)
);

NAND2x1p5_ASAP7_75t_L g3392 ( 
.A(n_3250),
.B(n_352),
.Y(n_3392)
);

OR2x2_ASAP7_75t_L g3393 ( 
.A(n_3257),
.B(n_352),
.Y(n_3393)
);

AND2x2_ASAP7_75t_L g3394 ( 
.A(n_3187),
.B(n_354),
.Y(n_3394)
);

AND2x4_ASAP7_75t_L g3395 ( 
.A(n_3197),
.B(n_355),
.Y(n_3395)
);

INVx1_ASAP7_75t_SL g3396 ( 
.A(n_3284),
.Y(n_3396)
);

INVx1_ASAP7_75t_SL g3397 ( 
.A(n_3271),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3234),
.B(n_3244),
.Y(n_3398)
);

INVx1_ASAP7_75t_L g3399 ( 
.A(n_3249),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3265),
.B(n_356),
.Y(n_3400)
);

NOR3xp33_ASAP7_75t_SL g3401 ( 
.A(n_3291),
.B(n_357),
.C(n_358),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_SL g3402 ( 
.A(n_3199),
.B(n_3182),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3229),
.Y(n_3403)
);

NAND2xp5_ASAP7_75t_L g3404 ( 
.A(n_3279),
.B(n_357),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3170),
.Y(n_3405)
);

OR2x2_ASAP7_75t_L g3406 ( 
.A(n_3281),
.B(n_359),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3251),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3215),
.B(n_360),
.Y(n_3408)
);

AND2x2_ASAP7_75t_L g3409 ( 
.A(n_3175),
.B(n_360),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3240),
.B(n_361),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3204),
.Y(n_3411)
);

INVx1_ASAP7_75t_SL g3412 ( 
.A(n_3175),
.Y(n_3412)
);

NAND2xp33_ASAP7_75t_SL g3413 ( 
.A(n_3198),
.B(n_361),
.Y(n_3413)
);

INVx1_ASAP7_75t_L g3414 ( 
.A(n_3204),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3240),
.B(n_362),
.Y(n_3415)
);

INVxp67_ASAP7_75t_SL g3416 ( 
.A(n_3216),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3204),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_3204),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_3204),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3240),
.B(n_363),
.Y(n_3420)
);

AND2x2_ASAP7_75t_L g3421 ( 
.A(n_3175),
.B(n_364),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3175),
.B(n_365),
.Y(n_3422)
);

AND2x2_ASAP7_75t_L g3423 ( 
.A(n_3175),
.B(n_367),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_3175),
.B(n_368),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3240),
.B(n_369),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3175),
.B(n_370),
.Y(n_3426)
);

NAND2x1p5_ASAP7_75t_L g3427 ( 
.A(n_3198),
.B(n_371),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3204),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3240),
.B(n_372),
.Y(n_3429)
);

BUFx2_ASAP7_75t_SL g3430 ( 
.A(n_3175),
.Y(n_3430)
);

NAND2xp33_ASAP7_75t_SL g3431 ( 
.A(n_3198),
.B(n_372),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_3204),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3204),
.Y(n_3433)
);

NAND3xp33_ASAP7_75t_L g3434 ( 
.A(n_3286),
.B(n_373),
.C(n_374),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3204),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3204),
.Y(n_3436)
);

INVxp67_ASAP7_75t_L g3437 ( 
.A(n_3198),
.Y(n_3437)
);

INVx1_ASAP7_75t_L g3438 ( 
.A(n_3204),
.Y(n_3438)
);

A2O1A1Ixp33_ASAP7_75t_L g3439 ( 
.A1(n_3177),
.A2(n_375),
.B(n_373),
.C(n_374),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3204),
.Y(n_3440)
);

OAI22xp5_ASAP7_75t_L g3441 ( 
.A1(n_3175),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_3441)
);

INVxp67_ASAP7_75t_SL g3442 ( 
.A(n_3216),
.Y(n_3442)
);

INVx1_ASAP7_75t_SL g3443 ( 
.A(n_3175),
.Y(n_3443)
);

AND2x2_ASAP7_75t_L g3444 ( 
.A(n_3175),
.B(n_376),
.Y(n_3444)
);

INVx2_ASAP7_75t_SL g3445 ( 
.A(n_3427),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3412),
.B(n_378),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_3307),
.B(n_379),
.Y(n_3447)
);

OAI21xp33_ASAP7_75t_L g3448 ( 
.A1(n_3443),
.A2(n_379),
.B(n_381),
.Y(n_3448)
);

XOR2xp5_ASAP7_75t_L g3449 ( 
.A(n_3314),
.B(n_3430),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3310),
.B(n_382),
.Y(n_3450)
);

NOR3xp33_ASAP7_75t_SL g3451 ( 
.A(n_3434),
.B(n_382),
.C(n_384),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3406),
.Y(n_3452)
);

OAI21xp33_ASAP7_75t_L g3453 ( 
.A1(n_3294),
.A2(n_384),
.B(n_386),
.Y(n_3453)
);

AND2x2_ASAP7_75t_L g3454 ( 
.A(n_3316),
.B(n_387),
.Y(n_3454)
);

OAI211xp5_ASAP7_75t_L g3455 ( 
.A1(n_3357),
.A2(n_389),
.B(n_387),
.C(n_388),
.Y(n_3455)
);

A2O1A1Ixp33_ASAP7_75t_L g3456 ( 
.A1(n_3330),
.A2(n_3305),
.B(n_3440),
.C(n_3292),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3409),
.Y(n_3457)
);

NAND2xp33_ASAP7_75t_SL g3458 ( 
.A(n_3354),
.B(n_388),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_3343),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3313),
.B(n_390),
.Y(n_3460)
);

INVx3_ASAP7_75t_SL g3461 ( 
.A(n_3396),
.Y(n_3461)
);

NOR2xp33_ASAP7_75t_L g3462 ( 
.A(n_3331),
.B(n_390),
.Y(n_3462)
);

INVx1_ASAP7_75t_SL g3463 ( 
.A(n_3413),
.Y(n_3463)
);

AOI21xp33_ASAP7_75t_L g3464 ( 
.A1(n_3335),
.A2(n_391),
.B(n_394),
.Y(n_3464)
);

AND2x4_ASAP7_75t_L g3465 ( 
.A(n_3298),
.B(n_394),
.Y(n_3465)
);

BUFx3_ASAP7_75t_L g3466 ( 
.A(n_3421),
.Y(n_3466)
);

A2O1A1Ixp33_ASAP7_75t_L g3467 ( 
.A1(n_3292),
.A2(n_399),
.B(n_395),
.C(n_397),
.Y(n_3467)
);

NAND2xp5_ASAP7_75t_L g3468 ( 
.A(n_3340),
.B(n_399),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3422),
.Y(n_3469)
);

INVx1_ASAP7_75t_SL g3470 ( 
.A(n_3431),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3423),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_3426),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3444),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3342),
.Y(n_3474)
);

INVx1_ASAP7_75t_SL g3475 ( 
.A(n_3296),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_3401),
.B(n_3374),
.Y(n_3476)
);

NOR2xp33_ASAP7_75t_L g3477 ( 
.A(n_3392),
.B(n_400),
.Y(n_3477)
);

OAI211xp5_ASAP7_75t_L g3478 ( 
.A1(n_3437),
.A2(n_402),
.B(n_400),
.C(n_401),
.Y(n_3478)
);

HB1xp67_ASAP7_75t_L g3479 ( 
.A(n_3440),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3299),
.Y(n_3480)
);

NOR2xp33_ASAP7_75t_L g3481 ( 
.A(n_3337),
.B(n_401),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_3374),
.B(n_3302),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3410),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_L g3484 ( 
.A(n_3349),
.B(n_403),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_L g3485 ( 
.A(n_3311),
.B(n_403),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_3415),
.Y(n_3486)
);

INVxp67_ASAP7_75t_SL g3487 ( 
.A(n_3322),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3325),
.B(n_404),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3327),
.Y(n_3489)
);

AND2x2_ASAP7_75t_SL g3490 ( 
.A(n_3371),
.B(n_404),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3420),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_R g3492 ( 
.A(n_3320),
.B(n_408),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3341),
.B(n_408),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3425),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_3429),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3344),
.B(n_3350),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3295),
.B(n_410),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3300),
.B(n_410),
.Y(n_3498)
);

NOR4xp25_ASAP7_75t_SL g3499 ( 
.A(n_3338),
.B(n_414),
.C(n_411),
.D(n_412),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3411),
.B(n_411),
.Y(n_3500)
);

OR2x2_ASAP7_75t_L g3501 ( 
.A(n_3353),
.B(n_412),
.Y(n_3501)
);

XNOR2xp5_ASAP7_75t_L g3502 ( 
.A(n_3297),
.B(n_415),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3378),
.Y(n_3503)
);

A2O1A1Ixp33_ASAP7_75t_L g3504 ( 
.A1(n_3414),
.A2(n_418),
.B(n_415),
.C(n_416),
.Y(n_3504)
);

XOR2x2_ASAP7_75t_L g3505 ( 
.A(n_3364),
.B(n_416),
.Y(n_3505)
);

NAND3xp33_ASAP7_75t_L g3506 ( 
.A(n_3417),
.B(n_419),
.C(n_420),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3383),
.Y(n_3507)
);

NOR3xp33_ASAP7_75t_L g3508 ( 
.A(n_3346),
.B(n_421),
.C(n_422),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_L g3509 ( 
.A(n_3418),
.B(n_421),
.Y(n_3509)
);

HB1xp67_ASAP7_75t_L g3510 ( 
.A(n_3315),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_SL g3511 ( 
.A1(n_3419),
.A2(n_426),
.B1(n_422),
.B2(n_424),
.Y(n_3511)
);

NOR2xp33_ASAP7_75t_L g3512 ( 
.A(n_3347),
.B(n_424),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3408),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3352),
.Y(n_3514)
);

INVxp67_ASAP7_75t_L g3515 ( 
.A(n_3428),
.Y(n_3515)
);

AOI221xp5_ASAP7_75t_L g3516 ( 
.A1(n_3432),
.A2(n_427),
.B1(n_428),
.B2(n_429),
.C(n_430),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3433),
.B(n_429),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3395),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3435),
.B(n_3436),
.Y(n_3519)
);

NAND2xp5_ASAP7_75t_L g3520 ( 
.A(n_3438),
.B(n_430),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_3339),
.Y(n_3521)
);

INVx1_ASAP7_75t_SL g3522 ( 
.A(n_3308),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3361),
.Y(n_3523)
);

INVx1_ASAP7_75t_L g3524 ( 
.A(n_3373),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3380),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_3321),
.B(n_431),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_L g3527 ( 
.A(n_3359),
.B(n_431),
.Y(n_3527)
);

AOI21xp33_ASAP7_75t_L g3528 ( 
.A1(n_3345),
.A2(n_432),
.B(n_433),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3394),
.B(n_3326),
.Y(n_3529)
);

NOR2xp33_ASAP7_75t_L g3530 ( 
.A(n_3424),
.B(n_433),
.Y(n_3530)
);

INVx3_ASAP7_75t_L g3531 ( 
.A(n_3356),
.Y(n_3531)
);

AOI221xp5_ASAP7_75t_SL g3532 ( 
.A1(n_3304),
.A2(n_434),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3363),
.Y(n_3533)
);

INVx1_ASAP7_75t_SL g3534 ( 
.A(n_3384),
.Y(n_3534)
);

AND2x2_ASAP7_75t_L g3535 ( 
.A(n_3416),
.B(n_438),
.Y(n_3535)
);

NOR3x1_ASAP7_75t_L g3536 ( 
.A(n_3506),
.B(n_3442),
.C(n_3355),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3461),
.B(n_3293),
.Y(n_3537)
);

NOR2xp33_ASAP7_75t_L g3538 ( 
.A(n_3463),
.B(n_3370),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_SL g3539 ( 
.A(n_3465),
.B(n_3348),
.Y(n_3539)
);

NAND2x1_ASAP7_75t_L g3540 ( 
.A(n_3531),
.B(n_3365),
.Y(n_3540)
);

INVx2_ASAP7_75t_SL g3541 ( 
.A(n_3510),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_L g3542 ( 
.A(n_3465),
.B(n_3395),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3449),
.Y(n_3543)
);

O2A1O1Ixp33_ASAP7_75t_SL g3544 ( 
.A1(n_3479),
.A2(n_3306),
.B(n_3439),
.C(n_3367),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3454),
.Y(n_3545)
);

OAI211xp5_ASAP7_75t_SL g3546 ( 
.A1(n_3456),
.A2(n_3366),
.B(n_3368),
.C(n_3372),
.Y(n_3546)
);

BUFx6f_ASAP7_75t_L g3547 ( 
.A(n_3531),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_3535),
.Y(n_3548)
);

NOR3xp33_ASAP7_75t_L g3549 ( 
.A(n_3464),
.B(n_3362),
.C(n_3360),
.Y(n_3549)
);

NAND2xp5_ASAP7_75t_L g3550 ( 
.A(n_3459),
.B(n_3358),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3445),
.B(n_3470),
.Y(n_3551)
);

NOR2xp67_ASAP7_75t_SL g3552 ( 
.A(n_3533),
.B(n_3501),
.Y(n_3552)
);

NAND4xp25_ASAP7_75t_SL g3553 ( 
.A(n_3519),
.B(n_3407),
.C(n_3397),
.D(n_3385),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_3532),
.B(n_3312),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3466),
.B(n_3475),
.Y(n_3555)
);

O2A1O1Ixp33_ASAP7_75t_L g3556 ( 
.A1(n_3467),
.A2(n_3504),
.B(n_3498),
.C(n_3500),
.Y(n_3556)
);

NOR3x1_ASAP7_75t_L g3557 ( 
.A(n_3487),
.B(n_3377),
.C(n_3324),
.Y(n_3557)
);

INVx1_ASAP7_75t_L g3558 ( 
.A(n_3496),
.Y(n_3558)
);

NOR2xp33_ASAP7_75t_L g3559 ( 
.A(n_3455),
.B(n_3386),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3488),
.Y(n_3560)
);

INVx1_ASAP7_75t_L g3561 ( 
.A(n_3493),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_L g3562 ( 
.A(n_3534),
.B(n_3317),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3526),
.B(n_3381),
.Y(n_3563)
);

NOR3xp33_ASAP7_75t_L g3564 ( 
.A(n_3497),
.B(n_3328),
.C(n_3323),
.Y(n_3564)
);

AND2x2_ASAP7_75t_L g3565 ( 
.A(n_3446),
.B(n_3398),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3447),
.Y(n_3566)
);

OAI22xp5_ASAP7_75t_L g3567 ( 
.A1(n_3515),
.A2(n_3390),
.B1(n_3336),
.B2(n_3329),
.Y(n_3567)
);

AOI221xp5_ASAP7_75t_L g3568 ( 
.A1(n_3452),
.A2(n_3402),
.B1(n_3334),
.B2(n_3376),
.C(n_3375),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3489),
.B(n_3332),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3477),
.B(n_3333),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3533),
.B(n_3511),
.Y(n_3571)
);

AOI222xp33_ASAP7_75t_L g3572 ( 
.A1(n_3490),
.A2(n_3309),
.B1(n_3403),
.B2(n_3387),
.C1(n_3399),
.C2(n_3391),
.Y(n_3572)
);

INVx3_ASAP7_75t_L g3573 ( 
.A(n_3474),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_SL g3574 ( 
.A(n_3458),
.B(n_3369),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3478),
.B(n_3393),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_3505),
.Y(n_3576)
);

NOR3x1_ASAP7_75t_L g3577 ( 
.A(n_3509),
.B(n_3319),
.C(n_3318),
.Y(n_3577)
);

A2O1A1Ixp33_ASAP7_75t_SL g3578 ( 
.A1(n_3482),
.A2(n_3405),
.B(n_3379),
.C(n_3351),
.Y(n_3578)
);

AOI221x1_ASAP7_75t_L g3579 ( 
.A1(n_3517),
.A2(n_3441),
.B1(n_3388),
.B2(n_3389),
.C(n_3404),
.Y(n_3579)
);

NAND4xp25_ASAP7_75t_L g3580 ( 
.A(n_3529),
.B(n_3382),
.C(n_3303),
.D(n_3400),
.Y(n_3580)
);

AOI221x1_ASAP7_75t_L g3581 ( 
.A1(n_3520),
.A2(n_3301),
.B1(n_440),
.B2(n_441),
.C(n_442),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3457),
.B(n_439),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_SL g3583 ( 
.A(n_3476),
.B(n_441),
.Y(n_3583)
);

AOI21xp5_ASAP7_75t_L g3584 ( 
.A1(n_3450),
.A2(n_443),
.B(n_444),
.Y(n_3584)
);

AOI221x1_ASAP7_75t_L g3585 ( 
.A1(n_3484),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.C(n_448),
.Y(n_3585)
);

NAND3xp33_ASAP7_75t_L g3586 ( 
.A(n_3462),
.B(n_446),
.C(n_448),
.Y(n_3586)
);

NOR2xp33_ASAP7_75t_L g3587 ( 
.A(n_3469),
.B(n_3471),
.Y(n_3587)
);

NAND3xp33_ASAP7_75t_L g3588 ( 
.A(n_3502),
.B(n_449),
.C(n_450),
.Y(n_3588)
);

NOR2xp33_ASAP7_75t_L g3589 ( 
.A(n_3472),
.B(n_450),
.Y(n_3589)
);

OAI22xp33_ASAP7_75t_L g3590 ( 
.A1(n_3468),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3518),
.Y(n_3591)
);

NAND2xp5_ASAP7_75t_SL g3592 ( 
.A(n_3516),
.B(n_453),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_SL g3593 ( 
.A(n_3473),
.B(n_455),
.Y(n_3593)
);

NOR2xp33_ASAP7_75t_SL g3594 ( 
.A(n_3448),
.B(n_456),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_SL g3595 ( 
.A(n_3547),
.B(n_3508),
.Y(n_3595)
);

INVxp33_ASAP7_75t_L g3596 ( 
.A(n_3552),
.Y(n_3596)
);

OR2x2_ASAP7_75t_L g3597 ( 
.A(n_3541),
.B(n_3460),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_3547),
.B(n_3499),
.Y(n_3598)
);

OAI211xp5_ASAP7_75t_SL g3599 ( 
.A1(n_3543),
.A2(n_3513),
.B(n_3507),
.C(n_3503),
.Y(n_3599)
);

NOR2xp33_ASAP7_75t_SL g3600 ( 
.A(n_3537),
.B(n_3453),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_SL g3601 ( 
.A(n_3547),
.B(n_3492),
.Y(n_3601)
);

NOR3xp33_ASAP7_75t_L g3602 ( 
.A(n_3546),
.B(n_3527),
.C(n_3512),
.Y(n_3602)
);

NAND3x1_ASAP7_75t_L g3603 ( 
.A(n_3555),
.B(n_3481),
.C(n_3485),
.Y(n_3603)
);

OAI211xp5_ASAP7_75t_L g3604 ( 
.A1(n_3540),
.A2(n_3524),
.B(n_3525),
.C(n_3523),
.Y(n_3604)
);

NOR3xp33_ASAP7_75t_L g3605 ( 
.A(n_3553),
.B(n_3514),
.C(n_3521),
.Y(n_3605)
);

NAND2xp5_ASAP7_75t_SL g3606 ( 
.A(n_3573),
.B(n_3451),
.Y(n_3606)
);

OAI221xp5_ASAP7_75t_L g3607 ( 
.A1(n_3571),
.A2(n_3494),
.B1(n_3483),
.B2(n_3486),
.C(n_3495),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_3565),
.B(n_3522),
.Y(n_3608)
);

OAI21xp5_ASAP7_75t_L g3609 ( 
.A1(n_3556),
.A2(n_3491),
.B(n_3480),
.Y(n_3609)
);

OAI211xp5_ASAP7_75t_SL g3610 ( 
.A1(n_3551),
.A2(n_3568),
.B(n_3562),
.C(n_3544),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_3591),
.Y(n_3611)
);

AOI33xp33_ASAP7_75t_L g3612 ( 
.A1(n_3558),
.A2(n_3528),
.A3(n_3530),
.B1(n_459),
.B2(n_460),
.B3(n_461),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3585),
.B(n_457),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3573),
.A2(n_3554),
.B1(n_3587),
.B2(n_3550),
.Y(n_3614)
);

A2O1A1Ixp33_ASAP7_75t_L g3615 ( 
.A1(n_3538),
.A2(n_457),
.B(n_458),
.C(n_459),
.Y(n_3615)
);

AO21x1_ASAP7_75t_L g3616 ( 
.A1(n_3567),
.A2(n_3593),
.B(n_3583),
.Y(n_3616)
);

NOR3xp33_ASAP7_75t_L g3617 ( 
.A(n_3569),
.B(n_458),
.C(n_460),
.Y(n_3617)
);

NOR3xp33_ASAP7_75t_SL g3618 ( 
.A(n_3574),
.B(n_461),
.C(n_462),
.Y(n_3618)
);

NOR3x1_ASAP7_75t_L g3619 ( 
.A(n_3578),
.B(n_462),
.C(n_463),
.Y(n_3619)
);

NOR2xp33_ASAP7_75t_L g3620 ( 
.A(n_3542),
.B(n_463),
.Y(n_3620)
);

INVx1_ASAP7_75t_L g3621 ( 
.A(n_3545),
.Y(n_3621)
);

AOI211xp5_ASAP7_75t_SL g3622 ( 
.A1(n_3570),
.A2(n_3559),
.B(n_3575),
.C(n_3589),
.Y(n_3622)
);

NOR2xp67_ASAP7_75t_L g3623 ( 
.A(n_3584),
.B(n_465),
.Y(n_3623)
);

AND2x2_ASAP7_75t_L g3624 ( 
.A(n_3536),
.B(n_466),
.Y(n_3624)
);

AOI221xp5_ASAP7_75t_L g3625 ( 
.A1(n_3564),
.A2(n_466),
.B1(n_468),
.B2(n_469),
.C(n_471),
.Y(n_3625)
);

NAND4xp25_ASAP7_75t_L g3626 ( 
.A(n_3557),
.B(n_469),
.C(n_472),
.D(n_473),
.Y(n_3626)
);

OAI222xp33_ASAP7_75t_L g3627 ( 
.A1(n_3539),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.C1(n_475),
.C2(n_476),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_SL g3628 ( 
.A(n_3590),
.B(n_476),
.Y(n_3628)
);

INVxp67_ASAP7_75t_L g3629 ( 
.A(n_3563),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3548),
.B(n_477),
.Y(n_3630)
);

NAND4xp75_ASAP7_75t_L g3631 ( 
.A(n_3619),
.B(n_3577),
.C(n_3579),
.D(n_3581),
.Y(n_3631)
);

AO22x2_ASAP7_75t_L g3632 ( 
.A1(n_3614),
.A2(n_3588),
.B1(n_3576),
.B2(n_3560),
.Y(n_3632)
);

AOI21xp33_ASAP7_75t_SL g3633 ( 
.A1(n_3596),
.A2(n_3586),
.B(n_3582),
.Y(n_3633)
);

AOI221xp5_ASAP7_75t_L g3634 ( 
.A1(n_3611),
.A2(n_3549),
.B1(n_3566),
.B2(n_3561),
.C(n_3580),
.Y(n_3634)
);

AOI22xp5_ASAP7_75t_SL g3635 ( 
.A1(n_3629),
.A2(n_3594),
.B1(n_3592),
.B2(n_3572),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3608),
.Y(n_3636)
);

INVx1_ASAP7_75t_L g3637 ( 
.A(n_3613),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_SL g3638 ( 
.A(n_3627),
.B(n_477),
.Y(n_3638)
);

NAND4xp75_ASAP7_75t_L g3639 ( 
.A(n_3616),
.B(n_478),
.C(n_479),
.D(n_480),
.Y(n_3639)
);

OAI21xp5_ASAP7_75t_L g3640 ( 
.A1(n_3603),
.A2(n_479),
.B(n_481),
.Y(n_3640)
);

AND3x2_ASAP7_75t_L g3641 ( 
.A(n_3605),
.B(n_481),
.C(n_482),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3618),
.B(n_482),
.Y(n_3642)
);

NOR2x1_ASAP7_75t_L g3643 ( 
.A(n_3610),
.B(n_483),
.Y(n_3643)
);

AOI211xp5_ASAP7_75t_SL g3644 ( 
.A1(n_3604),
.A2(n_483),
.B(n_484),
.C(n_485),
.Y(n_3644)
);

INVx1_ASAP7_75t_L g3645 ( 
.A(n_3624),
.Y(n_3645)
);

INVx1_ASAP7_75t_SL g3646 ( 
.A(n_3597),
.Y(n_3646)
);

INVx1_ASAP7_75t_L g3647 ( 
.A(n_3612),
.Y(n_3647)
);

NAND3xp33_ASAP7_75t_L g3648 ( 
.A(n_3622),
.B(n_484),
.C(n_485),
.Y(n_3648)
);

AO22x2_ASAP7_75t_L g3649 ( 
.A1(n_3601),
.A2(n_486),
.B1(n_489),
.B2(n_490),
.Y(n_3649)
);

NAND4xp75_ASAP7_75t_L g3650 ( 
.A(n_3643),
.B(n_3609),
.C(n_3595),
.D(n_3598),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3641),
.B(n_3623),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_3646),
.B(n_3602),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_SL g3653 ( 
.A(n_3636),
.B(n_3621),
.Y(n_3653)
);

AOI22xp5_ASAP7_75t_L g3654 ( 
.A1(n_3645),
.A2(n_3606),
.B1(n_3600),
.B2(n_3599),
.Y(n_3654)
);

INVx2_ASAP7_75t_SL g3655 ( 
.A(n_3649),
.Y(n_3655)
);

INVx2_ASAP7_75t_L g3656 ( 
.A(n_3631),
.Y(n_3656)
);

AND2x2_ASAP7_75t_L g3657 ( 
.A(n_3644),
.B(n_3620),
.Y(n_3657)
);

AND3x4_ASAP7_75t_L g3658 ( 
.A(n_3635),
.B(n_3617),
.C(n_3607),
.Y(n_3658)
);

OR2x2_ASAP7_75t_L g3659 ( 
.A(n_3642),
.B(n_3626),
.Y(n_3659)
);

NOR2x1_ASAP7_75t_L g3660 ( 
.A(n_3648),
.B(n_3630),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3639),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_L g3662 ( 
.A(n_3637),
.B(n_3615),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3657),
.Y(n_3663)
);

OR2x2_ASAP7_75t_L g3664 ( 
.A(n_3656),
.B(n_3647),
.Y(n_3664)
);

CKINVDCx16_ASAP7_75t_R g3665 ( 
.A(n_3654),
.Y(n_3665)
);

NOR2xp33_ASAP7_75t_L g3666 ( 
.A(n_3651),
.B(n_3638),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3655),
.B(n_3632),
.Y(n_3667)
);

NOR2x1_ASAP7_75t_L g3668 ( 
.A(n_3658),
.B(n_3640),
.Y(n_3668)
);

NAND3xp33_ASAP7_75t_L g3669 ( 
.A(n_3652),
.B(n_3634),
.C(n_3633),
.Y(n_3669)
);

AOI221xp5_ASAP7_75t_L g3670 ( 
.A1(n_3653),
.A2(n_3628),
.B1(n_3625),
.B2(n_492),
.C(n_493),
.Y(n_3670)
);

AND2x4_ASAP7_75t_L g3671 ( 
.A(n_3661),
.B(n_486),
.Y(n_3671)
);

NOR3xp33_ASAP7_75t_L g3672 ( 
.A(n_3650),
.B(n_491),
.C(n_494),
.Y(n_3672)
);

OR2x2_ASAP7_75t_L g3673 ( 
.A(n_3665),
.B(n_3659),
.Y(n_3673)
);

AOI22xp5_ASAP7_75t_L g3674 ( 
.A1(n_3667),
.A2(n_3660),
.B1(n_3662),
.B2(n_495),
.Y(n_3674)
);

NOR2x1_ASAP7_75t_R g3675 ( 
.A(n_3663),
.B(n_491),
.Y(n_3675)
);

INVx2_ASAP7_75t_L g3676 ( 
.A(n_3668),
.Y(n_3676)
);

NAND4xp25_ASAP7_75t_L g3677 ( 
.A(n_3673),
.B(n_3669),
.C(n_3666),
.D(n_3664),
.Y(n_3677)
);

INVx2_ASAP7_75t_SL g3678 ( 
.A(n_3676),
.Y(n_3678)
);

BUFx2_ASAP7_75t_L g3679 ( 
.A(n_3675),
.Y(n_3679)
);

AOI22xp33_ASAP7_75t_L g3680 ( 
.A1(n_3678),
.A2(n_3672),
.B1(n_3670),
.B2(n_3674),
.Y(n_3680)
);

OAI211xp5_ASAP7_75t_SL g3681 ( 
.A1(n_3680),
.A2(n_3677),
.B(n_3679),
.C(n_3671),
.Y(n_3681)
);

INVx1_ASAP7_75t_L g3682 ( 
.A(n_3681),
.Y(n_3682)
);

OAI21xp5_ASAP7_75t_L g3683 ( 
.A1(n_3682),
.A2(n_494),
.B(n_496),
.Y(n_3683)
);

OAI22x1_ASAP7_75t_L g3684 ( 
.A1(n_3683),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_3684)
);

AO22x2_ASAP7_75t_L g3685 ( 
.A1(n_3684),
.A2(n_497),
.B1(n_498),
.B2(n_499),
.Y(n_3685)
);

OAI21xp33_ASAP7_75t_L g3686 ( 
.A1(n_3685),
.A2(n_500),
.B(n_501),
.Y(n_3686)
);

INVxp67_ASAP7_75t_SL g3687 ( 
.A(n_3686),
.Y(n_3687)
);

AND2x2_ASAP7_75t_L g3688 ( 
.A(n_3687),
.B(n_500),
.Y(n_3688)
);

AOI221xp5_ASAP7_75t_L g3689 ( 
.A1(n_3688),
.A2(n_501),
.B1(n_502),
.B2(n_504),
.C(n_505),
.Y(n_3689)
);

AOI211xp5_ASAP7_75t_L g3690 ( 
.A1(n_3689),
.A2(n_502),
.B(n_504),
.C(n_505),
.Y(n_3690)
);


endmodule