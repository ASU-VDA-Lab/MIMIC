module fake_ariane_1618_n_1886 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1886);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1886;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1654;
wire n_1560;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_590;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_16),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_139),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_24),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_10),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_36),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_75),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_108),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_141),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_43),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_40),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_18),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_81),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_2),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_54),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_103),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_158),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_44),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_123),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_65),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_22),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_0),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_38),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_62),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_91),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_150),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_22),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_92),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_34),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_72),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_153),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_100),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_50),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_51),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_16),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_55),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_171),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_96),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_20),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_127),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_152),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_174),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_47),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_97),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_49),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_163),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_111),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_166),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_32),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_105),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_42),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_20),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_119),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_15),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_25),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_175),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_66),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_129),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_84),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_124),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_90),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_40),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_101),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_39),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_118),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_167),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_126),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_143),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_146),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_19),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_74),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_79),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_60),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_106),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_19),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_42),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_149),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_55),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_115),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_78),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_93),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_68),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_107),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_50),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_133),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_56),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_1),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_63),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_109),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_140),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_62),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_8),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_44),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_121),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_87),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_64),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_27),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_98),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_104),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_54),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_138),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_85),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_24),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_35),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_110),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_82),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_38),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_73),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_33),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_48),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_43),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_131),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_170),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_89),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_157),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_45),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_102),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_48),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_8),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_28),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_137),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_31),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_2),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_4),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_134),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_160),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_34),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_12),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_169),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_159),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_52),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_113),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_86),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_70),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_125),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_122),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_162),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_39),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_83),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_9),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_112),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_46),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_148),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_3),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_14),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_145),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_31),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_7),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_250),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_195),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_288),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_195),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_330),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_195),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_R g363 ( 
.A(n_180),
.B(n_196),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_195),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_195),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_239),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_307),
.Y(n_367)
);

OR2x2_ASAP7_75t_L g368 ( 
.A(n_218),
.B(n_0),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_195),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_195),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_328),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_179),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_182),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_225),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_195),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_245),
.B(n_3),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_229),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_230),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_242),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_249),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_183),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_253),
.Y(n_382)
);

NOR2xp67_ASAP7_75t_L g383 ( 
.A(n_240),
.B(n_4),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_264),
.Y(n_384)
);

NAND2xp33_ASAP7_75t_R g385 ( 
.A(n_185),
.B(n_186),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_211),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_273),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_211),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g389 ( 
.A(n_240),
.B(n_5),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_269),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_211),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_252),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_276),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_189),
.B(n_5),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_211),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_211),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_296),
.B(n_7),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_290),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_290),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_279),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_179),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_290),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_191),
.B(n_10),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_184),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_290),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_281),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_247),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_326),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_247),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_192),
.B(n_11),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_290),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_285),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_207),
.B(n_11),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_296),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_301),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_301),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_291),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_317),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_317),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_297),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_303),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_273),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_306),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_273),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_247),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_310),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_335),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_356),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_208),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_193),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_184),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_332),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_183),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_274),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_197),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_332),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_274),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_274),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_213),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_220),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_227),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_197),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_209),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_362),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_401),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_358),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_360),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_217),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_360),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_381),
.B(n_231),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_357),
.Y(n_461)
);

OAI21x1_ASAP7_75t_L g462 ( 
.A1(n_365),
.A2(n_226),
.B(n_223),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_361),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_401),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_369),
.B(n_234),
.Y(n_466)
);

INVx6_ASAP7_75t_L g467 ( 
.A(n_389),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_370),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_370),
.B(n_238),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_375),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_373),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_386),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_388),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_376),
.B(n_268),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_368),
.A2(n_355),
.B1(n_214),
.B2(n_353),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_243),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_391),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_444),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_395),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_431),
.B(n_244),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_363),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_443),
.B(n_232),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_434),
.B(n_268),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_434),
.B(n_248),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_396),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_398),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_436),
.B(n_251),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_405),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_411),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_436),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_444),
.B(n_235),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_440),
.B(n_236),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_440),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_414),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_415),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_415),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_416),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_366),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_416),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_418),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_419),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_359),
.A2(n_181),
.B1(n_194),
.B2(n_300),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_422),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_394),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_426),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_426),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_429),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_429),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_430),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_430),
.Y(n_524)
);

INVx4_ASAP7_75t_L g525 ( 
.A(n_454),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_505),
.Y(n_526)
);

CKINVDCx6p67_ASAP7_75t_R g527 ( 
.A(n_461),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_458),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_482),
.B(n_387),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_467),
.B(n_368),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_458),
.Y(n_531)
);

INVxp33_ASAP7_75t_L g532 ( 
.A(n_451),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_505),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_458),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_472),
.Y(n_536)
);

AND2x6_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_489),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_517),
.B(n_377),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_387),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_482),
.B(n_404),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_467),
.A2(n_403),
.B1(n_410),
.B2(n_389),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_451),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_465),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_454),
.B(n_379),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_454),
.B(n_517),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_465),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_467),
.B(n_380),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_467),
.B(n_382),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_454),
.B(n_384),
.Y(n_549)
);

INVx6_ASAP7_75t_L g550 ( 
.A(n_454),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_464),
.B(n_407),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_467),
.A2(n_413),
.B1(n_383),
.B2(n_397),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_465),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_468),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_468),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_465),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_467),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_448),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_475),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_472),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_475),
.Y(n_561)
);

BUFx8_ASAP7_75t_SL g562 ( 
.A(n_509),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_448),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_482),
.B(n_467),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_448),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_486),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_475),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_476),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_462),
.A2(n_265),
.B(n_263),
.Y(n_571)
);

BUFx4f_ASAP7_75t_L g572 ( 
.A(n_505),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_476),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_479),
.B(n_385),
.C(n_390),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_463),
.B(n_393),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_476),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_495),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_463),
.B(n_400),
.Y(n_579)
);

CKINVDCx16_ASAP7_75t_R g580 ( 
.A(n_463),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_459),
.B(n_433),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_495),
.Y(n_582)
);

NAND3xp33_ASAP7_75t_L g583 ( 
.A(n_479),
.B(n_412),
.C(n_406),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_495),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_502),
.B(n_435),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_478),
.A2(n_446),
.B1(n_372),
.B2(n_437),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_502),
.B(n_439),
.Y(n_587)
);

BUFx4f_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_221),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_505),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_454),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_449),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_478),
.B(n_417),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_447),
.B(n_420),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_450),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_450),
.B(n_421),
.Y(n_597)
);

INVxp67_ASAP7_75t_SL g598 ( 
.A(n_468),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_447),
.B(n_424),
.Y(n_600)
);

BUFx3_ASAP7_75t_L g601 ( 
.A(n_452),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_452),
.B(n_428),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_489),
.B(n_432),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_452),
.B(n_409),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_453),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_489),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_489),
.A2(n_316),
.B1(n_254),
.B2(n_261),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_453),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_468),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_459),
.B(n_488),
.Y(n_610)
);

INVx4_ASAP7_75t_L g611 ( 
.A(n_468),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_453),
.B(n_427),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_449),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_456),
.B(n_442),
.Y(n_614)
);

INVxp67_ASAP7_75t_SL g615 ( 
.A(n_455),
.Y(n_615)
);

AND3x1_ASAP7_75t_L g616 ( 
.A(n_515),
.B(n_271),
.C(n_262),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_456),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_445),
.Y(n_618)
);

BUFx10_ASAP7_75t_L g619 ( 
.A(n_464),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_456),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_505),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_489),
.A2(n_515),
.B1(n_502),
.B2(n_501),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_492),
.A2(n_347),
.B1(n_325),
.B2(n_345),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_457),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_488),
.B(n_277),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_457),
.B(n_187),
.Y(n_626)
);

BUFx10_ASAP7_75t_L g627 ( 
.A(n_492),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_505),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_449),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_457),
.B(n_299),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_488),
.B(n_501),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_460),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_455),
.B(n_423),
.Y(n_634)
);

BUFx8_ASAP7_75t_SL g635 ( 
.A(n_501),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_460),
.B(n_185),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_507),
.B(n_287),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_449),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_449),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_460),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_470),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_507),
.B(n_292),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_470),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_471),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_505),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_471),
.Y(n_647)
);

CKINVDCx11_ASAP7_75t_R g648 ( 
.A(n_505),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_471),
.B(n_186),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_487),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_487),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_480),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_466),
.A2(n_334),
.B1(n_347),
.B2(n_214),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_481),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_511),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_480),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_481),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_500),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_R g661 ( 
.A(n_485),
.B(n_425),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_500),
.B(n_438),
.Y(n_662)
);

NOR2x1p5_ASAP7_75t_L g663 ( 
.A(n_507),
.B(n_198),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_466),
.A2(n_212),
.B1(n_355),
.B2(n_210),
.Y(n_664)
);

AND3x2_ASAP7_75t_L g665 ( 
.A(n_500),
.B(n_260),
.C(n_348),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_506),
.A2(n_309),
.B1(n_324),
.B2(n_295),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_491),
.Y(n_667)
);

AO22x2_ASAP7_75t_L g668 ( 
.A1(n_506),
.A2(n_272),
.B1(n_313),
.B2(n_329),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_507),
.B(n_322),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_481),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_491),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_493),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_493),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_469),
.B(n_507),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_503),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_469),
.B(n_188),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_481),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_660),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_668),
.A2(n_537),
.B1(n_622),
.B2(n_652),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_580),
.B(n_352),
.C(n_199),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_658),
.B(n_518),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_674),
.A2(n_462),
.B(n_485),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_569),
.B(n_441),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_558),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_650),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_558),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_634),
.B(n_539),
.Y(n_687)
);

AOI221xp5_ASAP7_75t_L g688 ( 
.A1(n_623),
.A2(n_338),
.B1(n_334),
.B2(n_331),
.C(n_325),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_563),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_595),
.B(n_600),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_658),
.B(n_615),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_564),
.B(n_518),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_564),
.B(n_518),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_660),
.B(n_462),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_563),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_631),
.B(n_518),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_597),
.B(n_518),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_532),
.B(n_367),
.Y(n_698)
);

BUFx5_ASAP7_75t_L g699 ( 
.A(n_537),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_530),
.B(n_490),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_651),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_667),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_671),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_660),
.B(n_462),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_537),
.A2(n_272),
.B1(n_188),
.B2(n_333),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_601),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_602),
.B(n_518),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_569),
.B(n_371),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_662),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_611),
.B(n_511),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_594),
.B(n_374),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_611),
.B(n_511),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_606),
.B(n_506),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_611),
.B(n_511),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_671),
.Y(n_717)
);

OAI221xp5_ASAP7_75t_L g718 ( 
.A1(n_541),
.A2(n_345),
.B1(n_350),
.B2(n_338),
.C(n_353),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_574),
.B(n_378),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_672),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_530),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_606),
.B(n_524),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_530),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_557),
.B(n_654),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_557),
.B(n_511),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_529),
.B(n_392),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_565),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_538),
.B(n_408),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_547),
.B(n_490),
.Y(n_729)
);

INVxp33_ASAP7_75t_L g730 ( 
.A(n_529),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_672),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_585),
.B(n_587),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_673),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_673),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_631),
.B(n_508),
.Y(n_735)
);

OR2x2_ASAP7_75t_SL g736 ( 
.A(n_583),
.B(n_494),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_575),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_548),
.B(n_494),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_614),
.B(n_198),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_604),
.B(n_508),
.Y(n_740)
);

INVxp67_ASAP7_75t_L g741 ( 
.A(n_551),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_567),
.B(n_199),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_612),
.B(n_626),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_630),
.B(n_524),
.Y(n_744)
);

BUFx5_ASAP7_75t_L g745 ( 
.A(n_537),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_551),
.B(n_201),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_537),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_654),
.B(n_511),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_601),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_544),
.B(n_524),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_575),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_549),
.B(n_508),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_585),
.B(n_512),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_530),
.A2(n_331),
.B1(n_205),
.B2(n_203),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_537),
.B(n_512),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_624),
.Y(n_756)
);

INVxp67_ASAP7_75t_L g757 ( 
.A(n_562),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_537),
.B(n_512),
.Y(n_758)
);

NAND2xp33_ASAP7_75t_L g759 ( 
.A(n_526),
.B(n_201),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_566),
.B(n_202),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_624),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_653),
.A2(n_212),
.B1(n_210),
.B2(n_205),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_642),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_526),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_587),
.B(n_513),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_542),
.B(n_527),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_663),
.A2(n_190),
.B1(n_200),
.B2(n_204),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_668),
.A2(n_523),
.B1(n_521),
.B2(n_513),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_528),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_654),
.B(n_511),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_523),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_528),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_576),
.B(n_202),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_566),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_535),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_554),
.B(n_511),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_581),
.B(n_523),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_535),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_581),
.B(n_610),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_546),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_579),
.B(n_203),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_642),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_603),
.B(n_315),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_619),
.B(n_315),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_610),
.A2(n_222),
.B1(n_190),
.B2(n_200),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_619),
.B(n_350),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_546),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_619),
.B(n_513),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_610),
.B(n_521),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_598),
.B(n_609),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_637),
.B(n_521),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_627),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_554),
.B(n_514),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_559),
.Y(n_794)
);

A2O1A1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_571),
.A2(n_503),
.B(n_510),
.C(n_519),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_540),
.B(n_504),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_559),
.Y(n_797)
);

AOI22xp33_ASAP7_75t_L g798 ( 
.A1(n_668),
.A2(n_520),
.B1(n_514),
.B2(n_516),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_540),
.B(n_504),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_637),
.B(n_503),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_536),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_627),
.B(n_504),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_554),
.B(n_514),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_555),
.B(n_514),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_553),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_643),
.B(n_503),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_676),
.B(n_504),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_668),
.A2(n_514),
.B1(n_520),
.B2(n_516),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_561),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_661),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_607),
.A2(n_514),
.B1(n_520),
.B2(n_516),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_643),
.B(n_510),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_618),
.B(n_510),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_552),
.A2(n_222),
.B1(n_354),
.B2(n_351),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_586),
.B(n_340),
.C(n_206),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_555),
.B(n_514),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_553),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_664),
.B(n_522),
.C(n_519),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_669),
.B(n_510),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_669),
.B(n_519),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_555),
.B(n_514),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_635),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_599),
.B(n_514),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_527),
.B(n_519),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_618),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_545),
.B(n_522),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_599),
.B(n_522),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_556),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_618),
.B(n_522),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_625),
.B(n_516),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_556),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_636),
.A2(n_219),
.B1(n_354),
.B2(n_351),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_599),
.B(n_516),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_561),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_625),
.B(n_666),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_536),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_649),
.B(n_516),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_L g839 ( 
.A1(n_589),
.A2(n_520),
.B1(n_516),
.B2(n_499),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_638),
.B(n_516),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_638),
.B(n_516),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_638),
.B(n_593),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_526),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_616),
.B(n_520),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_593),
.B(n_520),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_589),
.A2(n_520),
.B1(n_499),
.B2(n_498),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_596),
.A2(n_499),
.B(n_498),
.C(n_497),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_596),
.B(n_520),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_690),
.B(n_605),
.Y(n_849)
);

OAI321xp33_ASAP7_75t_L g850 ( 
.A1(n_711),
.A2(n_675),
.A3(n_570),
.B1(n_584),
.B2(n_582),
.C(n_578),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_687),
.B(n_605),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_732),
.B(n_617),
.C(n_608),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_694),
.A2(n_588),
.B(n_572),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_SL g854 ( 
.A1(n_678),
.A2(n_640),
.B(n_608),
.C(n_645),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_694),
.A2(n_588),
.B(n_572),
.Y(n_855)
);

OA22x2_ASAP7_75t_L g856 ( 
.A1(n_826),
.A2(n_665),
.B1(n_675),
.B2(n_560),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_743),
.B(n_617),
.Y(n_857)
);

BUFx8_ASAP7_75t_L g858 ( 
.A(n_710),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_691),
.B(n_620),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_706),
.A2(n_588),
.B(n_572),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_721),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_757),
.B(n_560),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_706),
.A2(n_632),
.B(n_620),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_750),
.A2(n_752),
.B(n_827),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_774),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_747),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_730),
.B(n_632),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_721),
.B(n_640),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_764),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_735),
.A2(n_644),
.B(n_641),
.C(n_645),
.Y(n_870)
);

OAI22xp5_ASAP7_75t_L g871 ( 
.A1(n_747),
.A2(n_644),
.B1(n_641),
.B2(n_647),
.Y(n_871)
);

INVx8_ASAP7_75t_L g872 ( 
.A(n_700),
.Y(n_872)
);

BUFx12f_ASAP7_75t_L g873 ( 
.A(n_774),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_730),
.B(n_525),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_791),
.A2(n_647),
.B(n_584),
.C(n_578),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_723),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_685),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_842),
.A2(n_591),
.B(n_525),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_800),
.A2(n_582),
.B(n_573),
.C(n_577),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_842),
.A2(n_591),
.B(n_525),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_729),
.B(n_531),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_698),
.B(n_713),
.Y(n_882)
);

CKINVDCx10_ASAP7_75t_R g883 ( 
.A(n_801),
.Y(n_883)
);

AND2x2_ASAP7_75t_SL g884 ( 
.A(n_679),
.B(n_270),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_712),
.A2(n_591),
.B(n_534),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_738),
.B(n_531),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_747),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_814),
.B(n_534),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_712),
.A2(n_543),
.B(n_656),
.Y(n_889)
);

INVxp67_ASAP7_75t_SL g890 ( 
.A(n_779),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_714),
.A2(n_543),
.B(n_656),
.Y(n_891)
);

INVx2_ASAP7_75t_SL g892 ( 
.A(n_766),
.Y(n_892)
);

CKINVDCx10_ASAP7_75t_R g893 ( 
.A(n_837),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_714),
.A2(n_657),
.B(n_656),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_716),
.A2(n_657),
.B(n_613),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_723),
.B(n_526),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_678),
.B(n_526),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_716),
.A2(n_657),
.B(n_613),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_788),
.B(n_568),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_840),
.A2(n_570),
.B(n_568),
.Y(n_900)
);

INVx3_ASAP7_75t_L g901 ( 
.A(n_708),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_753),
.B(n_592),
.Y(n_902)
);

A2O1A1Ixp33_ASAP7_75t_L g903 ( 
.A1(n_739),
.A2(n_573),
.B(n_577),
.C(n_629),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_719),
.B(n_741),
.Y(n_904)
);

CKINVDCx16_ASAP7_75t_R g905 ( 
.A(n_683),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_784),
.B(n_786),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_765),
.B(n_592),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_796),
.B(n_629),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_748),
.A2(n_633),
.B(n_639),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_748),
.A2(n_633),
.B(n_639),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_799),
.B(n_589),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_699),
.B(n_533),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_830),
.B(n_589),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_700),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_764),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_696),
.B(n_589),
.Y(n_916)
);

BUFx3_ASAP7_75t_L g917 ( 
.A(n_726),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_764),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_770),
.A2(n_628),
.B(n_590),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_770),
.A2(n_628),
.B(n_590),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_696),
.B(n_589),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_697),
.A2(n_628),
.B(n_590),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_708),
.A2(n_550),
.B1(n_533),
.B2(n_621),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_696),
.B(n_589),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_709),
.A2(n_628),
.B(n_590),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_838),
.A2(n_628),
.B(n_590),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_771),
.B(n_655),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_777),
.B(n_655),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_807),
.A2(n_813),
.B(n_821),
.C(n_820),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_840),
.A2(n_841),
.B(n_834),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_841),
.A2(n_646),
.B(n_621),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_828),
.A2(n_646),
.B(n_621),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_728),
.B(n_648),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_699),
.B(n_533),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_802),
.B(n_659),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_746),
.B(n_520),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_724),
.A2(n_646),
.B(n_621),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_742),
.B(n_659),
.Y(n_938)
);

AOI21xp33_ASAP7_75t_L g939 ( 
.A1(n_773),
.A2(n_677),
.B(n_670),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_760),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_708),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_740),
.B(n_670),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_684),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_789),
.A2(n_677),
.B(n_499),
.C(n_498),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_686),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_724),
.A2(n_646),
.B(n_621),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_790),
.A2(n_646),
.B(n_533),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_831),
.B(n_550),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_701),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_845),
.A2(n_533),
.B(n_550),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_848),
.A2(n_550),
.B(n_342),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_702),
.A2(n_319),
.B(n_343),
.C(n_280),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_744),
.A2(n_215),
.B(n_206),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_688),
.B(n_336),
.C(n_215),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_836),
.B(n_497),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_831),
.B(n_204),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_686),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_755),
.A2(n_216),
.B(n_219),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_758),
.A2(n_216),
.B(n_312),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_681),
.A2(n_312),
.B(n_314),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_776),
.A2(n_314),
.B(n_318),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_776),
.A2(n_318),
.B(n_321),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_760),
.Y(n_963)
);

OAI21xp5_ASAP7_75t_L g964 ( 
.A1(n_682),
.A2(n_498),
.B(n_497),
.Y(n_964)
);

NAND2xp33_ASAP7_75t_L g965 ( 
.A(n_699),
.B(n_745),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_793),
.A2(n_321),
.B(n_333),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_831),
.B(n_336),
.Y(n_967)
);

AOI21x1_ASAP7_75t_L g968 ( 
.A1(n_793),
.A2(n_497),
.B(n_473),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_692),
.B(n_339),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_693),
.B(n_339),
.Y(n_970)
);

BUFx3_ASAP7_75t_L g971 ( 
.A(n_792),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_803),
.A2(n_340),
.B(n_341),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_803),
.A2(n_341),
.B(n_342),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_804),
.B(n_283),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_718),
.A2(n_302),
.B(n_311),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_805),
.A2(n_822),
.B(n_817),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_699),
.B(n_224),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_700),
.B(n_473),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_805),
.A2(n_289),
.B(n_228),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_699),
.B(n_233),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_703),
.B(n_473),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_817),
.A2(n_293),
.B(n_246),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_822),
.A2(n_294),
.B(n_255),
.Y(n_983)
);

O2A1O1Ixp5_ASAP7_75t_L g984 ( 
.A1(n_725),
.A2(n_320),
.B(n_337),
.C(n_344),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_764),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_825),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_824),
.A2(n_286),
.B(n_237),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_843),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_699),
.B(n_241),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_689),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_SL g991 ( 
.A1(n_704),
.A2(n_346),
.B(n_349),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_792),
.B(n_256),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_794),
.A2(n_835),
.B1(n_797),
.B2(n_810),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_717),
.B(n_473),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_720),
.B(n_474),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_824),
.A2(n_284),
.B(n_259),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_731),
.A2(n_474),
.B(n_484),
.C(n_483),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_725),
.A2(n_298),
.B(n_266),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_798),
.A2(n_474),
.B1(n_484),
.B2(n_483),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_715),
.A2(n_304),
.B(n_267),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_733),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_734),
.A2(n_474),
.B(n_484),
.C(n_483),
.Y(n_1002)
);

AOI33xp33_ASAP7_75t_L g1003 ( 
.A1(n_762),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_17),
.B3(n_21),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_843),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_700),
.A2(n_305),
.B1(n_257),
.B2(n_258),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_795),
.A2(n_308),
.B(n_275),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_722),
.A2(n_496),
.B1(n_484),
.B2(n_483),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_749),
.B(n_278),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_781),
.B(n_282),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_756),
.A2(n_496),
.B1(n_484),
.B2(n_483),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_844),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_699),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_769),
.A2(n_484),
.B(n_483),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_769),
.A2(n_484),
.B(n_483),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_783),
.A2(n_496),
.B1(n_484),
.B2(n_483),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_761),
.B(n_13),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_763),
.B(n_782),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_843),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_833),
.B(n_815),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_768),
.B(n_17),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_811),
.B(n_496),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_772),
.A2(n_484),
.B(n_483),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_695),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_816),
.B(n_21),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_772),
.A2(n_496),
.B(n_477),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_808),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_745),
.B(n_496),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_795),
.A2(n_496),
.B(n_477),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_775),
.A2(n_780),
.B(n_787),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_775),
.Y(n_1030)
);

OA22x2_ASAP7_75t_L g1031 ( 
.A1(n_754),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_778),
.A2(n_477),
.B(n_496),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_707),
.A2(n_496),
.B1(n_477),
.B2(n_323),
.Y(n_1033)
);

OAI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_847),
.A2(n_477),
.B(n_323),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_695),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_819),
.B(n_23),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_785),
.B(n_26),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_778),
.A2(n_477),
.B(n_323),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_877),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_849),
.A2(n_759),
.B(n_843),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_917),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_906),
.B(n_767),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_869),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_SL g1044 ( 
.A1(n_884),
.A2(n_745),
.B1(n_759),
.B2(n_809),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_R g1045 ( 
.A(n_963),
.B(n_823),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_943),
.Y(n_1046)
);

INVxp67_ASAP7_75t_SL g1047 ( 
.A(n_890),
.Y(n_1047)
);

BUFx12f_ASAP7_75t_L g1048 ( 
.A(n_873),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_882),
.B(n_736),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_904),
.B(n_680),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_949),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_SL g1052 ( 
.A(n_862),
.B(n_933),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_864),
.A2(n_780),
.B(n_787),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_905),
.B(n_27),
.C(n_28),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_904),
.B(n_806),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_SL g1056 ( 
.A1(n_899),
.A2(n_806),
.B(n_818),
.C(n_832),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_945),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_899),
.A2(n_1009),
.B(n_1019),
.C(n_851),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_865),
.B(n_745),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_SL g1060 ( 
.A1(n_857),
.A2(n_832),
.B(n_829),
.C(n_818),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_986),
.B(n_829),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_872),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_940),
.B(n_745),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_1001),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_890),
.B(n_867),
.Y(n_1065)
);

AOI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_852),
.A2(n_745),
.B1(n_812),
.B2(n_839),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1036),
.A2(n_751),
.B(n_737),
.C(n_727),
.Y(n_1067)
);

OAI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_881),
.A2(n_727),
.B1(n_751),
.B2(n_737),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_884),
.A2(n_705),
.B1(n_745),
.B2(n_846),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_867),
.B(n_705),
.Y(n_1070)
);

NAND2x1p5_ASAP7_75t_L g1071 ( 
.A(n_866),
.B(n_477),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_1024),
.A2(n_1026),
.B(n_852),
.C(n_929),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_856),
.A2(n_975),
.B1(n_1011),
.B2(n_1020),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_957),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1026),
.B(n_29),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_886),
.A2(n_477),
.B1(n_323),
.B2(n_221),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1017),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1030),
.Y(n_1078)
);

NOR3xp33_ASAP7_75t_SL g1079 ( 
.A(n_993),
.B(n_29),
.C(n_30),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_986),
.B(n_30),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_929),
.A2(n_477),
.B(n_323),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_990),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_1023),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_859),
.A2(n_874),
.B1(n_902),
.B2(n_907),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_869),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_938),
.B(n_861),
.Y(n_1086)
);

BUFx12f_ASAP7_75t_L g1087 ( 
.A(n_858),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_SL g1088 ( 
.A(n_858),
.B(n_221),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_883),
.B(n_80),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_872),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_SL g1091 ( 
.A(n_892),
.B(n_221),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1035),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_R g1093 ( 
.A(n_893),
.B(n_77),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_861),
.B(n_33),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_955),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_876),
.B(n_992),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_863),
.A2(n_879),
.B(n_875),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_971),
.B(n_35),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_876),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_850),
.B(n_221),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1016),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1029),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_974),
.B(n_36),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_930),
.A2(n_37),
.B(n_41),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1005),
.B(n_37),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_908),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_888),
.B(n_41),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1021),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_969),
.B(n_45),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_981),
.Y(n_1110)
);

CKINVDCx16_ASAP7_75t_R g1111 ( 
.A(n_978),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_901),
.B(n_46),
.Y(n_1112)
);

OA22x2_ASAP7_75t_L g1113 ( 
.A1(n_1037),
.A2(n_914),
.B1(n_978),
.B2(n_956),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_869),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_970),
.B(n_51),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_942),
.B(n_53),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_978),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_914),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_856),
.Y(n_1119)
);

INVx1_ASAP7_75t_SL g1120 ( 
.A(n_1021),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_869),
.Y(n_1121)
);

AO221x2_ASAP7_75t_L g1122 ( 
.A1(n_991),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.C(n_61),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_872),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1031),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_1124)
);

NAND2x1p5_ASAP7_75t_L g1125 ( 
.A(n_866),
.B(n_887),
.Y(n_1125)
);

O2A1O1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_903),
.A2(n_61),
.B(n_63),
.C(n_67),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_916),
.B(n_921),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_901),
.B(n_69),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_954),
.B(n_88),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_994),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_948),
.A2(n_94),
.B1(n_95),
.B2(n_114),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_871),
.A2(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_900),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_936),
.B(n_130),
.Y(n_1134)
);

AND2x6_ASAP7_75t_L g1135 ( 
.A(n_887),
.B(n_915),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_941),
.B(n_135),
.Y(n_1136)
);

NAND2x1p5_ASAP7_75t_L g1137 ( 
.A(n_1004),
.B(n_161),
.Y(n_1137)
);

O2A1O1Ixp5_ASAP7_75t_L g1138 ( 
.A1(n_1028),
.A2(n_164),
.B(n_165),
.C(n_173),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1003),
.B(n_176),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_941),
.B(n_177),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_924),
.B(n_1004),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_915),
.B(n_918),
.Y(n_1142)
);

BUFx2_ASAP7_75t_SL g1143 ( 
.A(n_915),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_967),
.A2(n_870),
.B1(n_875),
.B2(n_879),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_870),
.A2(n_952),
.B(n_944),
.C(n_854),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_926),
.A2(n_922),
.B(n_925),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_913),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_853),
.A2(n_855),
.B(n_860),
.Y(n_1148)
);

AOI21x1_ASAP7_75t_L g1149 ( 
.A1(n_968),
.A2(n_964),
.B(n_947),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_995),
.Y(n_1150)
);

AND2x4_ASAP7_75t_L g1151 ( 
.A(n_915),
.B(n_918),
.Y(n_1151)
);

O2A1O1Ixp5_ASAP7_75t_L g1152 ( 
.A1(n_1034),
.A2(n_984),
.B(n_1006),
.C(n_897),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_911),
.A2(n_935),
.B1(n_927),
.B2(n_928),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_868),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_997),
.A2(n_1002),
.B(n_1038),
.Y(n_1155)
);

OAI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_923),
.A2(n_988),
.B1(n_918),
.B2(n_985),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_918),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_985),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_965),
.A2(n_932),
.B(n_950),
.Y(n_1159)
);

AO22x1_ASAP7_75t_L g1160 ( 
.A1(n_1031),
.A2(n_1008),
.B1(n_1018),
.B2(n_985),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_976),
.A2(n_889),
.B(n_891),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_919),
.A2(n_931),
.B(n_920),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_896),
.Y(n_1163)
);

OAI21xp33_ASAP7_75t_SL g1164 ( 
.A1(n_1012),
.A2(n_1027),
.B(n_912),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_985),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_944),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_894),
.A2(n_885),
.B(n_895),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_988),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_898),
.A2(n_909),
.B(n_910),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_937),
.A2(n_946),
.B(n_1013),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_988),
.B(n_1018),
.Y(n_1171)
);

BUFx12f_ASAP7_75t_L g1172 ( 
.A(n_988),
.Y(n_1172)
);

NAND3xp33_ASAP7_75t_SL g1173 ( 
.A(n_953),
.B(n_984),
.C(n_960),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_878),
.A2(n_880),
.B(n_951),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1010),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_1033),
.A2(n_1012),
.B1(n_961),
.B2(n_962),
.Y(n_1176)
);

O2A1O1Ixp33_ASAP7_75t_L g1177 ( 
.A1(n_939),
.A2(n_1007),
.B(n_1000),
.C(n_972),
.Y(n_1177)
);

NOR4xp25_ASAP7_75t_SL g1178 ( 
.A(n_977),
.B(n_989),
.C(n_980),
.D(n_934),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1018),
.B(n_966),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_973),
.B(n_999),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_958),
.A2(n_959),
.B(n_1018),
.Y(n_1181)
);

NOR3xp33_ASAP7_75t_SL g1182 ( 
.A(n_979),
.B(n_982),
.C(n_983),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_999),
.B(n_987),
.Y(n_1183)
);

O2A1O1Ixp33_ASAP7_75t_SL g1184 ( 
.A1(n_996),
.A2(n_998),
.B(n_1015),
.C(n_1014),
.Y(n_1184)
);

AOI221xp5_ASAP7_75t_L g1185 ( 
.A1(n_1032),
.A2(n_690),
.B1(n_906),
.B2(n_882),
.C(n_711),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1022),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1025),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_865),
.B(n_696),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_906),
.B(n_690),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_882),
.B(n_690),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_906),
.A2(n_690),
.B(n_687),
.C(n_882),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_882),
.B(n_732),
.Y(n_1192)
);

INVx8_ASAP7_75t_L g1193 ( 
.A(n_872),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_906),
.A2(n_690),
.B(n_687),
.C(n_882),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_906),
.B(n_690),
.Y(n_1195)
);

NOR4xp25_ASAP7_75t_L g1196 ( 
.A(n_906),
.B(n_690),
.C(n_1003),
.D(n_975),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_849),
.A2(n_690),
.B(n_864),
.Y(n_1197)
);

BUFx10_ASAP7_75t_L g1198 ( 
.A(n_1188),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_1191),
.Y(n_1199)
);

O2A1O1Ixp5_ASAP7_75t_L g1200 ( 
.A1(n_1194),
.A2(n_1195),
.B(n_1104),
.C(n_1197),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1047),
.A2(n_1081),
.B(n_1159),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1072),
.A2(n_1097),
.B(n_1081),
.Y(n_1202)
);

AOI221xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1185),
.A2(n_1103),
.B1(n_1144),
.B2(n_1126),
.C(n_1042),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1047),
.A2(n_1159),
.B(n_1097),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1152),
.A2(n_1100),
.B(n_1183),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1084),
.A2(n_1146),
.B(n_1148),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_1170),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_L g1208 ( 
.A1(n_1049),
.A2(n_1161),
.B(n_1152),
.C(n_1174),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1192),
.B(n_1055),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1146),
.A2(n_1162),
.B(n_1169),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1174),
.A2(n_1040),
.B(n_1167),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1039),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1185),
.A2(n_1129),
.B(n_1126),
.C(n_1115),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_SL g1214 ( 
.A(n_1088),
.B(n_1087),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1050),
.B(n_1052),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1040),
.A2(n_1153),
.B(n_1053),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1188),
.B(n_1099),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_1075),
.A2(n_1107),
.B(n_1128),
.C(n_1109),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1134),
.A2(n_1065),
.B(n_1184),
.Y(n_1219)
);

AOI221x1_ASAP7_75t_L g1220 ( 
.A1(n_1132),
.A2(n_1173),
.B1(n_1096),
.B2(n_1076),
.C(n_1181),
.Y(n_1220)
);

AOI221x1_ASAP7_75t_L g1221 ( 
.A1(n_1173),
.A2(n_1181),
.B1(n_1166),
.B2(n_1101),
.C(n_1116),
.Y(n_1221)
);

AOI21xp33_ASAP7_75t_L g1222 ( 
.A1(n_1113),
.A2(n_1073),
.B(n_1067),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1145),
.A2(n_1044),
.B(n_1105),
.C(n_1079),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1045),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1124),
.A2(n_1145),
.B1(n_1139),
.B2(n_1112),
.C(n_1080),
.Y(n_1225)
);

INVx5_ASAP7_75t_L g1226 ( 
.A(n_1135),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1048),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1156),
.A2(n_1060),
.B(n_1056),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1095),
.B(n_1077),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1062),
.B(n_1123),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1177),
.A2(n_1067),
.B(n_1136),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1051),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1064),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1175),
.A2(n_1196),
.B(n_1138),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1078),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1187),
.A2(n_1155),
.B(n_1138),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1041),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1186),
.A2(n_1176),
.B(n_1070),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1177),
.A2(n_1164),
.B(n_1140),
.Y(n_1239)
);

NAND2x1p5_ASAP7_75t_L g1240 ( 
.A(n_1062),
.B(n_1090),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1110),
.A2(n_1130),
.B(n_1179),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1125),
.A2(n_1178),
.B(n_1066),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1121),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1086),
.B(n_1106),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1155),
.A2(n_1137),
.B(n_1142),
.Y(n_1245)
);

BUFx10_ASAP7_75t_L g1246 ( 
.A(n_1098),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1044),
.A2(n_1079),
.B1(n_1094),
.B2(n_1098),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1172),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1137),
.A2(n_1125),
.B(n_1063),
.Y(n_1249)
);

AO21x2_ASAP7_75t_L g1250 ( 
.A1(n_1180),
.A2(n_1182),
.B(n_1147),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1069),
.A2(n_1150),
.B(n_1071),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_L g1252 ( 
.A(n_1099),
.B(n_1118),
.Y(n_1252)
);

BUFx12f_ASAP7_75t_L g1253 ( 
.A(n_1043),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1061),
.B(n_1111),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1069),
.A2(n_1071),
.B(n_1171),
.Y(n_1255)
);

BUFx3_ASAP7_75t_L g1256 ( 
.A(n_1193),
.Y(n_1256)
);

OAI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1054),
.A2(n_1154),
.B1(n_1163),
.B2(n_1091),
.C(n_1119),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1168),
.A2(n_1059),
.B(n_1113),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1193),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1182),
.A2(n_1147),
.B(n_1127),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1127),
.B(n_1141),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1168),
.A2(n_1165),
.B(n_1157),
.Y(n_1262)
);

AOI221x1_ASAP7_75t_L g1263 ( 
.A1(n_1131),
.A2(n_1108),
.B1(n_1092),
.B2(n_1082),
.C(n_1141),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1046),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1117),
.A2(n_1120),
.B1(n_1122),
.B2(n_1193),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1054),
.A2(n_1122),
.B1(n_1143),
.B2(n_1151),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1151),
.A2(n_1171),
.B(n_1160),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1043),
.A2(n_1158),
.B(n_1114),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1057),
.A2(n_1083),
.A3(n_1074),
.B1(n_1043),
.B2(n_1085),
.Y(n_1269)
);

OA21x2_ASAP7_75t_L g1270 ( 
.A1(n_1135),
.A2(n_1085),
.B(n_1114),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1158),
.B(n_1114),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1135),
.A2(n_1089),
.B(n_1093),
.Y(n_1272)
);

NOR2xp67_ASAP7_75t_L g1273 ( 
.A(n_1135),
.B(n_873),
.Y(n_1273)
);

AO32x2_ASAP7_75t_L g1274 ( 
.A1(n_1135),
.A2(n_1144),
.A3(n_1084),
.B1(n_1153),
.B2(n_1068),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_SL g1277 ( 
.A1(n_1058),
.A2(n_1047),
.B(n_1084),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1039),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_1087),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1096),
.B(n_873),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1039),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1192),
.B(n_905),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_L g1283 ( 
.A1(n_1190),
.A2(n_690),
.B(n_906),
.C(n_1191),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_SL g1284 ( 
.A(n_1058),
.B(n_1047),
.Y(n_1284)
);

AO21x1_ASAP7_75t_L g1285 ( 
.A1(n_1047),
.A2(n_690),
.B(n_906),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1144),
.A2(n_1084),
.A3(n_1153),
.B1(n_1068),
.B2(n_1156),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1041),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1039),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1188),
.Y(n_1295)
);

A2O1A1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1190),
.A2(n_690),
.B(n_906),
.C(n_882),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1297)
);

O2A1O1Ixp33_ASAP7_75t_SL g1298 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1058),
.C(n_690),
.Y(n_1298)
);

AOI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1190),
.A2(n_690),
.B1(n_906),
.B2(n_882),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1041),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_1159),
.Y(n_1301)
);

AND2x2_ASAP7_75t_SL g1302 ( 
.A(n_1111),
.B(n_884),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1081),
.A2(n_1148),
.B(n_1146),
.Y(n_1305)
);

CKINVDCx20_ASAP7_75t_R g1306 ( 
.A(n_1089),
.Y(n_1306)
);

AOI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1081),
.A2(n_1149),
.B(n_1148),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1190),
.B(n_1189),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_1159),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_1159),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1039),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1039),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1191),
.A2(n_1194),
.B1(n_1190),
.B2(n_1058),
.C(n_1189),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1089),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1058),
.A2(n_1194),
.B(n_1191),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1039),
.Y(n_1319)
);

O2A1O1Ixp33_ASAP7_75t_SL g1320 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1058),
.C(n_690),
.Y(n_1320)
);

AO22x2_ASAP7_75t_L g1321 ( 
.A1(n_1047),
.A2(n_1144),
.B1(n_1065),
.B2(n_1101),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_1048),
.Y(n_1322)
);

AOI21xp33_ASAP7_75t_L g1323 ( 
.A1(n_1190),
.A2(n_690),
.B(n_906),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1121),
.Y(n_1324)
);

CKINVDCx16_ASAP7_75t_R g1325 ( 
.A(n_1087),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1190),
.A2(n_690),
.B(n_906),
.C(n_882),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1089),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1099),
.Y(n_1328)
);

INVxp67_ASAP7_75t_L g1329 ( 
.A(n_1041),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_1087),
.Y(n_1331)
);

BUFx2_ASAP7_75t_L g1332 ( 
.A(n_1188),
.Y(n_1332)
);

OAI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1058),
.A2(n_1194),
.B(n_1191),
.Y(n_1333)
);

AOI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1081),
.A2(n_1149),
.B(n_1148),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1062),
.B(n_1188),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1190),
.C(n_690),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1197),
.A2(n_1058),
.B(n_864),
.Y(n_1337)
);

OA21x2_ASAP7_75t_L g1338 ( 
.A1(n_1081),
.A2(n_1148),
.B(n_1146),
.Y(n_1338)
);

O2A1O1Ixp33_ASAP7_75t_SL g1339 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1058),
.C(n_690),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1039),
.Y(n_1340)
);

O2A1O1Ixp33_ASAP7_75t_L g1341 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1190),
.C(n_690),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1188),
.Y(n_1342)
);

BUFx8_ASAP7_75t_SL g1343 ( 
.A(n_1087),
.Y(n_1343)
);

O2A1O1Ixp33_ASAP7_75t_SL g1344 ( 
.A1(n_1191),
.A2(n_1194),
.B(n_1058),
.C(n_690),
.Y(n_1344)
);

AOI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1189),
.A2(n_1195),
.B(n_1103),
.Y(n_1345)
);

NAND3xp33_ASAP7_75t_SL g1346 ( 
.A(n_1190),
.B(n_1194),
.C(n_1191),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1062),
.B(n_1188),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1058),
.A2(n_1194),
.B(n_1191),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1081),
.A2(n_1102),
.A3(n_1133),
.B(n_1146),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1149),
.A2(n_1148),
.B(n_1159),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1212),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1250),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1302),
.A2(n_1346),
.B1(n_1299),
.B2(n_1247),
.Y(n_1353)
);

BUFx10_ASAP7_75t_L g1354 ( 
.A(n_1224),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1248),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1299),
.A2(n_1326),
.B1(n_1296),
.B2(n_1323),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1237),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1247),
.A2(n_1265),
.B1(n_1215),
.B2(n_1317),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1343),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1232),
.Y(n_1360)
);

INVx6_ASAP7_75t_L g1361 ( 
.A(n_1198),
.Y(n_1361)
);

INVx3_ASAP7_75t_SL g1362 ( 
.A(n_1279),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1226),
.Y(n_1363)
);

CKINVDCx11_ASAP7_75t_R g1364 ( 
.A(n_1325),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1237),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1331),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1284),
.A2(n_1321),
.B1(n_1348),
.B2(n_1333),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1336),
.A2(n_1341),
.B1(n_1333),
.B2(n_1317),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1233),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1348),
.A2(n_1222),
.B1(n_1284),
.B2(n_1209),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_1306),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1321),
.A2(n_1257),
.B1(n_1310),
.B2(n_1282),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1202),
.A2(n_1254),
.B1(n_1285),
.B2(n_1244),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1213),
.A2(n_1223),
.B1(n_1277),
.B2(n_1199),
.Y(n_1374)
);

INVx6_ASAP7_75t_L g1375 ( 
.A(n_1198),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1300),
.A2(n_1329),
.B1(n_1202),
.B2(n_1252),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1229),
.A2(n_1314),
.B1(n_1293),
.B2(n_1319),
.Y(n_1377)
);

INVx3_ASAP7_75t_L g1378 ( 
.A(n_1253),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1217),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1278),
.Y(n_1380)
);

INVxp67_ASAP7_75t_SL g1381 ( 
.A(n_1204),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1227),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1290),
.Y(n_1383)
);

BUFx12f_ASAP7_75t_L g1384 ( 
.A(n_1324),
.Y(n_1384)
);

OAI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1214),
.A2(n_1266),
.B1(n_1290),
.B2(n_1313),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_SL g1386 ( 
.A1(n_1214),
.A2(n_1266),
.B1(n_1205),
.B2(n_1225),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_SL g1387 ( 
.A1(n_1205),
.A2(n_1225),
.B1(n_1203),
.B2(n_1239),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1203),
.A2(n_1242),
.B1(n_1250),
.B2(n_1340),
.Y(n_1388)
);

BUFx8_ASAP7_75t_L g1389 ( 
.A(n_1243),
.Y(n_1389)
);

CKINVDCx11_ASAP7_75t_R g1390 ( 
.A(n_1316),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1281),
.A2(n_1235),
.B1(n_1264),
.B2(n_1261),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1315),
.B(n_1328),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1260),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1270),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1234),
.A2(n_1260),
.B1(n_1315),
.B2(n_1246),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1324),
.Y(n_1396)
);

INVx6_ASAP7_75t_L g1397 ( 
.A(n_1335),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1241),
.A2(n_1280),
.B1(n_1234),
.B2(n_1342),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1259),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1238),
.A2(n_1251),
.B1(n_1272),
.B2(n_1274),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1269),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1269),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1295),
.B(n_1332),
.Y(n_1404)
);

BUFx3_ASAP7_75t_L g1405 ( 
.A(n_1256),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1327),
.Y(n_1406)
);

CKINVDCx11_ASAP7_75t_R g1407 ( 
.A(n_1322),
.Y(n_1407)
);

INVx2_ASAP7_75t_R g1408 ( 
.A(n_1208),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1262),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1258),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1298),
.B(n_1320),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_SL g1412 ( 
.A1(n_1238),
.A2(n_1274),
.B1(n_1255),
.B2(n_1286),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1274),
.A2(n_1286),
.B1(n_1275),
.B2(n_1288),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1230),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1339),
.B(n_1344),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1289),
.A2(n_1337),
.B1(n_1292),
.B2(n_1294),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1230),
.B(n_1347),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1335),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1271),
.Y(n_1419)
);

BUFx8_ASAP7_75t_SL g1420 ( 
.A(n_1259),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1291),
.A2(n_1304),
.B1(n_1330),
.B2(n_1318),
.Y(n_1421)
);

BUFx2_ASAP7_75t_L g1422 ( 
.A(n_1347),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1240),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1276),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1286),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1308),
.A2(n_1231),
.B1(n_1219),
.B2(n_1273),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1268),
.Y(n_1427)
);

CKINVDCx11_ASAP7_75t_R g1428 ( 
.A(n_1345),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1276),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1240),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1270),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1283),
.A2(n_1206),
.B1(n_1201),
.B2(n_1216),
.Y(n_1432)
);

CKINVDCx6p67_ASAP7_75t_R g1433 ( 
.A(n_1218),
.Y(n_1433)
);

BUFx4f_ASAP7_75t_SL g1434 ( 
.A(n_1221),
.Y(n_1434)
);

CKINVDCx20_ASAP7_75t_R g1435 ( 
.A(n_1267),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1287),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1200),
.B(n_1249),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1297),
.B(n_1303),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1305),
.A2(n_1338),
.B1(n_1228),
.B2(n_1211),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1297),
.Y(n_1440)
);

INVx3_ASAP7_75t_L g1441 ( 
.A(n_1245),
.Y(n_1441)
);

BUFx12f_ASAP7_75t_L g1442 ( 
.A(n_1263),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1303),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1220),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1309),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1305),
.A2(n_1338),
.B1(n_1210),
.B2(n_1236),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1210),
.A2(n_1312),
.B1(n_1350),
.B2(n_1301),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1349),
.B(n_1311),
.Y(n_1448)
);

BUFx6f_ASAP7_75t_SL g1449 ( 
.A(n_1349),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1334),
.A2(n_1299),
.B1(n_1190),
.B2(n_1296),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1307),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1207),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1212),
.Y(n_1453)
);

NAND2x1p5_ASAP7_75t_L g1454 ( 
.A(n_1226),
.B(n_1270),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1299),
.A2(n_1190),
.B1(n_1326),
.B2(n_1296),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1302),
.A2(n_884),
.B1(n_690),
.B2(n_1190),
.Y(n_1456)
);

BUFx4f_ASAP7_75t_SL g1457 ( 
.A(n_1306),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1302),
.A2(n_884),
.B1(n_1122),
.B2(n_690),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1302),
.A2(n_884),
.B1(n_690),
.B2(n_1190),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1302),
.A2(n_884),
.B1(n_690),
.B2(n_1190),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1299),
.A2(n_1284),
.B1(n_1189),
.B2(n_1195),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1302),
.A2(n_884),
.B1(n_690),
.B2(n_1190),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1248),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1343),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1198),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1212),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1299),
.A2(n_1190),
.B1(n_1326),
.B2(n_1296),
.Y(n_1467)
);

BUFx8_ASAP7_75t_L g1468 ( 
.A(n_1243),
.Y(n_1468)
);

INVx5_ASAP7_75t_L g1469 ( 
.A(n_1226),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1212),
.Y(n_1470)
);

CKINVDCx11_ASAP7_75t_R g1471 ( 
.A(n_1325),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1410),
.Y(n_1472)
);

AOI21xp33_ASAP7_75t_L g1473 ( 
.A1(n_1461),
.A2(n_1374),
.B(n_1456),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1359),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1437),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1432),
.A2(n_1439),
.B(n_1446),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1357),
.B(n_1365),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1376),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1424),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1429),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1379),
.B(n_1401),
.Y(n_1481)
);

OA21x2_ASAP7_75t_L g1482 ( 
.A1(n_1439),
.A2(n_1446),
.B(n_1421),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1431),
.B(n_1469),
.Y(n_1483)
);

AOI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1451),
.A2(n_1450),
.B(n_1448),
.Y(n_1484)
);

AOI21xp5_ASAP7_75t_SL g1485 ( 
.A1(n_1461),
.A2(n_1368),
.B(n_1385),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1416),
.A2(n_1421),
.B(n_1426),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1436),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1443),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1445),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1469),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1367),
.B(n_1412),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1409),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1440),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1455),
.A2(n_1467),
.B(n_1356),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1438),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1418),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1497)
);

CKINVDCx16_ASAP7_75t_R g1498 ( 
.A(n_1384),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1416),
.A2(n_1426),
.B(n_1441),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1351),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1431),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1367),
.A2(n_1381),
.B(n_1413),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1360),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1394),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1369),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1392),
.B(n_1352),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1364),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1394),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1381),
.A2(n_1413),
.B(n_1411),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1352),
.A2(n_1452),
.B(n_1393),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1380),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1444),
.Y(n_1512)
);

OAI21x1_ASAP7_75t_L g1513 ( 
.A1(n_1415),
.A2(n_1454),
.B(n_1398),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1453),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1383),
.Y(n_1515)
);

INVx3_ASAP7_75t_SL g1516 ( 
.A(n_1433),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1466),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1412),
.B(n_1470),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1449),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1425),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1373),
.B(n_1393),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1373),
.B(n_1387),
.Y(n_1522)
);

INVx3_ASAP7_75t_L g1523 ( 
.A(n_1434),
.Y(n_1523)
);

BUFx2_ASAP7_75t_L g1524 ( 
.A(n_1434),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1377),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1377),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1366),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1419),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1388),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1456),
.A2(n_1462),
.B(n_1460),
.C(n_1459),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1388),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1387),
.A2(n_1353),
.B(n_1386),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1353),
.B(n_1358),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1358),
.B(n_1372),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1370),
.B(n_1408),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1442),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1370),
.B(n_1408),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1400),
.A2(n_1404),
.B(n_1447),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1400),
.B(n_1395),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1391),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_SL g1541 ( 
.A(n_1389),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1427),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1391),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1447),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1395),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1458),
.B(n_1372),
.Y(n_1546)
);

AO31x2_ASAP7_75t_L g1547 ( 
.A1(n_1430),
.A2(n_1422),
.A3(n_1414),
.B(n_1417),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1398),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1423),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1363),
.B(n_1399),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1464),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1435),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1397),
.B(n_1399),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1428),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1361),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1516),
.B(n_1362),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1524),
.B(n_1405),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1524),
.B(n_1405),
.Y(n_1558)
);

OR2x2_ASAP7_75t_SL g1559 ( 
.A(n_1554),
.B(n_1396),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1552),
.B(n_1355),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1552),
.B(n_1463),
.Y(n_1561)
);

OAI211xp5_ASAP7_75t_L g1562 ( 
.A1(n_1494),
.A2(n_1471),
.B(n_1407),
.C(n_1390),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1481),
.B(n_1362),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1516),
.B(n_1457),
.Y(n_1564)
);

AO32x2_ASAP7_75t_L g1565 ( 
.A1(n_1478),
.A2(n_1389),
.A3(n_1468),
.B1(n_1420),
.B2(n_1375),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1515),
.B(n_1378),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_SL g1567 ( 
.A1(n_1530),
.A2(n_1468),
.B(n_1354),
.Y(n_1567)
);

INVxp67_ASAP7_75t_L g1568 ( 
.A(n_1477),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1515),
.B(n_1378),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1516),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1473),
.A2(n_1371),
.B(n_1406),
.C(n_1457),
.Y(n_1571)
);

OAI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1485),
.A2(n_1354),
.B(n_1361),
.Y(n_1572)
);

NOR2x1_ASAP7_75t_L g1573 ( 
.A(n_1554),
.B(n_1382),
.Y(n_1573)
);

AO32x2_ASAP7_75t_L g1574 ( 
.A1(n_1518),
.A2(n_1375),
.A3(n_1465),
.B1(n_1475),
.B2(n_1506),
.Y(n_1574)
);

AND2x6_ASAP7_75t_L g1575 ( 
.A(n_1539),
.B(n_1465),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1532),
.A2(n_1533),
.B1(n_1545),
.B2(n_1522),
.Y(n_1576)
);

AO32x2_ASAP7_75t_L g1577 ( 
.A1(n_1518),
.A2(n_1475),
.A3(n_1506),
.B1(n_1491),
.B2(n_1497),
.Y(n_1577)
);

OAI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1545),
.A2(n_1485),
.B1(n_1534),
.B2(n_1523),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1528),
.B(n_1542),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1500),
.Y(n_1580)
);

AOI221xp5_ASAP7_75t_L g1581 ( 
.A1(n_1546),
.A2(n_1521),
.B1(n_1539),
.B2(n_1502),
.C(n_1529),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1500),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1483),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1498),
.B(n_1507),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1483),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1523),
.B(n_1520),
.Y(n_1586)
);

OA21x2_ASAP7_75t_L g1587 ( 
.A1(n_1476),
.A2(n_1509),
.B(n_1499),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1503),
.Y(n_1588)
);

AND2x4_ASAP7_75t_L g1589 ( 
.A(n_1547),
.B(n_1483),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1536),
.B(n_1512),
.Y(n_1590)
);

CKINVDCx14_ASAP7_75t_R g1591 ( 
.A(n_1474),
.Y(n_1591)
);

OA21x2_ASAP7_75t_L g1592 ( 
.A1(n_1476),
.A2(n_1499),
.B(n_1544),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_SL g1593 ( 
.A1(n_1551),
.A2(n_1541),
.B(n_1512),
.C(n_1534),
.Y(n_1593)
);

CKINVDCx20_ASAP7_75t_R g1594 ( 
.A(n_1527),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1536),
.B(n_1512),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1486),
.A2(n_1535),
.B(n_1537),
.Y(n_1596)
);

INVx4_ASAP7_75t_L g1597 ( 
.A(n_1550),
.Y(n_1597)
);

AO32x2_ASAP7_75t_L g1598 ( 
.A1(n_1491),
.A2(n_1497),
.A3(n_1495),
.B1(n_1547),
.B2(n_1521),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1505),
.B(n_1511),
.Y(n_1599)
);

O2A1O1Ixp33_ASAP7_75t_SL g1600 ( 
.A1(n_1512),
.A2(n_1555),
.B(n_1542),
.C(n_1544),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1511),
.B(n_1514),
.Y(n_1601)
);

BUFx8_ASAP7_75t_L g1602 ( 
.A(n_1549),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1546),
.A2(n_1529),
.B1(n_1531),
.B2(n_1537),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1498),
.B(n_1496),
.Y(n_1604)
);

A2O1A1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1531),
.A2(n_1535),
.B(n_1548),
.C(n_1543),
.Y(n_1605)
);

OAI211xp5_ASAP7_75t_L g1606 ( 
.A1(n_1548),
.A2(n_1486),
.B(n_1482),
.C(n_1526),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1514),
.Y(n_1607)
);

BUFx8_ASAP7_75t_SL g1608 ( 
.A(n_1553),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1517),
.B(n_1525),
.Y(n_1609)
);

OAI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1578),
.A2(n_1513),
.B(n_1540),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1577),
.B(n_1482),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1583),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1582),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1510),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1577),
.B(n_1482),
.Y(n_1615)
);

INVx1_ASAP7_75t_SL g1616 ( 
.A(n_1563),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1577),
.B(n_1482),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1574),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1574),
.B(n_1501),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1510),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1581),
.A2(n_1538),
.B1(n_1517),
.B2(n_1519),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1574),
.B(n_1501),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1607),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1501),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1587),
.B(n_1484),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_1597),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1580),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1599),
.B(n_1538),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1576),
.A2(n_1603),
.B1(n_1575),
.B2(n_1538),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1601),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1609),
.B(n_1493),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1592),
.B(n_1493),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1598),
.B(n_1484),
.Y(n_1634)
);

AOI222xp33_ASAP7_75t_L g1635 ( 
.A1(n_1605),
.A2(n_1488),
.B1(n_1489),
.B2(n_1487),
.C1(n_1479),
.C2(n_1480),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_1472),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1592),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1602),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1598),
.B(n_1472),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1632),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1624),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1620),
.B(n_1596),
.Y(n_1644)
);

AOI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1622),
.A2(n_1630),
.B1(n_1611),
.B2(n_1615),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1636),
.B(n_1606),
.Y(n_1646)
);

NAND5xp2_ASAP7_75t_SL g1647 ( 
.A(n_1622),
.B(n_1562),
.C(n_1572),
.D(n_1571),
.E(n_1557),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1624),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1633),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1613),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1633),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1633),
.Y(n_1652)
);

AOI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1619),
.A2(n_1593),
.B1(n_1568),
.B2(n_1600),
.C(n_1567),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1632),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1617),
.Y(n_1655)
);

OAI211xp5_ASAP7_75t_L g1656 ( 
.A1(n_1630),
.A2(n_1591),
.B(n_1570),
.C(n_1566),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1620),
.B(n_1585),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1620),
.B(n_1585),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1628),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1623),
.B(n_1589),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1635),
.A2(n_1575),
.B1(n_1610),
.B2(n_1618),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1616),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1617),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1556),
.C(n_1564),
.D(n_1584),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1640),
.B(n_1492),
.Y(n_1667)
);

AOI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1610),
.A2(n_1611),
.B1(n_1615),
.B2(n_1618),
.C1(n_1634),
.C2(n_1575),
.Y(n_1668)
);

OAI211xp5_ASAP7_75t_L g1669 ( 
.A1(n_1619),
.A2(n_1569),
.B(n_1558),
.C(n_1573),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1639),
.A2(n_1559),
.B1(n_1565),
.B2(n_1594),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1640),
.B(n_1492),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1623),
.B(n_1586),
.Y(n_1672)
);

OAI31xp33_ASAP7_75t_SL g1673 ( 
.A1(n_1615),
.A2(n_1595),
.A3(n_1590),
.B(n_1565),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1612),
.Y(n_1674)
);

AO21x2_ASAP7_75t_L g1675 ( 
.A1(n_1638),
.A2(n_1504),
.B(n_1508),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1646),
.B(n_1621),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1644),
.B(n_1640),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1644),
.B(n_1618),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1634),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1661),
.Y(n_1680)
);

NOR2x1_ASAP7_75t_L g1681 ( 
.A(n_1666),
.B(n_1639),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1660),
.B(n_1634),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1674),
.B(n_1625),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1675),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1675),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1655),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1657),
.B(n_1625),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1658),
.B(n_1637),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_SL g1689 ( 
.A(n_1653),
.Y(n_1689)
);

NAND2x1p5_ASAP7_75t_L g1690 ( 
.A(n_1663),
.B(n_1626),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1641),
.B(n_1642),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1675),
.Y(n_1692)
);

AO21x1_ASAP7_75t_SL g1693 ( 
.A1(n_1646),
.A2(n_1614),
.B(n_1631),
.Y(n_1693)
);

AND2x4_ASAP7_75t_L g1694 ( 
.A(n_1674),
.B(n_1627),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1675),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1649),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1673),
.B(n_1626),
.C(n_1614),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.B(n_1662),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_L g1699 ( 
.A(n_1669),
.B(n_1638),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1654),
.B(n_1631),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1643),
.B(n_1631),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1649),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1643),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1650),
.Y(n_1704)
);

HB1xp67_ASAP7_75t_L g1705 ( 
.A(n_1648),
.Y(n_1705)
);

INVxp67_ASAP7_75t_SL g1706 ( 
.A(n_1649),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1648),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1651),
.Y(n_1708)
);

OAI31xp33_ASAP7_75t_L g1709 ( 
.A1(n_1690),
.A2(n_1697),
.A3(n_1656),
.B(n_1669),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1703),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1679),
.B(n_1664),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1667),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1703),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1698),
.B(n_1673),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1705),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1705),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1707),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1698),
.B(n_1672),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1689),
.Y(n_1719)
);

NOR2x1_ASAP7_75t_L g1720 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1720)
);

NAND2x1p5_ASAP7_75t_L g1721 ( 
.A(n_1681),
.B(n_1663),
.Y(n_1721)
);

OR2x6_ASAP7_75t_L g1722 ( 
.A(n_1690),
.B(n_1670),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1698),
.B(n_1672),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1707),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1687),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1701),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1701),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1700),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1687),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1679),
.B(n_1664),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1681),
.B(n_1670),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1676),
.B(n_1667),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1700),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1689),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1679),
.B(n_1671),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1680),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1680),
.Y(n_1737)
);

INVxp67_ASAP7_75t_L g1738 ( 
.A(n_1693),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

AOI221xp5_ASAP7_75t_L g1740 ( 
.A1(n_1697),
.A2(n_1647),
.B1(n_1645),
.B2(n_1656),
.C(n_1652),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1691),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1687),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1687),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1698),
.B(n_1672),
.Y(n_1744)
);

NAND2x1p5_ASAP7_75t_L g1745 ( 
.A(n_1686),
.B(n_1655),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1676),
.B(n_1671),
.Y(n_1746)
);

AND2x2_ASAP7_75t_SL g1747 ( 
.A(n_1686),
.B(n_1653),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1704),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1677),
.B(n_1662),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1682),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1677),
.B(n_1659),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1710),
.Y(n_1752)
);

INVxp67_ASAP7_75t_SL g1753 ( 
.A(n_1721),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1725),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

AND3x1_ASAP7_75t_L g1756 ( 
.A(n_1709),
.B(n_1679),
.C(n_1647),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1739),
.B(n_1741),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1608),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.B(n_1677),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_SL g1761 ( 
.A(n_1720),
.B(n_1699),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1678),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1734),
.Y(n_1763)
);

XNOR2xp5_ASAP7_75t_L g1764 ( 
.A(n_1747),
.B(n_1690),
.Y(n_1764)
);

O2A1O1Ixp33_ASAP7_75t_L g1765 ( 
.A1(n_1731),
.A2(n_1690),
.B(n_1699),
.C(n_1668),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1712),
.B(n_1678),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1749),
.B(n_1688),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1710),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1713),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1712),
.B(n_1678),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1713),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1747),
.B(n_1678),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1715),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1715),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1716),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1721),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1716),
.Y(n_1777)
);

NOR2xp67_ASAP7_75t_L g1778 ( 
.A(n_1738),
.B(n_1699),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1717),
.Y(n_1779)
);

OR2x2_ASAP7_75t_L g1780 ( 
.A(n_1732),
.B(n_1690),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1728),
.B(n_1733),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1749),
.B(n_1688),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1728),
.B(n_1686),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1718),
.B(n_1688),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1717),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1733),
.B(n_1668),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1718),
.B(n_1688),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1752),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1756),
.B(n_1740),
.C(n_1722),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_SL g1790 ( 
.A(n_1756),
.B(n_1721),
.Y(n_1790)
);

OAI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1764),
.A2(n_1722),
.B(n_1745),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1752),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1763),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1768),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1765),
.B(n_1722),
.C(n_1736),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1772),
.B(n_1763),
.Y(n_1796)
);

OAI21xp5_ASAP7_75t_L g1797 ( 
.A1(n_1764),
.A2(n_1722),
.B(n_1745),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1768),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1763),
.B(n_1711),
.Y(n_1799)
);

O2A1O1Ixp5_ASAP7_75t_L g1800 ( 
.A1(n_1761),
.A2(n_1737),
.B(n_1736),
.C(n_1724),
.Y(n_1800)
);

OAI21xp33_ASAP7_75t_L g1801 ( 
.A1(n_1786),
.A2(n_1730),
.B(n_1751),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1769),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1767),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1753),
.B(n_1737),
.Y(n_1804)
);

AOI22xp5_ASAP7_75t_L g1805 ( 
.A1(n_1778),
.A2(n_1638),
.B1(n_1682),
.B2(n_1626),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_SL g1806 ( 
.A1(n_1758),
.A2(n_1745),
.B(n_1751),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_SL g1807 ( 
.A(n_1759),
.B(n_1724),
.C(n_1735),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1778),
.B(n_1727),
.C(n_1726),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1758),
.B(n_1723),
.Y(n_1809)
);

OAI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1780),
.A2(n_1776),
.B1(n_1762),
.B2(n_1766),
.Y(n_1810)
);

NOR2xp67_ASAP7_75t_SL g1811 ( 
.A(n_1776),
.B(n_1490),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1769),
.Y(n_1812)
);

A2O1A1Ixp33_ASAP7_75t_L g1813 ( 
.A1(n_1780),
.A2(n_1682),
.B(n_1706),
.C(n_1746),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1771),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1800),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1789),
.B(n_1760),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1793),
.Y(n_1817)
);

AOI222xp33_ASAP7_75t_L g1818 ( 
.A1(n_1790),
.A2(n_1776),
.B1(n_1760),
.B2(n_1706),
.C1(n_1695),
.C2(n_1684),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1809),
.B(n_1767),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1788),
.Y(n_1820)
);

OAI222xp33_ASAP7_75t_L g1821 ( 
.A1(n_1790),
.A2(n_1766),
.B1(n_1770),
.B2(n_1757),
.C1(n_1781),
.C2(n_1754),
.Y(n_1821)
);

OR2x2_ASAP7_75t_L g1822 ( 
.A(n_1796),
.B(n_1770),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1799),
.Y(n_1823)
);

OAI22xp5_ASAP7_75t_L g1824 ( 
.A1(n_1807),
.A2(n_1742),
.B1(n_1743),
.B2(n_1729),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_L g1825 ( 
.A1(n_1795),
.A2(n_1757),
.B(n_1771),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1800),
.A2(n_1783),
.B(n_1755),
.Y(n_1826)
);

AOI332xp33_ASAP7_75t_L g1827 ( 
.A1(n_1792),
.A2(n_1774),
.A3(n_1785),
.B1(n_1773),
.B2(n_1775),
.B3(n_1779),
.C1(n_1777),
.C2(n_1755),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1804),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1801),
.B(n_1784),
.Y(n_1829)
);

A2O1A1Ixp33_ASAP7_75t_L g1830 ( 
.A1(n_1791),
.A2(n_1732),
.B(n_1746),
.C(n_1684),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1803),
.B(n_1782),
.Y(n_1831)
);

OAI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1797),
.A2(n_1750),
.B1(n_1629),
.B2(n_1742),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1807),
.Y(n_1833)
);

XOR2x2_ASAP7_75t_L g1834 ( 
.A(n_1816),
.B(n_1808),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1823),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1822),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1822),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1819),
.B(n_1810),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1831),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1815),
.B(n_1794),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1831),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1820),
.Y(n_1842)
);

AOI221x1_ASAP7_75t_L g1843 ( 
.A1(n_1815),
.A2(n_1814),
.B1(n_1798),
.B2(n_1812),
.C(n_1802),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1821),
.B(n_1820),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1839),
.B(n_1828),
.Y(n_1845)
);

NOR3xp33_ASAP7_75t_L g1846 ( 
.A(n_1844),
.B(n_1833),
.C(n_1825),
.Y(n_1846)
);

INVxp67_ASAP7_75t_L g1847 ( 
.A(n_1838),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1841),
.Y(n_1848)
);

AOI211x1_ASAP7_75t_L g1849 ( 
.A1(n_1840),
.A2(n_1826),
.B(n_1829),
.C(n_1810),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1836),
.Y(n_1850)
);

AOI221xp5_ASAP7_75t_L g1851 ( 
.A1(n_1840),
.A2(n_1830),
.B1(n_1817),
.B2(n_1832),
.C(n_1813),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1837),
.B(n_1819),
.Y(n_1852)
);

OAI211xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1835),
.A2(n_1806),
.B(n_1818),
.C(n_1827),
.Y(n_1853)
);

NAND3xp33_ASAP7_75t_SL g1854 ( 
.A(n_1842),
.B(n_1817),
.C(n_1813),
.Y(n_1854)
);

AOI21xp5_ASAP7_75t_L g1855 ( 
.A1(n_1846),
.A2(n_1834),
.B(n_1843),
.Y(n_1855)
);

NOR3xp33_ASAP7_75t_SL g1856 ( 
.A(n_1853),
.B(n_1824),
.C(n_1774),
.Y(n_1856)
);

NAND2xp33_ASAP7_75t_SL g1857 ( 
.A(n_1852),
.B(n_1773),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1849),
.A2(n_1805),
.B1(n_1775),
.B2(n_1777),
.C(n_1785),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1850),
.Y(n_1859)
);

AOI22xp5_ASAP7_75t_L g1860 ( 
.A1(n_1856),
.A2(n_1847),
.B1(n_1851),
.B2(n_1854),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1855),
.A2(n_1848),
.B1(n_1845),
.B2(n_1779),
.C(n_1754),
.Y(n_1861)
);

OAI22xp5_ASAP7_75t_L g1862 ( 
.A1(n_1858),
.A2(n_1750),
.B1(n_1743),
.B2(n_1729),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1859),
.B(n_1811),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1857),
.B(n_1782),
.Y(n_1864)
);

NOR3xp33_ASAP7_75t_L g1865 ( 
.A(n_1855),
.B(n_1685),
.C(n_1684),
.Y(n_1865)
);

NOR2x1_ASAP7_75t_L g1866 ( 
.A(n_1864),
.B(n_1863),
.Y(n_1866)
);

NAND4xp75_ASAP7_75t_L g1867 ( 
.A(n_1860),
.B(n_1787),
.C(n_1784),
.D(n_1723),
.Y(n_1867)
);

NAND4xp75_ASAP7_75t_L g1868 ( 
.A(n_1861),
.B(n_1787),
.C(n_1744),
.D(n_1727),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1865),
.A2(n_1726),
.B1(n_1682),
.B2(n_1748),
.Y(n_1869)
);

AND3x2_ASAP7_75t_L g1870 ( 
.A(n_1862),
.B(n_1744),
.C(n_1748),
.Y(n_1870)
);

HB1xp67_ASAP7_75t_L g1871 ( 
.A(n_1866),
.Y(n_1871)
);

AOI21xp33_ASAP7_75t_SL g1872 ( 
.A1(n_1869),
.A2(n_1702),
.B(n_1696),
.Y(n_1872)
);

OAI211xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1868),
.A2(n_1692),
.B(n_1684),
.C(n_1695),
.Y(n_1873)
);

AOI21xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1871),
.A2(n_1867),
.B(n_1870),
.Y(n_1874)
);

OA22x2_ASAP7_75t_L g1875 ( 
.A1(n_1874),
.A2(n_1873),
.B1(n_1872),
.B2(n_1694),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1708),
.B1(n_1696),
.B2(n_1702),
.Y(n_1876)
);

NOR3xp33_ASAP7_75t_L g1877 ( 
.A(n_1875),
.B(n_1692),
.C(n_1685),
.Y(n_1877)
);

AOI22x1_ASAP7_75t_L g1878 ( 
.A1(n_1877),
.A2(n_1665),
.B1(n_1659),
.B2(n_1683),
.Y(n_1878)
);

AOI21xp5_ASAP7_75t_L g1879 ( 
.A1(n_1876),
.A2(n_1702),
.B(n_1696),
.Y(n_1879)
);

AO22x2_ASAP7_75t_L g1880 ( 
.A1(n_1879),
.A2(n_1708),
.B1(n_1702),
.B2(n_1696),
.Y(n_1880)
);

AOI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1878),
.A2(n_1708),
.B(n_1692),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1881),
.A2(n_1692),
.B(n_1685),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1882),
.B(n_1880),
.Y(n_1883)
);

O2A1O1Ixp33_ASAP7_75t_L g1884 ( 
.A1(n_1883),
.A2(n_1565),
.B(n_1685),
.C(n_1695),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_R g1885 ( 
.A1(n_1884),
.A2(n_1693),
.B1(n_1683),
.B2(n_1602),
.C(n_1665),
.Y(n_1885)
);

AOI211xp5_ASAP7_75t_L g1886 ( 
.A1(n_1885),
.A2(n_1604),
.B(n_1560),
.C(n_1561),
.Y(n_1886)
);


endmodule