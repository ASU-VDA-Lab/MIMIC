module fake_jpeg_2923_n_101 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_101);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_101;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_35),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_31),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_36),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_37),
.B1(n_38),
.B2(n_36),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_51),
.A2(n_55),
.B1(n_56),
.B2(n_59),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_38),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_33),
.B1(n_29),
.B2(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_1),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_58),
.A2(n_47),
.B1(n_30),
.B2(n_49),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_64),
.A2(n_69),
.B(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_43),
.B1(n_30),
.B2(n_40),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_26),
.B1(n_25),
.B2(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_40),
.B1(n_30),
.B2(n_49),
.Y(n_67)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_67),
.A2(n_34),
.B1(n_12),
.B2(n_14),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_2),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_3),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_76),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_75),
.A2(n_67),
.B1(n_6),
.B2(n_7),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_4),
.Y(n_77)
);

AOI322xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_78),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_4),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_81),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_82),
.B(n_83),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_64),
.C(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_88),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_94),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_86),
.B(n_87),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

OAI221xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_85),
.B1(n_90),
.B2(n_92),
.C(n_81),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_91),
.B(n_84),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_15),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_19),
.C(n_20),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_21),
.C(n_10),
.Y(n_101)
);


endmodule