module fake_jpeg_9479_n_67 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_14),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_27),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_39),
.B(n_4),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_49),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_25),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_44),
.C(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_5),
.Y(n_44)
);

AO21x2_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_6),
.B(n_7),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_47),
.B1(n_40),
.B2(n_46),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_24),
.B1(n_10),
.B2(n_11),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_9),
.C(n_13),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_16),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_51),
.B(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_53),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_45),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_56),
.B(n_50),
.Y(n_61)
);

XNOR2x1_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_59),
.Y(n_64)
);

AOI31xp67_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_56),
.A3(n_45),
.B(n_55),
.Y(n_65)
);

AOI322xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_43),
.A3(n_58),
.B1(n_57),
.B2(n_52),
.C1(n_41),
.C2(n_23),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_22),
.Y(n_67)
);


endmodule