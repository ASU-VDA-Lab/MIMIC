module fake_jpeg_30618_n_324 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_0),
.B(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx8_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx2_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_40),
.Y(n_86)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_15),
.B(n_13),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_45),
.B(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_20),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_22),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_54),
.Y(n_96)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_57),
.Y(n_95)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_62),
.Y(n_88)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_64),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_16),
.B(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_23),
.Y(n_78)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_22),
.B1(n_34),
.B2(n_32),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_72),
.A2(n_112),
.B1(n_113),
.B2(n_86),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_30),
.B1(n_25),
.B2(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_73),
.A2(n_75),
.B1(n_90),
.B2(n_94),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_25),
.B1(n_30),
.B2(n_28),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_23),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_85),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_67),
.A2(n_25),
.B1(n_36),
.B2(n_19),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_89),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_18),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_46),
.B(n_36),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_91),
.B(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_51),
.A2(n_30),
.B1(n_18),
.B2(n_34),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_57),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_52),
.B(n_28),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_105),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_56),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_26),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_61),
.A2(n_31),
.B1(n_24),
.B2(n_34),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_44),
.A2(n_37),
.B1(n_29),
.B2(n_21),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_57),
.A2(n_37),
.B1(n_29),
.B2(n_21),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_18),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_7),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_62),
.A2(n_7),
.B1(n_10),
.B2(n_8),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_10),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_154),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_114),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_119),
.B(n_140),
.Y(n_155)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_4),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_123),
.B(n_138),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

BUFx4f_ASAP7_75t_SL g182 ( 
.A(n_124),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_128),
.Y(n_188)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_82),
.Y(n_132)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_4),
.C(n_8),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_106),
.Y(n_164)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_147),
.Y(n_156)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_137),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_12),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_86),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_74),
.B(n_76),
.Y(n_168)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_149),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_72),
.A2(n_112),
.B1(n_113),
.B2(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_145),
.B1(n_106),
.B2(n_89),
.Y(n_158)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_144),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_100),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_82),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_1),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_153),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_96),
.B(n_2),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_108),
.Y(n_181)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_109),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_158),
.A2(n_161),
.B1(n_166),
.B2(n_180),
.Y(n_209)
);

BUFx24_ASAP7_75t_SL g160 ( 
.A(n_150),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_178),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_121),
.A2(n_101),
.B1(n_103),
.B2(n_102),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_102),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_164),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_101),
.B1(n_103),
.B2(n_81),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_73),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_167),
.B(n_174),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_173),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_71),
.Y(n_173)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_90),
.Y(n_174)
);

AND2x6_ASAP7_75t_L g178 ( 
.A(n_125),
.B(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_81),
.B1(n_77),
.B2(n_94),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_136),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_80),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_187),
.C(n_126),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_133),
.B(n_71),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_186),
.B(n_154),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_139),
.B(n_80),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_179),
.A2(n_145),
.B1(n_147),
.B2(n_146),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_162),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_193),
.B(n_196),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_134),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_187),
.B(n_129),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_198),
.Y(n_234)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_159),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_132),
.B(n_148),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_220),
.B(n_156),
.Y(n_236)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_165),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_155),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_210),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_157),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_211),
.Y(n_235)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_157),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_215),
.B(n_180),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_174),
.A2(n_130),
.B1(n_122),
.B2(n_153),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_217),
.Y(n_240)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_167),
.A2(n_136),
.B1(n_126),
.B2(n_128),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_219),
.B1(n_158),
.B2(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_161),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_230),
.A2(n_218),
.B1(n_216),
.B2(n_219),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_178),
.C(n_168),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_236),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_193),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_237),
.B(n_245),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_201),
.A2(n_221),
.B(n_197),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_239),
.A2(n_199),
.B(n_190),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_188),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_236),
.B(n_191),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_221),
.B(n_207),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_252),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_253),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_227),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_254),
.B(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_206),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_209),
.Y(n_257)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_223),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_259),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_200),
.Y(n_260)
);

AOI221xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.C(n_264),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_213),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_223),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_211),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_250),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_257),
.A2(n_264),
.B1(n_259),
.B2(n_258),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_269),
.B1(n_270),
.B2(n_263),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_267),
.B(n_280),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_230),
.B1(n_240),
.B2(n_225),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_240),
.B1(n_223),
.B2(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_245),
.C(n_237),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_272),
.B(n_278),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_251),
.C(n_232),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_225),
.C(n_222),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_273),
.B(n_254),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_283),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_256),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_288),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_274),
.A2(n_265),
.B1(n_252),
.B2(n_247),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_287),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_275),
.Y(n_287)
);

NOR3xp33_ASAP7_75t_SL g288 ( 
.A(n_277),
.B(n_249),
.C(n_255),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_289),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_271),
.A2(n_260),
.B1(n_261),
.B2(n_253),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_268),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_291),
.A2(n_292),
.B(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_269),
.B(n_228),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_262),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_277),
.B(n_266),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_294),
.B(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_272),
.C(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_301),
.C(n_285),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_271),
.C(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_270),
.C(n_274),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_276),
.B(n_248),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_304),
.B(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_309),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_283),
.B1(n_289),
.B2(n_276),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_310),
.Y(n_313)
);

OA21x2_ASAP7_75t_SL g308 ( 
.A1(n_303),
.A2(n_235),
.B(n_242),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_311),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_295),
.A2(n_241),
.B1(n_229),
.B2(n_244),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_301),
.C(n_297),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_299),
.B1(n_300),
.B2(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_314),
.B(n_311),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_306),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_316),
.B(n_318),
.Y(n_320)
);

AOI322xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_313),
.A3(n_314),
.B1(n_217),
.B2(n_208),
.C1(n_182),
.C2(n_244),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_315),
.B(n_305),
.C(n_241),
.Y(n_318)
);

AOI322xp5_ASAP7_75t_L g321 ( 
.A1(n_319),
.A2(n_182),
.A3(n_177),
.B1(n_154),
.B2(n_195),
.C1(n_185),
.C2(n_198),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_182),
.B(n_320),
.Y(n_322)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_198),
.B(n_203),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_128),
.Y(n_324)
);


endmodule