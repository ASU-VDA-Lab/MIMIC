module fake_netlist_1_7080_n_719 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_719);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_719;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g82 ( .A(n_10), .Y(n_82) );
INVx4_ASAP7_75t_R g83 ( .A(n_20), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_45), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_39), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_43), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_13), .Y(n_87) );
INVxp67_ASAP7_75t_SL g88 ( .A(n_10), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_8), .Y(n_89) );
CKINVDCx14_ASAP7_75t_R g90 ( .A(n_70), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_2), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_60), .Y(n_93) );
INVxp67_ASAP7_75t_L g94 ( .A(n_49), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_2), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_75), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_57), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_14), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_78), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_74), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_41), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_68), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_22), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_32), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_56), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_44), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_65), .Y(n_107) );
INVxp33_ASAP7_75t_L g108 ( .A(n_20), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_38), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_23), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_50), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_4), .Y(n_113) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_14), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_79), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_73), .B(n_62), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_28), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_63), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_35), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_24), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_33), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_52), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_17), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_69), .Y(n_125) );
INVx1_ASAP7_75t_SL g126 ( .A(n_59), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_46), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_40), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_23), .Y(n_129) );
INVxp33_ASAP7_75t_SL g130 ( .A(n_16), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_21), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_114), .B(n_0), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_82), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_97), .Y(n_134) );
CKINVDCx20_ASAP7_75t_R g135 ( .A(n_101), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_110), .B(n_0), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
OR2x6_ASAP7_75t_L g139 ( .A(n_91), .B(n_1), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_85), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_118), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g143 ( .A(n_112), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_117), .Y(n_144) );
INVxp67_ASAP7_75t_SL g145 ( .A(n_108), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_122), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_115), .B(n_1), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_111), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_90), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_86), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_92), .B(n_3), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_92), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_98), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_93), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_93), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_82), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_91), .B(n_3), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_130), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g162 ( .A(n_82), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_82), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_87), .B(n_4), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_104), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_107), .B(n_31), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_96), .Y(n_167) );
CKINVDCx20_ASAP7_75t_R g168 ( .A(n_82), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_99), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_99), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_87), .B(n_5), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_100), .Y(n_172) );
NAND2x1_ASAP7_75t_L g173 ( .A(n_83), .B(n_5), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_89), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_100), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_102), .Y(n_176) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_171), .B(n_164), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
INVxp67_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_171), .B(n_131), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_149), .B(n_94), .Y(n_183) );
INVx8_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_138), .B(n_125), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_142), .Y(n_187) );
AO22x2_ASAP7_75t_L g188 ( .A1(n_171), .A2(n_102), .B1(n_105), .B2(n_106), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_135), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_138), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_140), .B(n_128), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_170), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_165), .B(n_109), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_140), .B(n_119), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_163), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_174), .A2(n_131), .B1(n_129), .B2(n_89), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_171), .B(n_119), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_141), .B(n_120), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_162), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_168), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_139), .B(n_129), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_154), .B(n_120), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_141), .B(n_106), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_170), .Y(n_206) );
AO22x2_ASAP7_75t_L g207 ( .A1(n_173), .A2(n_105), .B1(n_95), .B2(n_124), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_142), .Y(n_208) );
INVxp67_ASAP7_75t_SL g209 ( .A(n_150), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_150), .B(n_95), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_139), .A2(n_103), .B1(n_124), .B2(n_123), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
BUFx2_ASAP7_75t_L g214 ( .A(n_139), .Y(n_214) );
INVxp67_ASAP7_75t_L g215 ( .A(n_161), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_139), .A2(n_103), .B1(n_123), .B2(n_113), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_134), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_170), .Y(n_219) );
INVxp67_ASAP7_75t_L g220 ( .A(n_144), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_133), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_153), .B(n_127), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_153), .B(n_113), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_160), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_133), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_133), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_160), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_133), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_156), .B(n_126), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_157), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_160), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_160), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
NAND2xp33_ASAP7_75t_L g234 ( .A(n_156), .B(n_121), .Y(n_234) );
OAI22xp5_ASAP7_75t_L g235 ( .A1(n_132), .A2(n_88), .B1(n_116), .B2(n_8), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_167), .B(n_6), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_167), .B(n_6), .Y(n_237) );
INVx4_ASAP7_75t_L g238 ( .A(n_160), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_169), .B(n_36), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_157), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_169), .B(n_34), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_136), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_184), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_203), .B(n_164), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_184), .Y(n_245) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_190), .A2(n_172), .B(n_175), .Y(n_246) );
INVx5_ASAP7_75t_L g247 ( .A(n_199), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_209), .B(n_190), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_186), .B(n_175), .Y(n_249) );
NOR2xp33_ASAP7_75t_R g250 ( .A(n_189), .B(n_146), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_191), .B(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_223), .B(n_158), .Y(n_252) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_202), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_184), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_201), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_184), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_177), .B(n_137), .Y(n_257) );
NAND2xp33_ASAP7_75t_R g258 ( .A(n_214), .B(n_166), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_203), .Y(n_259) );
AO22x1_ASAP7_75t_L g260 ( .A1(n_203), .A2(n_158), .B1(n_136), .B2(n_155), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_236), .Y(n_262) );
BUFx2_ASAP7_75t_L g263 ( .A(n_214), .Y(n_263) );
INVx8_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_236), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_179), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_236), .Y(n_267) );
AND2x4_ASAP7_75t_L g268 ( .A(n_181), .B(n_173), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_223), .B(n_147), .Y(n_269) );
INVx4_ASAP7_75t_L g270 ( .A(n_199), .Y(n_270) );
NOR2xp33_ASAP7_75t_R g271 ( .A(n_189), .B(n_143), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_179), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_210), .B(n_159), .Y(n_273) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_178), .A2(n_152), .B1(n_159), .B2(n_155), .Y(n_274) );
AND2x4_ASAP7_75t_L g275 ( .A(n_181), .B(n_176), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_223), .B(n_176), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_187), .Y(n_277) );
CKINVDCx6p67_ASAP7_75t_R g278 ( .A(n_199), .Y(n_278) );
NAND2x1p5_ASAP7_75t_L g279 ( .A(n_181), .B(n_151), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_187), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_208), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_178), .B(n_151), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_242), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_210), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_208), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_178), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_199), .B(n_157), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_242), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_242), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_212), .B(n_157), .Y(n_291) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_180), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_188), .Y(n_293) );
INVx4_ASAP7_75t_L g294 ( .A(n_199), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_188), .Y(n_295) );
NOR3xp33_ASAP7_75t_SL g296 ( .A(n_235), .B(n_7), .C(n_9), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_198), .B(n_7), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_216), .Y(n_298) );
NAND2x1p5_ASAP7_75t_L g299 ( .A(n_194), .B(n_163), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_224), .Y(n_300) );
NOR2xp33_ASAP7_75t_R g301 ( .A(n_215), .B(n_42), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_217), .A2(n_163), .B1(n_11), .B2(n_12), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_188), .B(n_9), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_188), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_237), .Y(n_305) );
BUFx12f_ASAP7_75t_L g306 ( .A(n_199), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_239), .B(n_163), .Y(n_307) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_185), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_224), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_207), .Y(n_310) );
CKINVDCx20_ASAP7_75t_R g311 ( .A(n_220), .Y(n_311) );
AND3x1_ASAP7_75t_SL g312 ( .A(n_207), .B(n_12), .C(n_13), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_200), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_313), .B(n_207), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_310), .Y(n_315) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_293), .A2(n_207), .B1(n_234), .B2(n_222), .Y(n_316) );
INVx2_ASAP7_75t_SL g317 ( .A(n_256), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_284), .B(n_193), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_262), .Y(n_319) );
AOI22xp5_ASAP7_75t_L g320 ( .A1(n_310), .A2(n_234), .B1(n_205), .B2(n_204), .Y(n_320) );
NAND3xp33_ASAP7_75t_L g321 ( .A(n_296), .B(n_241), .C(n_238), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_313), .B(n_229), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_283), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_262), .Y(n_325) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_265), .A2(n_183), .B1(n_238), .B2(n_182), .Y(n_326) );
CKINVDCx8_ASAP7_75t_R g327 ( .A(n_264), .Y(n_327) );
INVx2_ASAP7_75t_SL g328 ( .A(n_256), .Y(n_328) );
BUFx2_ASAP7_75t_L g329 ( .A(n_256), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_270), .B(n_238), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_256), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_271), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_256), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g334 ( .A1(n_297), .A2(n_240), .B(n_221), .C(n_225), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_270), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_250), .Y(n_336) );
AND2x6_ASAP7_75t_L g337 ( .A(n_245), .B(n_195), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_253), .B(n_15), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_293), .A2(n_195), .B1(n_185), .B2(n_232), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_289), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_270), .B(n_232), .Y(n_341) );
INVx1_ASAP7_75t_SL g342 ( .A(n_263), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_289), .Y(n_343) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_264), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_244), .B(n_15), .Y(n_345) );
OR2x6_ASAP7_75t_L g346 ( .A(n_264), .B(n_227), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_249), .A2(n_219), .B(n_213), .Y(n_347) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_264), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_290), .Y(n_349) );
AND3x1_ASAP7_75t_SL g350 ( .A(n_311), .B(n_16), .C(n_17), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_306), .Y(n_351) );
BUFx3_ASAP7_75t_L g352 ( .A(n_306), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_295), .A2(n_304), .B1(n_268), .B2(n_303), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_290), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_266), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_265), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_266), .Y(n_357) );
INVx2_ASAP7_75t_SL g358 ( .A(n_245), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_279), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_278), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_272), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_244), .B(n_18), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_244), .B(n_18), .Y(n_363) );
INVx3_ASAP7_75t_L g364 ( .A(n_294), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_272), .Y(n_365) );
BUFx2_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
AND2x6_ASAP7_75t_L g367 ( .A(n_254), .B(n_219), .Y(n_367) );
INVx5_ASAP7_75t_L g368 ( .A(n_294), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g369 ( .A(n_311), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_322), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_345), .Y(n_371) );
AOI22xp33_ASAP7_75t_SL g372 ( .A1(n_342), .A2(n_303), .B1(n_297), .B2(n_304), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_355), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_355), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_369), .Y(n_375) );
AND2x4_ASAP7_75t_L g376 ( .A(n_359), .B(n_286), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_314), .A2(n_295), .B1(n_268), .B2(n_275), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_347), .A2(n_307), .B(n_246), .Y(n_378) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_320), .A2(n_267), .B1(n_252), .B2(n_279), .Y(n_379) );
INVx4_ASAP7_75t_SL g380 ( .A(n_337), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_353), .A2(n_279), .B1(n_278), .B2(n_286), .Y(n_381) );
AOI21xp5_ASAP7_75t_L g382 ( .A1(n_355), .A2(n_251), .B(n_248), .Y(n_382) );
OR2x6_ASAP7_75t_L g383 ( .A(n_315), .B(n_243), .Y(n_383) );
INVxp67_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_327), .Y(n_385) );
AOI21xp5_ASAP7_75t_SL g386 ( .A1(n_346), .A2(n_294), .B(n_243), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_345), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_336), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_359), .B(n_268), .Y(n_389) );
OR2x6_ASAP7_75t_L g390 ( .A(n_315), .B(n_260), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_357), .A2(n_305), .B(n_269), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_338), .B(n_257), .Y(n_392) );
BUFx12f_ASAP7_75t_L g393 ( .A(n_332), .Y(n_393) );
AOI221xp5_ASAP7_75t_L g394 ( .A1(n_318), .A2(n_255), .B1(n_261), .B2(n_273), .C(n_292), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_351), .B(n_263), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g396 ( .A1(n_320), .A2(n_259), .B1(n_305), .B2(n_275), .Y(n_396) );
AOI211x1_ASAP7_75t_L g397 ( .A1(n_314), .A2(n_260), .B(n_274), .C(n_282), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_363), .Y(n_398) );
INVx4_ASAP7_75t_L g399 ( .A(n_337), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_316), .A2(n_327), .B1(n_275), .B2(n_276), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_363), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_368), .B(n_247), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_334), .B(n_273), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_338), .B(n_291), .Y(n_404) );
AOI222xp33_ASAP7_75t_L g405 ( .A1(n_392), .A2(n_325), .B1(n_319), .B2(n_356), .C1(n_302), .C2(n_362), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_402), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_372), .B(n_319), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_394), .A2(n_379), .B1(n_403), .B2(n_401), .C(n_371), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_373), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_372), .A2(n_321), .B1(n_356), .B2(n_325), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_370), .B(n_323), .Y(n_413) );
INVx4_ASAP7_75t_L g414 ( .A(n_380), .Y(n_414) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_391), .A2(n_321), .B(n_326), .C(n_358), .Y(n_415) );
BUFx2_ASAP7_75t_L g416 ( .A(n_376), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_382), .A2(n_326), .B(n_349), .Y(n_417) );
AOI22xp33_ASAP7_75t_SL g418 ( .A1(n_390), .A2(n_366), .B1(n_350), .B2(n_301), .Y(n_418) );
AOI22xp33_ASAP7_75t_SL g419 ( .A1(n_390), .A2(n_366), .B1(n_351), .B2(n_352), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_374), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_376), .B(n_323), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g422 ( .A1(n_390), .A2(n_258), .B1(n_358), .B2(n_352), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_333), .B1(n_329), .B2(n_331), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_376), .B(n_323), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_396), .A2(n_333), .B1(n_331), .B2(n_329), .Y(n_425) );
OAI211xp5_ASAP7_75t_L g426 ( .A1(n_384), .A2(n_312), .B(n_339), .C(n_288), .Y(n_426) );
OR2x6_ASAP7_75t_L g427 ( .A(n_386), .B(n_346), .Y(n_427) );
INVxp33_ASAP7_75t_L g428 ( .A(n_395), .Y(n_428) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_387), .A2(n_349), .B1(n_340), .B2(n_343), .C(n_324), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_384), .Y(n_430) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_395), .A2(n_352), .B1(n_351), .B2(n_337), .Y(n_431) );
AO21x2_ASAP7_75t_L g432 ( .A1(n_378), .A2(n_324), .B(n_340), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g433 ( .A1(n_398), .A2(n_324), .B1(n_340), .B2(n_349), .C(n_354), .Y(n_433) );
AND4x1_ASAP7_75t_L g434 ( .A(n_375), .B(n_19), .C(n_21), .D(n_22), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_416), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_408), .B(n_377), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_427), .B(n_399), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_408), .B(n_397), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g440 ( .A(n_430), .Y(n_440) );
NOR2xp33_ASAP7_75t_SL g441 ( .A(n_427), .B(n_399), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g442 ( .A1(n_409), .A2(n_404), .B(n_377), .C(n_400), .Y(n_442) );
AOI222xp33_ASAP7_75t_L g443 ( .A1(n_412), .A2(n_389), .B1(n_381), .B2(n_393), .C1(n_380), .C2(n_385), .Y(n_443) );
NOR3xp33_ASAP7_75t_L g444 ( .A(n_418), .B(n_388), .C(n_385), .Y(n_444) );
AO21x2_ASAP7_75t_L g445 ( .A1(n_417), .A2(n_233), .B(n_227), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_432), .Y(n_446) );
OAI321xp33_ASAP7_75t_L g447 ( .A1(n_422), .A2(n_423), .A3(n_426), .B1(n_425), .B2(n_417), .C(n_416), .Y(n_447) );
NOR2xp33_ASAP7_75t_R g448 ( .A(n_407), .B(n_388), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_421), .B(n_389), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_407), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_432), .Y(n_451) );
INVx3_ASAP7_75t_SL g452 ( .A(n_407), .Y(n_452) );
OAI211xp5_ASAP7_75t_L g453 ( .A1(n_419), .A2(n_163), .B(n_343), .C(n_354), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_407), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_413), .A2(n_383), .B1(n_343), .B2(n_354), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_405), .A2(n_383), .B1(n_393), .B2(n_337), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_421), .B(n_380), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_413), .B(n_410), .Y(n_459) );
NOR4xp25_ASAP7_75t_SL g460 ( .A(n_410), .B(n_383), .C(n_19), .D(n_206), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_405), .A2(n_337), .B1(n_367), .B2(n_317), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_411), .B(n_357), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_411), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_424), .Y(n_464) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_428), .A2(n_360), .B1(n_368), .B2(n_317), .Y(n_465) );
OAI321xp33_ASAP7_75t_L g466 ( .A1(n_427), .A2(n_328), .A3(n_307), .B1(n_299), .B2(n_233), .C(n_231), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_424), .B(n_365), .Y(n_467) );
AOI21x1_ASAP7_75t_L g468 ( .A1(n_427), .A2(n_231), .B(n_182), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_432), .Y(n_469) );
INVx3_ASAP7_75t_L g470 ( .A(n_414), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_442), .A2(n_431), .B1(n_433), .B2(n_429), .Y(n_471) );
AOI221xp5_ASAP7_75t_L g472 ( .A1(n_457), .A2(n_420), .B1(n_434), .B2(n_415), .C(n_407), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_448), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_436), .B(n_420), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_438), .B(n_427), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_439), .B(n_414), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_438), .B(n_434), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_456), .B(n_414), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_456), .Y(n_479) );
BUFx2_ASAP7_75t_L g480 ( .A(n_435), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g481 ( .A1(n_455), .A2(n_414), .B1(n_337), .B2(n_367), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_436), .B(n_365), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_439), .B(n_365), .Y(n_483) );
INVx1_ASAP7_75t_SL g484 ( .A(n_452), .Y(n_484) );
BUFx2_ASAP7_75t_SL g485 ( .A(n_470), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_463), .B(n_357), .Y(n_486) );
BUFx2_ASAP7_75t_L g487 ( .A(n_435), .Y(n_487) );
NAND3xp33_ASAP7_75t_L g488 ( .A(n_443), .B(n_192), .C(n_206), .Y(n_488) );
INVx1_ASAP7_75t_SL g489 ( .A(n_452), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_463), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_459), .B(n_361), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_446), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_446), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_464), .B(n_361), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_452), .Y(n_496) );
BUFx2_ASAP7_75t_L g497 ( .A(n_455), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_467), .B(n_361), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_467), .B(n_25), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_449), .B(n_26), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_446), .Y(n_501) );
AOI22xp33_ASAP7_75t_SL g502 ( .A1(n_441), .A2(n_337), .B1(n_367), .B2(n_402), .Y(n_502) );
OAI31xp33_ASAP7_75t_L g503 ( .A1(n_453), .A2(n_402), .A3(n_328), .B(n_360), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_451), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_451), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_440), .B(n_368), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_454), .B(n_337), .Y(n_507) );
OAI31xp33_ASAP7_75t_L g508 ( .A1(n_461), .A2(n_444), .A3(n_441), .B(n_465), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_450), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_449), .B(n_27), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_462), .B(n_29), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_451), .Y(n_512) );
BUFx3_ASAP7_75t_L g513 ( .A(n_454), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_469), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_462), .B(n_30), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_469), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_469), .B(n_299), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_454), .B(n_37), .Y(n_518) );
HB1xp67_ASAP7_75t_L g519 ( .A(n_458), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_445), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_443), .B(n_367), .Y(n_521) );
OAI31xp33_ASAP7_75t_L g522 ( .A1(n_470), .A2(n_360), .A3(n_330), .B(n_364), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_492), .B(n_458), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_479), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_477), .B(n_490), .Y(n_525) );
INVx2_ASAP7_75t_SL g526 ( .A(n_473), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_473), .Y(n_527) );
NAND2x1_ASAP7_75t_L g528 ( .A(n_497), .B(n_437), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_474), .B(n_437), .Y(n_529) );
BUFx12f_ASAP7_75t_L g530 ( .A(n_498), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_519), .B(n_437), .Y(n_531) );
NAND2xp33_ASAP7_75t_SL g532 ( .A(n_497), .B(n_470), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_475), .B(n_445), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_477), .B(n_470), .Y(n_534) );
OAI211xp5_ASAP7_75t_SL g535 ( .A1(n_472), .A2(n_192), .B(n_196), .C(n_213), .Y(n_535) );
CKINVDCx16_ASAP7_75t_R g536 ( .A(n_509), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_474), .B(n_437), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_495), .B(n_460), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_486), .B(n_437), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_486), .B(n_460), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_475), .B(n_445), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_493), .B(n_445), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_509), .B(n_47), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_478), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_485), .Y(n_545) );
OAI211xp5_ASAP7_75t_L g546 ( .A1(n_472), .A2(n_468), .B(n_447), .C(n_196), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_478), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_488), .B(n_447), .C(n_466), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_495), .B(n_48), .Y(n_549) );
OR2x2_ASAP7_75t_L g550 ( .A(n_480), .B(n_51), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_493), .B(n_468), .Y(n_552) );
INVx3_ASAP7_75t_L g553 ( .A(n_504), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_488), .B(n_466), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_498), .B(n_53), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
NAND2xp33_ASAP7_75t_L g557 ( .A(n_521), .B(n_484), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_480), .B(n_54), .Y(n_558) );
NAND4xp25_ASAP7_75t_L g559 ( .A(n_508), .B(n_240), .C(n_221), .D(n_225), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_487), .B(n_58), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_494), .B(n_61), .Y(n_561) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_481), .A2(n_367), .B(n_307), .Y(n_562) );
NAND3x1_ASAP7_75t_L g563 ( .A(n_508), .B(n_335), .C(n_364), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_487), .B(n_491), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_483), .Y(n_565) );
OR2x2_ASAP7_75t_L g566 ( .A(n_482), .B(n_476), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_499), .B(n_64), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_484), .Y(n_568) );
BUFx4f_ASAP7_75t_L g569 ( .A(n_499), .Y(n_569) );
NOR3xp33_ASAP7_75t_SL g570 ( .A(n_506), .B(n_226), .C(n_228), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_483), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_476), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_489), .B(n_66), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_494), .B(n_67), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_471), .B(n_72), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_481), .B(n_368), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_521), .A2(n_367), .B1(n_346), .B2(n_341), .Y(n_577) );
NOR4xp25_ASAP7_75t_SL g578 ( .A(n_502), .B(n_76), .C(n_77), .D(n_80), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_489), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_504), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_482), .B(n_367), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_536), .B(n_496), .Y(n_582) );
INVxp67_ASAP7_75t_L g583 ( .A(n_526), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g584 ( .A1(n_575), .A2(n_471), .B(n_502), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_564), .B(n_525), .Y(n_585) );
NAND2xp5_ASAP7_75t_SL g586 ( .A(n_569), .B(n_496), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_569), .A2(n_485), .B1(n_500), .B2(n_510), .Y(n_587) );
AOI211x1_ASAP7_75t_L g588 ( .A1(n_534), .A2(n_500), .B(n_510), .C(n_507), .Y(n_588) );
NAND2xp33_ASAP7_75t_SL g589 ( .A(n_528), .B(n_518), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_524), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_569), .A2(n_503), .B(n_522), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_572), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_566), .B(n_544), .Y(n_593) );
OAI32xp33_ASAP7_75t_L g594 ( .A1(n_527), .A2(n_507), .A3(n_513), .B1(n_518), .B2(n_511), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_575), .A2(n_511), .B1(n_515), .B2(n_513), .Y(n_595) );
AOI322xp5_ASAP7_75t_L g596 ( .A1(n_548), .A2(n_515), .A3(n_514), .B1(n_501), .B2(n_516), .C1(n_505), .C2(n_512), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_547), .B(n_513), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_526), .B(n_81), .Y(n_598) );
NAND2xp33_ASAP7_75t_L g599 ( .A(n_563), .B(n_501), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_530), .B(n_576), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_565), .Y(n_601) );
O2A1O1Ixp33_ASAP7_75t_L g602 ( .A1(n_535), .A2(n_503), .B(n_522), .C(n_516), .Y(n_602) );
OAI21xp33_ASAP7_75t_L g603 ( .A1(n_554), .A2(n_514), .B(n_512), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_530), .B(n_512), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_571), .B(n_505), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_568), .B(n_505), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_551), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_523), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_576), .A2(n_517), .B(n_520), .C(n_368), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_563), .A2(n_520), .B1(n_517), .B2(n_367), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g611 ( .A1(n_554), .A2(n_346), .B1(n_341), .B2(n_330), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_537), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_579), .B(n_299), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_539), .B(n_346), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_531), .B(n_197), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_538), .A2(n_341), .B1(n_330), .B2(n_335), .Y(n_616) );
OAI322xp33_ASAP7_75t_L g617 ( .A1(n_529), .A2(n_197), .A3(n_211), .B1(n_226), .B2(n_228), .C1(n_230), .C2(n_298), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_540), .B(n_197), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_543), .B(n_335), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_556), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_580), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_533), .B(n_197), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_533), .B(n_197), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_552), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_545), .B(n_211), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_SL g626 ( .A1(n_546), .A2(n_364), .B(n_335), .C(n_230), .Y(n_626) );
OAI322xp33_ASAP7_75t_L g627 ( .A1(n_549), .A2(n_211), .A3(n_300), .B1(n_277), .B2(n_280), .C1(n_281), .C2(n_285), .Y(n_627) );
O2A1O1Ixp5_ASAP7_75t_L g628 ( .A1(n_532), .A2(n_341), .B(n_330), .C(n_277), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_538), .B(n_211), .C(n_308), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_570), .A2(n_364), .B(n_300), .C(n_280), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_541), .B(n_211), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_584), .B(n_557), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_608), .B(n_541), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_624), .B(n_553), .Y(n_634) );
XNOR2x1_ASAP7_75t_L g635 ( .A(n_593), .B(n_550), .Y(n_635) );
OR2x6_ASAP7_75t_L g636 ( .A(n_609), .B(n_552), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_612), .B(n_553), .Y(n_637) );
NOR2xp33_ASAP7_75t_R g638 ( .A(n_589), .B(n_532), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_606), .B(n_553), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_595), .A2(n_557), .B1(n_560), .B2(n_558), .Y(n_640) );
INVx1_ASAP7_75t_SL g641 ( .A(n_582), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_590), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_592), .B(n_542), .Y(n_643) );
BUFx2_ASAP7_75t_L g644 ( .A(n_583), .Y(n_644) );
NOR2xp33_ASAP7_75t_R g645 ( .A(n_599), .B(n_567), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_585), .B(n_542), .Y(n_646) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_629), .B(n_562), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_607), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_601), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_622), .B(n_561), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_604), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_591), .A2(n_577), .B1(n_581), .B2(n_573), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_597), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_600), .B(n_616), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_605), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_619), .B(n_555), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_620), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_586), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_588), .B(n_561), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_596), .B(n_574), .Y(n_660) );
AND2x2_ASAP7_75t_L g661 ( .A(n_631), .B(n_574), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_621), .B(n_577), .Y(n_662) );
XNOR2xp5_ASAP7_75t_L g663 ( .A(n_587), .B(n_559), .Y(n_663) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_609), .B(n_578), .Y(n_664) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_591), .B(n_368), .Y(n_665) );
AND2x2_ASAP7_75t_L g666 ( .A(n_639), .B(n_603), .Y(n_666) );
OAI31xp33_ASAP7_75t_L g667 ( .A1(n_632), .A2(n_626), .A3(n_598), .B(n_602), .Y(n_667) );
AOI322xp5_ASAP7_75t_L g668 ( .A1(n_632), .A2(n_611), .A3(n_610), .B1(n_623), .B2(n_618), .C1(n_615), .C2(n_625), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_663), .A2(n_628), .B1(n_602), .B2(n_630), .C(n_614), .Y(n_669) );
AOI21xp5_ASAP7_75t_L g670 ( .A1(n_664), .A2(n_628), .B(n_594), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_SL g671 ( .A1(n_654), .A2(n_630), .B(n_613), .C(n_617), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_655), .B(n_627), .Y(n_672) );
A2O1A1Ixp33_ASAP7_75t_SL g673 ( .A1(n_656), .A2(n_287), .B(n_309), .C(n_344), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_641), .A2(n_247), .A3(n_308), .B1(n_309), .B2(n_344), .C1(n_348), .C2(n_660), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_644), .B(n_308), .Y(n_675) );
INVxp67_ASAP7_75t_L g676 ( .A(n_649), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_653), .B(n_308), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_642), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_639), .B(n_308), .Y(n_679) );
INVx1_ASAP7_75t_SL g680 ( .A(n_645), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_648), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_657), .Y(n_682) );
AO22x2_ASAP7_75t_L g683 ( .A1(n_635), .A2(n_348), .B1(n_344), .B2(n_247), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_646), .Y(n_684) );
INVx2_ASAP7_75t_SL g685 ( .A(n_680), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_669), .A2(n_659), .B1(n_652), .B2(n_633), .C(n_643), .Y(n_686) );
NOR2xp33_ASAP7_75t_R g687 ( .A(n_672), .B(n_651), .Y(n_687) );
AOI211xp5_ASAP7_75t_L g688 ( .A1(n_670), .A2(n_645), .B(n_638), .C(n_658), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_683), .A2(n_635), .B1(n_640), .B2(n_636), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_683), .A2(n_636), .B(n_665), .Y(n_690) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_676), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_681), .A2(n_662), .B1(n_637), .B2(n_634), .C(n_638), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_667), .A2(n_671), .B1(n_665), .B2(n_674), .C(n_673), .Y(n_693) );
XNOR2xp5_ASAP7_75t_L g694 ( .A(n_683), .B(n_650), .Y(n_694) );
NOR2xp33_ASAP7_75t_R g695 ( .A(n_675), .B(n_656), .Y(n_695) );
OR2x6_ASAP7_75t_L g696 ( .A(n_675), .B(n_636), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_684), .B(n_634), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_682), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_666), .A2(n_647), .B1(n_650), .B2(n_661), .Y(n_699) );
INVx1_ASAP7_75t_SL g700 ( .A(n_677), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_678), .Y(n_701) );
NAND3xp33_ASAP7_75t_SL g702 ( .A(n_673), .B(n_344), .C(n_348), .Y(n_702) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_668), .A2(n_344), .B(n_348), .C(n_247), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_671), .B(n_667), .C(n_670), .D(n_669), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_679), .B(n_667), .C(n_670), .D(n_669), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_686), .B(n_705), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g707 ( .A(n_685), .Y(n_707) );
NAND2x1p5_ASAP7_75t_L g708 ( .A(n_690), .B(n_689), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_687), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_688), .B(n_700), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_708), .A2(n_704), .B1(n_693), .B2(n_696), .C(n_692), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_707), .Y(n_712) );
NOR4xp75_ASAP7_75t_L g713 ( .A(n_706), .B(n_699), .C(n_702), .D(n_697), .Y(n_713) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_712), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_711), .Y(n_715) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_708), .B1(n_709), .B2(n_707), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_714), .Y(n_717) );
AOI222xp33_ASAP7_75t_L g718 ( .A1(n_717), .A2(n_716), .B1(n_710), .B2(n_713), .C1(n_691), .C2(n_694), .Y(n_718) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_718), .A2(n_703), .B1(n_695), .B2(n_698), .C(n_701), .Y(n_719) );
endmodule