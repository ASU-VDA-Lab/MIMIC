module fake_jpeg_12970_n_40 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_40);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_17),
.B1(n_16),
.B2(n_7),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g25 ( 
.A(n_20),
.B(n_0),
.Y(n_25)
);

XNOR2x2_ASAP7_75t_SL g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_29),
.B(n_32),
.Y(n_34)
);

AO21x1_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_31),
.B(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_26),
.C(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_35),
.C(n_16),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_2),
.B(n_3),
.Y(n_37)
);

OA21x2_ASAP7_75t_SL g39 ( 
.A1(n_38),
.A2(n_37),
.B(n_6),
.Y(n_39)
);

O2A1O1Ixp33_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_4),
.B(n_8),
.C(n_9),
.Y(n_40)
);


endmodule