module fake_jpeg_14363_n_29 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_29);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_29;

wire n_13;
wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_15;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

OR2x2_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_9),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_5),
.B(n_6),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_12),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_17),
.Y(n_20)
);

OR2x4_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_18),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_21),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_24),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_20),
.A2(n_11),
.B1(n_14),
.B2(n_13),
.Y(n_24)
);

NOR3xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_11),
.C(n_2),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_24),
.B(n_25),
.Y(n_27)
);

OAI211xp5_ASAP7_75t_L g28 ( 
.A1(n_27),
.A2(n_1),
.B(n_3),
.C(n_7),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_10),
.Y(n_29)
);


endmodule