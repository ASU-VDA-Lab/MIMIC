module fake_jpeg_31541_n_443 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_443);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_443;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_46),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_48),
.B(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_58),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx4f_ASAP7_75t_SL g101 ( 
.A(n_59),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_60),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_20),
.B(n_9),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_80),
.Y(n_108)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_66),
.Y(n_109)
);

BUFx4f_ASAP7_75t_SL g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

BUFx12_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx4f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_81),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_78),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_24),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_79),
.B(n_44),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_24),
.B(n_10),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_19),
.B1(n_29),
.B2(n_37),
.Y(n_102)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_89),
.Y(n_135)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_36),
.B(n_43),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_92),
.Y(n_145)
);

OR2x4_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_43),
.Y(n_92)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_67),
.Y(n_100)
);

INVx13_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_28),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_58),
.A2(n_25),
.B1(n_37),
.B2(n_19),
.Y(n_119)
);

BUFx10_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_25),
.B1(n_37),
.B2(n_19),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_60),
.Y(n_125)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_54),
.B(n_25),
.C(n_44),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_78),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_59),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_129),
.B(n_59),
.Y(n_143)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_96),
.Y(n_138)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_101),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_141),
.B(n_143),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_28),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_144),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_136),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_147),
.Y(n_189)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_132),
.Y(n_148)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_155),
.Y(n_184)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_108),
.B(n_31),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_172),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_153),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_104),
.Y(n_154)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_76),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_156),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_73),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_157),
.B(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_158),
.Y(n_183)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_160),
.Y(n_198)
);

BUFx12f_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_162),
.Y(n_200)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_178)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

BUFx12_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_171),
.B1(n_173),
.B2(n_122),
.Y(n_196)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_101),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_135),
.B(n_23),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_102),
.B1(n_120),
.B2(n_119),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_192),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_168),
.A2(n_117),
.B1(n_128),
.B2(n_90),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_182),
.B1(n_122),
.B2(n_139),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_171),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_161),
.A2(n_128),
.B1(n_95),
.B2(n_111),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_145),
.B(n_23),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_31),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_167),
.A2(n_65),
.B1(n_57),
.B2(n_75),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_95),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_163),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_111),
.B1(n_118),
.B2(n_68),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_197),
.A2(n_126),
.B1(n_105),
.B2(n_118),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_204),
.Y(n_230)
);

OA22x2_ASAP7_75t_L g205 ( 
.A1(n_197),
.A2(n_167),
.B1(n_87),
.B2(n_150),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_206),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_195),
.B(n_167),
.Y(n_206)
);

NAND2x1_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_175),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_226),
.Y(n_242)
);

AND2x6_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_152),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_208),
.A2(n_180),
.B(n_199),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_145),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_183),
.C(n_174),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_211),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_202),
.B(n_18),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_137),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_216),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_185),
.B1(n_153),
.B2(n_170),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_140),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_221),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_180),
.Y(n_218)
);

INVx13_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_189),
.Y(n_219)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_137),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_152),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_165),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_22),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_224),
.Y(n_236)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_225),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_201),
.B(n_16),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_22),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_192),
.B1(n_185),
.B2(n_126),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_231),
.A2(n_232),
.B1(n_233),
.B2(n_253),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_206),
.A2(n_185),
.B1(n_105),
.B2(n_50),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_212),
.A2(n_205),
.B1(n_207),
.B2(n_216),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_209),
.B(n_199),
.C(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_237),
.B(n_252),
.C(n_217),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_243),
.A2(n_222),
.B(n_213),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_215),
.A2(n_212),
.B1(n_207),
.B2(n_205),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_209),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_187),
.B1(n_177),
.B2(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_207),
.B(n_188),
.C(n_174),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_154),
.B1(n_187),
.B2(n_84),
.Y(n_253)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_35),
.A3(n_94),
.B1(n_194),
.B2(n_130),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_254),
.A2(n_204),
.B(n_223),
.Y(n_259)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_255),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_256),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_269),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_226),
.B1(n_225),
.B2(n_194),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_258),
.A2(n_156),
.B1(n_244),
.B2(n_171),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_259),
.B(n_263),
.Y(n_309)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_276),
.B1(n_278),
.B2(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_210),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_221),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_267),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_208),
.B(n_212),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_265),
.A2(n_277),
.B(n_237),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_211),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_233),
.A2(n_214),
.B1(n_205),
.B2(n_218),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_270),
.A2(n_249),
.B1(n_214),
.B2(n_239),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_228),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_251),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_227),
.Y(n_273)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_238),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_281),
.Y(n_287)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_205),
.C(n_200),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_252),
.C(n_247),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_203),
.Y(n_280)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_280),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_238),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_234),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_236),
.B(n_224),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g307 ( 
.A1(n_283),
.A2(n_229),
.B(n_284),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_245),
.B(n_243),
.Y(n_284)
);

O2A1O1Ixp33_ASAP7_75t_L g285 ( 
.A1(n_262),
.A2(n_242),
.B(n_245),
.C(n_235),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_285),
.A2(n_265),
.B(n_277),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_298),
.C(n_306),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_273),
.B(n_240),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_281),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_230),
.Y(n_291)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_292),
.B(n_259),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_307),
.B1(n_278),
.B2(n_256),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_240),
.Y(n_294)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_294),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_296),
.A2(n_312),
.B1(n_280),
.B2(n_255),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_242),
.C(n_254),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_262),
.A2(n_205),
.B(n_200),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_303),
.A2(n_260),
.B(n_106),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_232),
.Y(n_305)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_305),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_231),
.C(n_198),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_310),
.B1(n_276),
.B2(n_268),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_229),
.B1(n_239),
.B2(n_179),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_257),
.B(n_198),
.C(n_179),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_266),
.C(n_268),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_282),
.A2(n_47),
.B1(n_72),
.B2(n_69),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_314),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_337),
.B1(n_300),
.B2(n_312),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_316),
.B(n_329),
.Y(n_351)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_317),
.Y(n_358)
);

AO21x1_ASAP7_75t_L g352 ( 
.A1(n_320),
.A2(n_332),
.B(n_291),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_321),
.A2(n_333),
.B(n_301),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_279),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_322),
.B(n_324),
.C(n_325),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_266),
.C(n_280),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_327),
.A2(n_328),
.B1(n_323),
.B2(n_333),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_328),
.A2(n_285),
.B(n_304),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_107),
.C(n_219),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_40),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g360 ( 
.A(n_330),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_311),
.B(n_107),
.C(n_219),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_289),
.B(n_14),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_303),
.A2(n_97),
.B(n_17),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_294),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_334),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_299),
.B(n_40),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_336),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_308),
.A2(n_35),
.B1(n_29),
.B2(n_99),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_166),
.C(n_162),
.Y(n_338)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_339),
.A2(n_345),
.B1(n_340),
.B2(n_343),
.Y(n_373)
);

AO21x1_ASAP7_75t_L g362 ( 
.A1(n_343),
.A2(n_348),
.B(n_352),
.Y(n_362)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_319),
.Y(n_344)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_327),
.A2(n_313),
.B1(n_309),
.B2(n_301),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_349),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_325),
.A2(n_298),
.B(n_313),
.Y(n_353)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_353),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_289),
.B1(n_300),
.B2(n_305),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_357),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_320),
.A2(n_292),
.B(n_287),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_356),
.A2(n_322),
.B(n_332),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_287),
.B1(n_297),
.B2(n_286),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_326),
.A2(n_297),
.B1(n_286),
.B2(n_302),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_317),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_324),
.A2(n_83),
.B1(n_62),
.B2(n_51),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_344),
.Y(n_363)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_342),
.A2(n_316),
.B1(n_329),
.B2(n_338),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_352),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_318),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_365),
.A2(n_376),
.B(n_377),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_367),
.B(n_369),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_375),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_331),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_318),
.C(n_7),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_371),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_346),
.A2(n_45),
.B1(n_13),
.B2(n_15),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g394 ( 
.A(n_373),
.B(n_358),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_166),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_374),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_346),
.B(n_162),
.Y(n_375)
);

NAND2x1_ASAP7_75t_SL g376 ( 
.A(n_350),
.B(n_160),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_339),
.A2(n_45),
.B1(n_16),
.B2(n_18),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_350),
.B(n_342),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_378),
.A2(n_345),
.B1(n_351),
.B2(n_358),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_347),
.C(n_341),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_384),
.C(n_372),
.Y(n_401)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_383),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_347),
.C(n_353),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_388),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_373),
.B(n_361),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_348),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_394),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_340),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_391),
.B(n_395),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_362),
.B(n_160),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_384),
.B(n_380),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_400),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_376),
.Y(n_399)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_399),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_380),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_401),
.B(n_403),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_396),
.A2(n_379),
.B1(n_381),
.B2(n_363),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_386),
.B(n_362),
.Y(n_405)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_393),
.A2(n_368),
.B1(n_131),
.B2(n_123),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_407),
.B(n_408),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_382),
.A2(n_131),
.B1(n_123),
.B2(n_45),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_392),
.B(n_123),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_55),
.Y(n_415)
);

A2O1A1Ixp33_ASAP7_75t_SL g411 ( 
.A1(n_406),
.A2(n_394),
.B(n_388),
.C(n_389),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_413),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_404),
.A2(n_385),
.B1(n_18),
.B2(n_8),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_415),
.B(n_417),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_13),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_13),
.B1(n_17),
.B2(n_8),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_418),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_406),
.B(n_17),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_420),
.A2(n_409),
.B(n_8),
.Y(n_423)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_412),
.A2(n_402),
.B(n_7),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_424),
.A2(n_425),
.B(n_426),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_419),
.A2(n_402),
.B(n_1),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_416),
.A2(n_131),
.B(n_114),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_410),
.A2(n_0),
.B(n_1),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_427),
.B(n_0),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g429 ( 
.A(n_428),
.Y(n_429)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_429),
.A2(n_434),
.A3(n_114),
.B1(n_64),
.B2(n_19),
.C1(n_73),
.C2(n_46),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_411),
.C(n_414),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_431),
.A2(n_432),
.B(n_433),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_411),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_435),
.Y(n_438)
);

AOI322xp5_ASAP7_75t_L g436 ( 
.A1(n_430),
.A2(n_64),
.A3(n_46),
.B1(n_3),
.B2(n_4),
.C1(n_2),
.C2(n_0),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_436),
.A2(n_437),
.B(n_0),
.Y(n_439)
);

AOI21x1_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_438),
.B(n_3),
.Y(n_440)
);

NAND3xp33_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_2),
.C(n_4),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_441),
.A2(n_4),
.B(n_46),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_442),
.B(n_4),
.Y(n_443)
);


endmodule