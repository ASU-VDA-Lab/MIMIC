module fake_jpeg_27887_n_328 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_47),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_31),
.Y(n_48)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_48),
.B(n_65),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_56),
.Y(n_80)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_46),
.A2(n_17),
.B1(n_27),
.B2(n_21),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_62),
.B1(n_75),
.B2(n_42),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_17),
.B1(n_27),
.B2(n_30),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_59),
.A2(n_20),
.B1(n_36),
.B2(n_38),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_27),
.B1(n_17),
.B2(n_34),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_18),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_76),
.B(n_35),
.C(n_22),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_35),
.B1(n_23),
.B2(n_22),
.Y(n_116)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_81),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_74),
.B(n_41),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_83),
.B(n_97),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_89),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_41),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_107),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_56),
.A2(n_42),
.B1(n_45),
.B2(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_104),
.B1(n_112),
.B2(n_116),
.Y(n_123)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_51),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_91),
.Y(n_136)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_49),
.A2(n_42),
.B1(n_37),
.B2(n_38),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_93),
.A2(n_106),
.B1(n_69),
.B2(n_72),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_102),
.B1(n_111),
.B2(n_112),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_98),
.B(n_103),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_28),
.B1(n_34),
.B2(n_30),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_66),
.A2(n_33),
.B1(n_25),
.B2(n_28),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_100),
.Y(n_132)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_20),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_60),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_49),
.A2(n_45),
.B1(n_41),
.B2(n_33),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_50),
.B(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_57),
.B(n_33),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_60),
.A2(n_45),
.B1(n_35),
.B2(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_57),
.B(n_25),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_61),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_118),
.A2(n_119),
.B1(n_121),
.B2(n_133),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_60),
.B1(n_69),
.B2(n_55),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_68),
.C(n_73),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_141),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_67),
.B1(n_72),
.B2(n_61),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_124),
.A2(n_111),
.B1(n_106),
.B2(n_89),
.Y(n_160)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_78),
.A2(n_72),
.B1(n_61),
.B2(n_29),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_81),
.B(n_96),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_140),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_116),
.A2(n_29),
.B1(n_24),
.B2(n_22),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_29),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_29),
.C(n_24),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_108),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_80),
.A2(n_24),
.B1(n_26),
.B2(n_8),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_80),
.A2(n_26),
.B1(n_7),
.B2(n_9),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_87),
.A2(n_26),
.B1(n_7),
.B2(n_9),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

A2O1A1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_94),
.B(n_103),
.C(n_87),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_148),
.A2(n_142),
.B(n_139),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_131),
.B(n_94),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_152),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_150),
.B(n_153),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_114),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_156),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_159),
.Y(n_208)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_132),
.B1(n_122),
.B2(n_145),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_163),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_135),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_162),
.Y(n_203)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_165),
.Y(n_185)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_128),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_166),
.B(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_117),
.B(n_77),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_118),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_178),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_126),
.A2(n_109),
.B(n_101),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_179),
.B(n_139),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_77),
.Y(n_175)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_79),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_136),
.B(n_79),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_173),
.A2(n_124),
.B1(n_123),
.B2(n_132),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_182),
.A2(n_195),
.B1(n_172),
.B2(n_154),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_120),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_184),
.C(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_120),
.C(n_136),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_188),
.A2(n_189),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_159),
.B(n_167),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_141),
.C(n_122),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_152),
.B(n_144),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_200),
.C(n_206),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_161),
.A2(n_123),
.B(n_127),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_179),
.B(n_155),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_137),
.B1(n_93),
.B2(n_86),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_199),
.B(n_176),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_142),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_201),
.B(n_0),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_147),
.Y(n_202)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_168),
.A2(n_86),
.B1(n_105),
.B2(n_115),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_204),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_151),
.B(n_113),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_163),
.A2(n_86),
.B1(n_98),
.B2(n_84),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_211),
.A2(n_170),
.B1(n_204),
.B2(n_178),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_148),
.C(n_149),
.Y(n_215)
);

AOI321xp33_ASAP7_75t_L g250 ( 
.A1(n_215),
.A2(n_222),
.A3(n_181),
.B1(n_10),
.B2(n_14),
.C(n_13),
.Y(n_250)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_185),
.Y(n_217)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_166),
.Y(n_219)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_220),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_190),
.B(n_165),
.Y(n_221)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_156),
.C(n_162),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_235),
.B(n_238),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_224),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_170),
.B1(n_157),
.B2(n_176),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_234),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_187),
.C(n_180),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_196),
.B(n_211),
.Y(n_249)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_147),
.A3(n_169),
.B1(n_134),
.B2(n_113),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_182),
.A2(n_110),
.B1(n_82),
.B2(n_9),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_82),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_110),
.B1(n_6),
.B2(n_10),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_194),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_237),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_198),
.B(n_6),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_209),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_183),
.C(n_184),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_242),
.C(n_244),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_200),
.C(n_191),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_206),
.C(n_193),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_189),
.C(n_187),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_246),
.C(n_247),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_192),
.C(n_201),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_188),
.C(n_210),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_230),
.B(n_218),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_235),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_224),
.B(n_181),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_251),
.B(n_226),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_186),
.C(n_14),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_256),
.C(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_186),
.C(n_12),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_11),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_232),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_264),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_276),
.B(n_225),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_258),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_265),
.B(n_269),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_267),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_275),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_245),
.B(n_246),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_233),
.Y(n_273)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_247),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_231),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_243),
.A2(n_213),
.B1(n_214),
.B2(n_234),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_0),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_214),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_264),
.A2(n_213),
.B1(n_255),
.B2(n_239),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_288),
.B(n_0),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_242),
.C(n_244),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_293),
.C(n_1),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_292),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_289),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_272),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_11),
.Y(n_293)
);

INVx6_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_298),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_270),
.Y(n_295)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_295),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_302),
.B(n_1),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_270),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_280),
.B(n_276),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_301),
.Y(n_309)
);

AOI31xp33_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_276),
.A3(n_266),
.B(n_261),
.Y(n_300)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_300),
.A2(n_281),
.B(n_3),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_11),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_5),
.B1(n_2),
.B2(n_3),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_303),
.A2(n_282),
.B1(n_281),
.B2(n_283),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_287),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_313),
.B(n_4),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_311),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_314),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_303),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_294),
.B1(n_297),
.B2(n_305),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_315),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_304),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_318),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_312),
.A2(n_302),
.B(n_4),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_319),
.Y(n_323)
);

NAND4xp25_ASAP7_75t_L g324 ( 
.A(n_317),
.B(n_308),
.C(n_306),
.D(n_309),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_324),
.A2(n_314),
.B(n_5),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_321),
.B(n_320),
.C(n_316),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.B(n_322),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_323),
.Y(n_328)
);


endmodule