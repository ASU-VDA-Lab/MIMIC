module fake_jpeg_3898_n_42 (n_3, n_2, n_1, n_0, n_4, n_5, n_42);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_42;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx6_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx5p33_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_19),
.B1(n_15),
.B2(n_21),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_11),
.A2(n_0),
.B(n_13),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_22),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_9),
.Y(n_21)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.C(n_27),
.Y(n_34)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_25),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_34),
.Y(n_36)
);

OAI321xp33_ASAP7_75t_L g37 ( 
.A1(n_33),
.A2(n_24),
.A3(n_17),
.B1(n_22),
.B2(n_26),
.C(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_26),
.B1(n_30),
.B2(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_38),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_14),
.C(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_39),
.Y(n_42)
);


endmodule