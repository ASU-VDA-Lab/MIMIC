module fake_jpeg_8784_n_169 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_41),
.Y(n_44)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_R g34 ( 
.A(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_28),
.B1(n_23),
.B2(n_31),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_21),
.B1(n_26),
.B2(n_22),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_25),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_16),
.Y(n_55)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_16),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_15),
.B1(n_23),
.B2(n_31),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_24),
.B1(n_27),
.B2(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_62),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_32),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_43),
.B1(n_15),
.B2(n_21),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_66),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_60),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_51),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_73),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_36),
.C(n_35),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_74),
.B(n_85),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_22),
.B1(n_17),
.B2(n_25),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_79),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_52),
.B(n_55),
.Y(n_79)
);

INVx5_ASAP7_75t_SL g81 ( 
.A(n_50),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

O2A1O1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_42),
.B(n_27),
.C(n_18),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_84),
.A2(n_87),
.B(n_27),
.Y(n_105)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_1),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_42),
.B1(n_24),
.B2(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_58),
.B1(n_54),
.B2(n_46),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_94),
.B1(n_102),
.B2(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_58),
.B1(n_48),
.B2(n_45),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_44),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_64),
.B(n_35),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_58),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_74),
.B1(n_64),
.B2(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_82),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_79),
.B(n_11),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_13),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_109),
.A2(n_120),
.B1(n_113),
.B2(n_89),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_113),
.Y(n_126)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_103),
.A2(n_85),
.B(n_73),
.C(n_80),
.D(n_36),
.Y(n_111)
);

NOR4xp25_ASAP7_75t_L g132 ( 
.A(n_111),
.B(n_101),
.C(n_106),
.D(n_12),
.Y(n_132)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_117),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_115),
.B(n_121),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_73),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_92),
.C(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_122),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_48),
.B1(n_86),
.B2(n_63),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_10),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_128),
.B1(n_133),
.B2(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_89),
.B1(n_105),
.B2(n_90),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_112),
.A2(n_93),
.B(n_95),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_129),
.B(n_108),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_130),
.B(n_131),
.C(n_110),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_93),
.C(n_91),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_132),
.B(n_111),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_97),
.B1(n_91),
.B2(n_61),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_9),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_135),
.B(n_10),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_137),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_124),
.B(n_83),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_107),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_129),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_107),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_144),
.A2(n_145),
.B1(n_143),
.B2(n_131),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_147),
.A2(n_151),
.B(n_9),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_140),
.A2(n_142),
.B1(n_139),
.B2(n_137),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_152),
.A2(n_153),
.B1(n_148),
.B2(n_150),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_141),
.A2(n_77),
.B1(n_72),
.B2(n_18),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_151),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_157),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_147),
.A2(n_1),
.B(n_2),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_2),
.C(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_152),
.B1(n_3),
.B2(n_6),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_159),
.B(n_161),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_8),
.B(n_6),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_160),
.C(n_7),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_161),
.B(n_155),
.Y(n_163)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_163),
.Y(n_167)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_7),
.B(n_8),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_164),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_167),
.Y(n_169)
);


endmodule