module real_aes_13169_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_923, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_923;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_905;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_860;
wire n_781;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_898;
wire n_115;
wire n_604;
wire n_110;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g190 ( .A(n_0), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_1), .Y(n_259) );
OA21x2_ASAP7_75t_L g138 ( .A1(n_2), .A2(n_49), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g198 ( .A(n_2), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_3), .B(n_187), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_4), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_5), .B(n_620), .Y(n_678) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_6), .B(n_149), .Y(n_591) );
AND2x2_ASAP7_75t_L g331 ( .A(n_7), .B(n_136), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_8), .B(n_148), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_9), .B(n_295), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_10), .B(n_295), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_11), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_12), .B(n_180), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_13), .B(n_235), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_14), .B(n_189), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_15), .Y(n_609) );
BUFx3_ASAP7_75t_L g146 ( .A(n_16), .Y(n_146) );
INVx1_ASAP7_75t_L g151 ( .A(n_16), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_17), .B(n_135), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_18), .B(n_322), .Y(n_658) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_19), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_20), .A2(n_124), .B1(n_911), .B2(n_912), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_20), .Y(n_911) );
BUFx10_ASAP7_75t_L g120 ( .A(n_21), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g654 ( .A(n_22), .B(n_216), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_23), .Y(n_603) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_24), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_25), .B(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g217 ( .A(n_26), .B(n_212), .C(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_27), .B(n_216), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_28), .B(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_29), .B(n_322), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_30), .Y(n_915) );
NAND2xp33_ASAP7_75t_L g681 ( .A(n_31), .B(n_176), .Y(n_681) );
INVx1_ASAP7_75t_L g169 ( .A(n_32), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_33), .A2(n_264), .B(n_324), .C(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_34), .B(n_179), .Y(n_178) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_35), .A2(n_100), .B1(n_113), .B2(n_920), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_36), .B(n_261), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_37), .B(n_187), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_38), .B(n_279), .Y(n_625) );
AND3x2_ASAP7_75t_L g108 ( .A(n_39), .B(n_109), .C(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g554 ( .A(n_39), .Y(n_554) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_40), .B(n_297), .Y(n_296) );
AO221x1_ASAP7_75t_L g661 ( .A1(n_41), .A2(n_82), .B1(n_175), .B2(n_216), .C(n_278), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_42), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_43), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g168 ( .A(n_44), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_45), .B(n_135), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_46), .B(n_164), .Y(n_184) );
NAND3xp33_ASAP7_75t_L g643 ( .A(n_47), .B(n_263), .C(n_264), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_48), .B(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g197 ( .A(n_49), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g328 ( .A(n_50), .Y(n_328) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_51), .A2(n_186), .B(n_188), .C(n_191), .Y(n_185) );
INVx1_ASAP7_75t_L g139 ( .A(n_52), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g565 ( .A1(n_53), .A2(n_566), .B(n_568), .C(n_570), .Y(n_565) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_54), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_55), .B(n_135), .Y(n_265) );
INVx2_ASAP7_75t_L g569 ( .A(n_56), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_57), .B(n_164), .Y(n_593) );
AND2x4_ASAP7_75t_L g106 ( .A(n_58), .B(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g245 ( .A(n_59), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g917 ( .A(n_60), .Y(n_917) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_61), .B(n_73), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_62), .B(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g107 ( .A(n_63), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_64), .B(n_143), .Y(n_159) );
INVx1_ASAP7_75t_L g277 ( .A(n_65), .Y(n_277) );
AND2x2_ASAP7_75t_L g627 ( .A(n_66), .B(n_164), .Y(n_627) );
INVx1_ASAP7_75t_L g666 ( .A(n_67), .Y(n_666) );
INVx2_ASAP7_75t_L g110 ( .A(n_68), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_69), .B(n_207), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_70), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_71), .B(n_218), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_72), .A2(n_75), .B1(n_575), .B2(n_620), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_74), .B(n_264), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_76), .A2(n_122), .B1(n_123), .B2(n_897), .Y(n_121) );
INVx1_ASAP7_75t_L g897 ( .A(n_76), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_77), .B(n_215), .Y(n_301) );
INVx1_ASAP7_75t_L g177 ( .A(n_78), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_79), .B(n_283), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_80), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_81), .B(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g577 ( .A(n_83), .B(n_136), .Y(n_577) );
INVx1_ASAP7_75t_L g154 ( .A(n_84), .Y(n_154) );
INVx1_ASAP7_75t_L g193 ( .A(n_84), .Y(n_193) );
BUFx3_ASAP7_75t_L g235 ( .A(n_84), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_85), .B(n_207), .Y(n_256) );
INVx1_ASAP7_75t_L g243 ( .A(n_86), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_87), .B(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_88), .B(n_195), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g299 ( .A(n_89), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_90), .B(n_136), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_91), .B(n_588), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_92), .B(n_164), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_93), .B(n_157), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_94), .Y(n_238) );
INVx1_ASAP7_75t_L g233 ( .A(n_95), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_96), .Y(n_645) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_97), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_98), .B(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
BUFx12f_ASAP7_75t_SL g921 ( .A(n_101), .Y(n_921) );
AND2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_108), .B(n_120), .Y(n_919) );
AND2x2_ASAP7_75t_L g118 ( .A(n_109), .B(n_111), .Y(n_118) );
BUFx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g908 ( .A(n_110), .Y(n_908) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_112), .B(n_554), .Y(n_909) );
OR2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_914), .Y(n_113) );
OAI21xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B(n_898), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
CKINVDCx11_ASAP7_75t_R g900 ( .A(n_120), .Y(n_900) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_549), .B1(n_555), .B2(n_895), .Y(n_123) );
INVx3_ASAP7_75t_L g912 ( .A(n_124), .Y(n_912) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_454), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_390), .C(n_425), .Y(n_125) );
NAND3xp33_ASAP7_75t_SL g126 ( .A(n_127), .B(n_332), .C(n_362), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_222), .B1(n_286), .B2(n_308), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_129), .B(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_170), .Y(n_129) );
AND2x2_ASAP7_75t_L g470 ( .A(n_130), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_130), .B(n_417), .Y(n_483) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_131), .B(n_267), .C(n_371), .Y(n_449) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g335 ( .A(n_132), .B(n_288), .Y(n_335) );
INVx2_ASAP7_75t_L g366 ( .A(n_132), .Y(n_366) );
OR2x2_ASAP7_75t_L g389 ( .A(n_132), .B(n_365), .Y(n_389) );
AND2x2_ASAP7_75t_L g405 ( .A(n_132), .B(n_201), .Y(n_405) );
BUFx2_ASAP7_75t_L g459 ( .A(n_132), .Y(n_459) );
AND2x4_ASAP7_75t_L g467 ( .A(n_132), .B(n_424), .Y(n_467) );
INVx2_ASAP7_75t_L g477 ( .A(n_132), .Y(n_477) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2x1_ASAP7_75t_L g133 ( .A(n_134), .B(n_140), .Y(n_133) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_135), .Y(n_307) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_138), .Y(n_164) );
BUFx2_ASAP7_75t_L g252 ( .A(n_138), .Y(n_252) );
INVx1_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
OAI21x1_ASAP7_75t_SL g140 ( .A1(n_141), .A2(n_155), .B(n_162), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_152), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_143), .A2(n_242), .B1(n_244), .B2(n_246), .Y(n_241) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_144), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
INVx1_ASAP7_75t_L g283 ( .A(n_145), .Y(n_283) );
INVx2_ASAP7_75t_L g575 ( .A(n_145), .Y(n_575) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx2_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx2_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVx2_ASAP7_75t_L g263 ( .A(n_150), .Y(n_263) );
INVx1_ASAP7_75t_L g567 ( .A(n_150), .Y(n_567) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_152), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_152), .B(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g240 ( .A(n_153), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_153), .A2(n_677), .B(n_678), .Y(n_676) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx3_ASAP7_75t_L g161 ( .A(n_154), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .B(n_160), .Y(n_155) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_161), .A2(n_294), .B(n_296), .Y(n_293) );
INVx1_ASAP7_75t_L g570 ( .A(n_161), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_161), .A2(n_680), .B(n_681), .Y(n_679) );
NOR2x1_ASAP7_75t_SL g162 ( .A(n_163), .B(n_165), .Y(n_162) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_163), .Y(n_291) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g203 ( .A(n_164), .Y(n_203) );
INVx2_ASAP7_75t_L g617 ( .A(n_164), .Y(n_617) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_164), .Y(n_651) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_164), .B(n_236), .Y(n_659) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_166), .B(n_196), .Y(n_599) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g220 ( .A(n_167), .Y(n_220) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g200 ( .A(n_168), .Y(n_200) );
INVx3_ASAP7_75t_L g236 ( .A(n_168), .Y(n_236) );
BUFx6f_ASAP7_75t_SL g284 ( .A(n_168), .Y(n_284) );
OR2x2_ASAP7_75t_L g462 ( .A(n_170), .B(n_341), .Y(n_462) );
INVx2_ASAP7_75t_L g520 ( .A(n_170), .Y(n_520) );
OR2x2_ASAP7_75t_SL g170 ( .A(n_171), .B(n_201), .Y(n_170) );
OR2x6_ASAP7_75t_L g303 ( .A(n_171), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g342 ( .A(n_171), .Y(n_342) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g338 ( .A(n_172), .Y(n_338) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_183), .B(n_194), .Y(n_172) );
AOI21x1_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_178), .B(n_182), .Y(n_173) );
OR2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_177), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g207 ( .A(n_176), .Y(n_207) );
INVx2_ASAP7_75t_L g261 ( .A(n_176), .Y(n_261) );
INVx2_ASAP7_75t_L g273 ( .A(n_176), .Y(n_273) );
INVx2_ASAP7_75t_L g295 ( .A(n_176), .Y(n_295) );
INVx3_ASAP7_75t_L g322 ( .A(n_176), .Y(n_322) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
INVx2_ASAP7_75t_L g297 ( .A(n_180), .Y(n_297) );
INVx2_ASAP7_75t_L g300 ( .A(n_180), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_180), .B(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
AOI22x1_ASAP7_75t_L g319 ( .A1(n_182), .A2(n_192), .B1(n_320), .B2(n_326), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_185), .Y(n_183) );
OAI21xp33_ASAP7_75t_L g194 ( .A1(n_184), .A2(n_195), .B(n_200), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_186), .A2(n_327), .B1(n_328), .B2(n_329), .Y(n_326) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
AOI21x1_ASAP7_75t_L g205 ( .A1(n_192), .A2(n_206), .B(n_208), .Y(n_205) );
AOI21xp5_ASAP7_75t_SL g618 ( .A1(n_192), .A2(n_619), .B(n_621), .Y(n_618) );
BUFx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g213 ( .A(n_193), .Y(n_213) );
INVxp67_ASAP7_75t_L g353 ( .A(n_195), .Y(n_353) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_196) );
AOI21x1_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_198), .B(n_199), .Y(n_229) );
INVx1_ASAP7_75t_L g355 ( .A(n_200), .Y(n_355) );
AND2x2_ASAP7_75t_L g471 ( .A(n_201), .B(n_338), .Y(n_471) );
OA21x2_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_221), .Y(n_201) );
OA21x2_ASAP7_75t_L g674 ( .A1(n_202), .A2(n_675), .B(n_682), .Y(n_674) );
INVx1_ASAP7_75t_SL g202 ( .A(n_203), .Y(n_202) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_204), .A2(n_221), .B(n_307), .Y(n_306) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_210), .B(n_220), .Y(n_204) );
O2A1O1Ixp5_ASAP7_75t_L g585 ( .A1(n_209), .A2(n_586), .B(n_587), .C(n_589), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_217), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
BUFx10_ASAP7_75t_L g257 ( .A(n_213), .Y(n_257) );
INVxp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_216), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g246 ( .A(n_216), .Y(n_246) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g279 ( .A(n_219), .Y(n_279) );
INVx2_ASAP7_75t_L g588 ( .A(n_219), .Y(n_588) );
INVx2_ASAP7_75t_L g620 ( .A(n_219), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_220), .A2(n_254), .B(n_258), .Y(n_253) );
AND2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_266), .Y(n_222) );
AND2x2_ASAP7_75t_L g442 ( .A(n_223), .B(n_372), .Y(n_442) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g495 ( .A(n_224), .Y(n_495) );
AND2x2_ASAP7_75t_L g543 ( .A(n_224), .B(n_382), .Y(n_543) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_249), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_226), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g377 ( .A(n_226), .B(n_378), .Y(n_377) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_247), .Y(n_226) );
AO21x2_ASAP7_75t_L g348 ( .A1(n_227), .A2(n_230), .B(n_247), .Y(n_348) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NOR2xp33_ASAP7_75t_SL g247 ( .A(n_228), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_228), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_R g664 ( .A(n_229), .B(n_236), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_241), .Y(n_230) );
AOI22xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_234), .B1(n_237), .B2(n_239), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NOR3xp33_ASAP7_75t_L g242 ( .A(n_235), .B(n_236), .C(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g264 ( .A(n_235), .Y(n_264) );
INVx2_ASAP7_75t_L g278 ( .A(n_235), .Y(n_278) );
INVx1_ASAP7_75t_L g589 ( .A(n_235), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_236), .B(n_240), .Y(n_239) );
NOR3xp33_ASAP7_75t_L g244 ( .A(n_236), .B(n_240), .C(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g580 ( .A(n_236), .Y(n_580) );
INVx2_ASAP7_75t_L g314 ( .A(n_249), .Y(n_314) );
INVx3_ASAP7_75t_L g356 ( .A(n_249), .Y(n_356) );
INVx1_ASAP7_75t_L g371 ( .A(n_249), .Y(n_371) );
AND2x2_ASAP7_75t_L g376 ( .A(n_249), .B(n_318), .Y(n_376) );
INVx3_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_253), .B(n_265), .Y(n_250) );
OAI21x1_ASAP7_75t_L g269 ( .A1(n_251), .A2(n_270), .B(n_285), .Y(n_269) );
OAI21x1_ASAP7_75t_L g583 ( .A1(n_251), .A2(n_584), .B(n_593), .Y(n_583) );
BUFx3_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_L g579 ( .A(n_252), .Y(n_579) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_257), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_281), .B(n_282), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_257), .A2(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_L g576 ( .A(n_257), .Y(n_576) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_257), .A2(n_591), .B(n_592), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g624 ( .A1(n_257), .A2(n_625), .B(n_626), .Y(n_624) );
O2A1O1Ixp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_260), .B(n_262), .C(n_264), .Y(n_258) );
OAI21xp5_ASAP7_75t_L g641 ( .A1(n_260), .A2(n_642), .B(n_643), .Y(n_641) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NOR2x1p5_ASAP7_75t_L g349 ( .A(n_266), .B(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g507 ( .A(n_267), .B(n_477), .Y(n_507) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_268), .Y(n_311) );
INVx3_ASAP7_75t_L g361 ( .A(n_268), .Y(n_361) );
INVx2_ASAP7_75t_L g378 ( .A(n_268), .Y(n_378) );
AND2x2_ASAP7_75t_L g384 ( .A(n_268), .B(n_347), .Y(n_384) );
AND2x2_ASAP7_75t_L g407 ( .A(n_268), .B(n_318), .Y(n_407) );
AND2x2_ASAP7_75t_L g436 ( .A(n_268), .B(n_348), .Y(n_436) );
INVx1_ASAP7_75t_L g505 ( .A(n_268), .Y(n_505) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_280), .B(n_284), .Y(n_270) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_272), .A2(n_274), .B(n_275), .Y(n_271) );
INVxp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVxp67_ASAP7_75t_L g327 ( .A(n_273), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_279), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
INVx1_ASAP7_75t_L g610 ( .A(n_278), .Y(n_610) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_284), .A2(n_293), .B(n_298), .Y(n_292) );
OAI21x1_ASAP7_75t_L g584 ( .A1(n_284), .A2(n_585), .B(n_590), .Y(n_584) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_303), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g337 ( .A(n_289), .B(n_338), .Y(n_337) );
BUFx3_ASAP7_75t_L g398 ( .A(n_289), .Y(n_398) );
AND2x4_ASAP7_75t_L g417 ( .A(n_289), .B(n_342), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_289), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_290), .Y(n_539) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_292), .B(n_302), .Y(n_290) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_291), .A2(n_319), .B(n_330), .Y(n_318) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_291), .A2(n_292), .B(n_302), .Y(n_341) );
INVx2_ASAP7_75t_L g324 ( .A(n_300), .Y(n_324) );
OR2x2_ASAP7_75t_L g458 ( .A(n_303), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g512 ( .A(n_303), .B(n_398), .Y(n_512) );
INVx2_ASAP7_75t_SL g530 ( .A(n_303), .Y(n_530) );
AND2x2_ASAP7_75t_L g412 ( .A(n_304), .B(n_341), .Y(n_412) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_305), .Y(n_365) );
INVx2_ASAP7_75t_L g424 ( .A(n_305), .Y(n_424) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_312), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND4xp25_ASAP7_75t_L g546 ( .A(n_311), .B(n_388), .C(n_467), .D(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_313), .B(n_407), .Y(n_541) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_314), .B(n_361), .Y(n_360) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_314), .B(n_396), .Y(n_419) );
NOR2x1_ASAP7_75t_L g498 ( .A(n_314), .B(n_347), .Y(n_498) );
AND2x2_ASAP7_75t_L g418 ( .A(n_315), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g359 ( .A(n_316), .B(n_360), .Y(n_359) );
NOR5xp2_ASAP7_75t_L g448 ( .A(n_317), .B(n_449), .C(n_450), .D(n_452), .E(n_453), .Y(n_448) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g430 ( .A(n_318), .B(n_356), .Y(n_430) );
INVx2_ASAP7_75t_L g352 ( .A(n_319), .Y(n_352) );
OAI22x1_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B1(n_324), .B2(n_325), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_331), .A2(n_352), .A3(n_353), .B(n_354), .Y(n_351) );
AO31x2_ASAP7_75t_L g383 ( .A1(n_331), .A2(n_352), .A3(n_353), .B(n_354), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_343), .B1(n_357), .B2(n_358), .Y(n_332) );
NAND3xp33_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .C(n_339), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g529 ( .A(n_335), .B(n_530), .Y(n_529) );
OR2x2_ASAP7_75t_L g526 ( .A(n_336), .B(n_389), .Y(n_526) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
AND2x2_ASAP7_75t_L g440 ( .A(n_337), .B(n_405), .Y(n_440) );
AND2x2_ASAP7_75t_L g476 ( .A(n_337), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g388 ( .A(n_338), .B(n_341), .Y(n_388) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_338), .Y(n_439) );
INVx1_ASAP7_75t_L g451 ( .A(n_338), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_338), .B(n_424), .Y(n_492) );
OAI22xp33_ASAP7_75t_SL g515 ( .A1(n_339), .A2(n_340), .B1(n_359), .B2(n_428), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_339), .A2(n_374), .B1(n_469), .B2(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g392 ( .A(n_340), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x4_ASAP7_75t_L g479 ( .A(n_341), .B(n_467), .Y(n_479) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g370 ( .A(n_346), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_346), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_347), .B(n_356), .Y(n_409) );
BUFx2_ASAP7_75t_L g452 ( .A(n_347), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_347), .B(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_349), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_415) );
INVx1_ASAP7_75t_L g428 ( .A(n_349), .Y(n_428) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_350), .Y(n_509) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_356), .Y(n_350) );
OR2x2_ASAP7_75t_L g373 ( .A(n_351), .B(n_361), .Y(n_373) );
BUFx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AO21x1_ASAP7_75t_L g456 ( .A1(n_360), .A2(n_457), .B(n_460), .Y(n_456) );
INVx2_ASAP7_75t_L g396 ( .A(n_361), .Y(n_396) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_367), .B1(n_379), .B2(n_385), .Y(n_362) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_364), .B(n_398), .Y(n_518) );
AND2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
BUFx2_ASAP7_75t_L g393 ( .A(n_366), .Y(n_393) );
INVx1_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_374), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_369), .A2(n_535), .B1(n_536), .B2(n_540), .C(n_544), .Y(n_534) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g548 ( .A(n_371), .Y(n_548) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
OR2x2_ASAP7_75t_L g414 ( .A(n_373), .B(n_409), .Y(n_414) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_377), .Y(n_375) );
INVx1_ASAP7_75t_L g401 ( .A(n_376), .Y(n_401) );
AND2x2_ASAP7_75t_L g487 ( .A(n_376), .B(n_436), .Y(n_487) );
AND2x2_ASAP7_75t_L g399 ( .A(n_377), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g464 ( .A(n_377), .B(n_381), .Y(n_464) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_381), .B(n_384), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g435 ( .A(n_382), .B(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g447 ( .A(n_383), .Y(n_447) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_388), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g432 ( .A(n_388), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g443 ( .A(n_388), .Y(n_443) );
NOR2x1_ASAP7_75t_L g465 ( .A(n_388), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g535 ( .A(n_388), .B(n_393), .Y(n_535) );
INVx2_ASAP7_75t_L g473 ( .A(n_389), .Y(n_473) );
OAI211xp5_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_401), .B(n_402), .C(n_415), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_394), .B(n_397), .Y(n_391) );
AND2x2_ASAP7_75t_L g416 ( .A(n_393), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g494 ( .A(n_396), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
OR2x2_ASAP7_75t_L g457 ( .A(n_398), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g421 ( .A(n_400), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_400), .B(n_461), .Y(n_460) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_400), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_406), .B1(n_410), .B2(n_413), .Y(n_402) );
OR2x2_ASAP7_75t_L g537 ( .A(n_404), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g533 ( .A(n_407), .Y(n_533) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g446 ( .A(n_409), .B(n_447), .Y(n_446) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g438 ( .A(n_412), .B(n_439), .Y(n_438) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_413), .A2(n_464), .B1(n_465), .B2(n_468), .C(n_474), .Y(n_463) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_417), .B(n_473), .Y(n_472) );
INVx3_ASAP7_75t_R g508 ( .A(n_417), .Y(n_508) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_423), .Y(n_433) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_424), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_431), .B1(n_434), .B2(n_437), .C(n_441), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_430), .B(n_436), .Y(n_480) );
AND2x2_ASAP7_75t_L g484 ( .A(n_430), .B(n_452), .Y(n_484) );
OAI32xp33_ASAP7_75t_L g501 ( .A1(n_430), .A2(n_462), .A3(n_475), .B1(n_497), .B2(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g522 ( .A(n_430), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_433), .Y(n_444) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221x1_ASAP7_75t_L g524 ( .A1(n_435), .A2(n_525), .B1(n_527), .B2(n_528), .C(n_531), .Y(n_524) );
AND2x2_ASAP7_75t_L g527 ( .A(n_436), .B(n_447), .Y(n_527) );
NOR2xp33_ASAP7_75t_SL g437 ( .A(n_438), .B(n_440), .Y(n_437) );
AOI321xp33_ASAP7_75t_L g441 ( .A1(n_438), .A2(n_442), .A3(n_443), .B1(n_444), .B2(n_445), .C(n_448), .Y(n_441) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g544 ( .A1(n_446), .A2(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_447), .B(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g513 ( .A(n_447), .B(n_504), .Y(n_513) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_499), .Y(n_454) );
NAND3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_463), .C(n_481), .Y(n_455) );
OR2x2_ASAP7_75t_L g545 ( .A(n_459), .B(n_492), .Y(n_545) );
INVx3_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_472), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_471), .B(n_477), .Y(n_510) );
INVx1_ASAP7_75t_L g493 ( .A(n_473), .Y(n_493) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_478), .B(n_480), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g490 ( .A(n_477), .Y(n_490) );
INVx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AOI211xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_485), .C(n_496), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B1(n_493), .B2(n_494), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
HB1xp67_ASAP7_75t_SL g511 ( .A(n_495), .Y(n_511) );
OR2x2_ASAP7_75t_L g532 ( .A(n_495), .B(n_533), .Y(n_532) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_514), .C(n_524), .D(n_534), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .Y(n_500) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_504), .Y(n_523) );
OAI322xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_508), .A3(n_509), .B1(n_510), .B2(n_511), .C1(n_512), .C2(n_513), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_521), .Y(n_517) );
INVx2_ASAP7_75t_SL g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
INVx11_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx8_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_SL g896 ( .A(n_552), .Y(n_896) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND4xp75_ASAP7_75t_L g556 ( .A(n_557), .B(n_794), .C(n_847), .D(n_881), .Y(n_556) );
AND4x1_ASAP7_75t_L g557 ( .A(n_558), .B(n_717), .C(n_750), .D(n_772), .Y(n_557) );
NOR2xp33_ASAP7_75t_SL g558 ( .A(n_559), .B(n_686), .Y(n_558) );
OAI222xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_633), .B1(n_667), .B2(n_670), .C1(n_683), .C2(n_923), .Y(n_559) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_628), .Y(n_560) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_594), .Y(n_561) );
OR2x2_ASAP7_75t_L g667 ( .A(n_562), .B(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_581), .Y(n_562) );
INVx1_ASAP7_75t_L g689 ( .A(n_563), .Y(n_689) );
OR2x2_ASAP7_75t_L g826 ( .A(n_563), .B(n_596), .Y(n_826) );
AND2x2_ASAP7_75t_L g837 ( .A(n_563), .B(n_596), .Y(n_837) );
AND2x2_ASAP7_75t_L g878 ( .A(n_563), .B(n_879), .Y(n_878) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g632 ( .A(n_564), .Y(n_632) );
AND2x2_ASAP7_75t_L g701 ( .A(n_564), .B(n_596), .Y(n_701) );
INVx1_ASAP7_75t_L g715 ( .A(n_564), .Y(n_715) );
OR2x2_ASAP7_75t_L g729 ( .A(n_564), .B(n_614), .Y(n_729) );
AND2x2_ASAP7_75t_L g740 ( .A(n_564), .B(n_613), .Y(n_740) );
AND2x2_ASAP7_75t_L g762 ( .A(n_564), .B(n_612), .Y(n_762) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_565), .A2(n_571), .B(n_578), .Y(n_564) );
NOR2xp67_ASAP7_75t_L g568 ( .A(n_566), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_567), .B(n_607), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B(n_577), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_575), .B(n_603), .Y(n_602) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_577), .A2(n_579), .B(n_580), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_579), .B(n_645), .Y(n_644) );
AND2x4_ASAP7_75t_L g616 ( .A(n_580), .B(n_617), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_580), .A2(n_676), .B(n_679), .Y(n_675) );
AND2x2_ASAP7_75t_L g631 ( .A(n_581), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g690 ( .A(n_581), .B(n_597), .Y(n_690) );
OR2x2_ASAP7_75t_L g725 ( .A(n_581), .B(n_612), .Y(n_725) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g685 ( .A(n_582), .Y(n_685) );
AND2x2_ASAP7_75t_L g705 ( .A(n_582), .B(n_614), .Y(n_705) );
INVx1_ASAP7_75t_L g778 ( .A(n_582), .Y(n_778) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g716 ( .A(n_583), .B(n_614), .Y(n_716) );
INVxp33_ASAP7_75t_L g879 ( .A(n_583), .Y(n_879) );
INVx2_ASAP7_75t_SL g622 ( .A(n_588), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g638 ( .A1(n_589), .A2(n_639), .B(n_640), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g656 ( .A1(n_589), .A2(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_612), .Y(n_594) );
BUFx2_ASAP7_75t_SL g743 ( .A(n_595), .Y(n_743) );
INVx2_ASAP7_75t_L g792 ( .A(n_595), .Y(n_792) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_597), .B(n_715), .Y(n_714) );
AO21x2_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_600), .B(n_604), .Y(n_597) );
AO21x1_ASAP7_75t_SL g669 ( .A1(n_598), .A2(n_600), .B(n_604), .Y(n_669) );
INVxp67_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
OAI21x1_ASAP7_75t_SL g604 ( .A1(n_599), .A2(n_605), .B(n_611), .Y(n_604) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_610), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_610), .A2(n_654), .B(n_655), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_612), .B(n_632), .Y(n_793) );
INVx2_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g630 ( .A(n_614), .Y(n_630) );
NAND2x1p5_ASAP7_75t_L g614 ( .A(n_615), .B(n_623), .Y(n_614) );
NAND2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
AOI21x1_ASAP7_75t_L g623 ( .A1(n_616), .A2(n_624), .B(n_627), .Y(n_623) );
O2A1O1Ixp5_ASAP7_75t_L g637 ( .A1(n_616), .A2(n_638), .B(n_641), .C(n_644), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g892 ( .A1(n_628), .A2(n_869), .B1(n_893), .B2(n_894), .Y(n_892) );
AND2x4_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g684 ( .A(n_630), .B(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_631), .Y(n_893) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_633), .A2(n_733), .B1(n_738), .B2(n_739), .Y(n_732) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_635), .B(n_646), .Y(n_634) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_635), .B(n_712), .Y(n_711) );
INVx2_ASAP7_75t_L g754 ( .A(n_635), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_635), .B(n_835), .Y(n_834) );
AND2x2_ASAP7_75t_L g860 ( .A(n_635), .B(n_699), .Y(n_860) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx2_ASAP7_75t_SL g671 ( .A(n_636), .Y(n_671) );
AND2x2_ASAP7_75t_L g695 ( .A(n_636), .B(n_674), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_636), .B(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g736 ( .A(n_636), .Y(n_736) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g737 ( .A(n_646), .Y(n_737) );
AND2x2_ASAP7_75t_L g780 ( .A(n_646), .B(n_722), .Y(n_780) );
AND2x4_ASAP7_75t_L g790 ( .A(n_646), .B(n_695), .Y(n_790) );
AND2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_660), .Y(n_646) );
INVx2_ASAP7_75t_L g710 ( .A(n_647), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_647), .B(n_736), .Y(n_747) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g699 ( .A(n_648), .B(n_674), .Y(n_699) );
OR2x2_ASAP7_75t_L g712 ( .A(n_648), .B(n_660), .Y(n_712) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_648), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_648), .B(n_674), .Y(n_784) );
AND2x2_ASAP7_75t_L g828 ( .A(n_648), .B(n_673), .Y(n_828) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .B(n_659), .Y(n_652) );
OR2x2_ASAP7_75t_L g672 ( .A(n_660), .B(n_673), .Y(n_672) );
BUFx3_ASAP7_75t_L g693 ( .A(n_660), .Y(n_693) );
INVx2_ASAP7_75t_SL g698 ( .A(n_660), .Y(n_698) );
AND2x2_ASAP7_75t_L g767 ( .A(n_660), .B(n_710), .Y(n_767) );
AND2x2_ASAP7_75t_L g785 ( .A(n_660), .B(n_736), .Y(n_785) );
AND2x2_ASAP7_75t_L g829 ( .A(n_660), .B(n_735), .Y(n_829) );
AO31x2_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .A3(n_664), .B(n_665), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_668), .B(n_684), .Y(n_683) );
INVx5_ASAP7_75t_L g724 ( .A(n_668), .Y(n_724) );
AND2x2_ASAP7_75t_L g755 ( .A(n_668), .B(n_693), .Y(n_755) );
AND2x2_ASAP7_75t_L g797 ( .A(n_668), .B(n_798), .Y(n_797) );
AND2x4_ASAP7_75t_L g859 ( .A(n_668), .B(n_762), .Y(n_859) );
AND2x4_ASAP7_75t_SL g866 ( .A(n_668), .B(n_867), .Y(n_866) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_L g704 ( .A(n_669), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_670), .B(n_851), .Y(n_850) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
NOR2x1_ASAP7_75t_SL g842 ( .A(n_671), .B(n_672), .Y(n_842) );
AND2x2_ASAP7_75t_L g884 ( .A(n_671), .B(n_699), .Y(n_884) );
OR2x2_ASAP7_75t_L g822 ( .A(n_672), .B(n_747), .Y(n_822) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g708 ( .A(n_674), .Y(n_708) );
INVx1_ASAP7_75t_L g746 ( .A(n_674), .Y(n_746) );
OAI33xp33_ASAP7_75t_L g741 ( .A1(n_684), .A2(n_694), .A3(n_742), .B1(n_744), .B2(n_748), .B3(n_749), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_684), .B(n_724), .Y(n_748) );
INVx1_ASAP7_75t_L g846 ( .A(n_684), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g881 ( .A1(n_684), .A2(n_882), .B(n_885), .Y(n_881) );
OR2x2_ASAP7_75t_L g770 ( .A(n_685), .B(n_729), .Y(n_770) );
INVx1_ASAP7_75t_L g810 ( .A(n_685), .Y(n_810) );
OAI221xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_691), .B1(n_696), .B2(n_700), .C(n_702), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_688), .A2(n_854), .B1(n_857), .B2(n_860), .Y(n_853) );
AND2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_690), .Y(n_688) );
NAND2x1_ASAP7_75t_L g852 ( .A(n_689), .B(n_787), .Y(n_852) );
OAI321xp33_ASAP7_75t_L g885 ( .A1(n_689), .A2(n_787), .A3(n_886), .B1(n_888), .B2(n_889), .C(n_892), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_690), .B(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g845 ( .A(n_690), .Y(n_845) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g749 ( .A(n_692), .Y(n_749) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_693), .B(n_699), .Y(n_758) );
A2O1A1Ixp33_ASAP7_75t_L g795 ( .A1(n_693), .A2(n_796), .B(n_799), .C(n_802), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_693), .B(n_787), .C(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_693), .Y(n_812) );
INVx2_ASAP7_75t_L g835 ( .A(n_693), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_694), .A2(n_862), .B1(n_868), .B2(n_870), .C(n_873), .Y(n_861) );
INVx2_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g730 ( .A(n_695), .B(n_731), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_695), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x4_ASAP7_75t_SL g697 ( .A(n_698), .B(n_699), .Y(n_697) );
AND2x2_ASAP7_75t_L g709 ( .A(n_698), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_698), .B(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g764 ( .A(n_699), .Y(n_764) );
NOR2xp33_ASAP7_75t_SL g871 ( .A(n_700), .B(n_725), .Y(n_871) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_701), .B(n_705), .Y(n_738) );
AND2x2_ASAP7_75t_L g769 ( .A(n_701), .B(n_716), .Y(n_769) );
AOI32xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_706), .A3(n_709), .B1(n_711), .B2(n_713), .Y(n_702) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_703), .Y(n_779) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_705), .A2(n_839), .B(n_840), .C(n_843), .Y(n_838) );
INVx1_ASAP7_75t_L g844 ( .A(n_705), .Y(n_844) );
BUFx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g722 ( .A(n_707), .Y(n_722) );
OR2x2_ASAP7_75t_L g816 ( .A(n_707), .B(n_712), .Y(n_816) );
AND2x2_ASAP7_75t_L g880 ( .A(n_709), .B(n_722), .Y(n_880) );
INVx1_ASAP7_75t_L g731 ( .A(n_710), .Y(n_731) );
INVx1_ASAP7_75t_L g856 ( .A(n_712), .Y(n_856) );
INVx2_ASAP7_75t_L g867 ( .A(n_712), .Y(n_867) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g776 ( .A(n_714), .Y(n_776) );
HB1xp67_ASAP7_75t_L g805 ( .A(n_714), .Y(n_805) );
INVx4_ASAP7_75t_L g788 ( .A(n_716), .Y(n_788) );
NOR3xp33_ASAP7_75t_L g717 ( .A(n_718), .B(n_732), .C(n_741), .Y(n_717) );
OAI21xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_723), .B(n_726), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_721), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g851 ( .A(n_722), .B(n_731), .Y(n_851) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
AND2x2_ASAP7_75t_L g727 ( .A(n_724), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g761 ( .A(n_724), .B(n_762), .Y(n_761) );
NAND2x1_ASAP7_75t_L g786 ( .A(n_724), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g819 ( .A(n_724), .B(n_820), .Y(n_819) );
AND2x4_ASAP7_75t_L g877 ( .A(n_724), .B(n_878), .Y(n_877) );
OAI322xp33_ASAP7_75t_L g751 ( .A1(n_725), .A2(n_752), .A3(n_756), .B1(n_758), .B2(n_759), .C1(n_760), .C2(n_763), .Y(n_751) );
INVx1_ASAP7_75t_L g820 ( .A(n_725), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
INVx1_ASAP7_75t_L g759 ( .A(n_727), .Y(n_759) );
INVx1_ASAP7_75t_L g876 ( .A(n_728), .Y(n_876) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g771 ( .A(n_730), .Y(n_771) );
OR2x2_ASAP7_75t_L g833 ( .A(n_731), .B(n_834), .Y(n_833) );
OR2x2_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
NAND2x1_ASAP7_75t_L g888 ( .A(n_734), .B(n_828), .Y(n_888) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AND2x4_ASAP7_75t_L g801 ( .A(n_740), .B(n_792), .Y(n_801) );
AND2x2_ASAP7_75t_L g809 ( .A(n_740), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g832 ( .A(n_740), .Y(n_832) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
OR2x2_ASAP7_75t_L g891 ( .A(n_743), .B(n_793), .Y(n_891) );
INVx1_ASAP7_75t_L g839 ( .A(n_744), .Y(n_839) );
OR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_747), .Y(n_744) );
INVx2_ASAP7_75t_L g757 ( .A(n_746), .Y(n_757) );
INVx2_ASAP7_75t_L g814 ( .A(n_747), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_749), .B(n_884), .Y(n_883) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_765), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_754), .B(n_767), .Y(n_766) );
INVx2_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g806 ( .A(n_757), .Y(n_806) );
AND2x4_ASAP7_75t_L g813 ( .A(n_757), .B(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AND2x2_ASAP7_75t_L g887 ( .A(n_764), .B(n_785), .Y(n_887) );
OAI22xp33_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_770), .B2(n_771), .Y(n_765) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g798 ( .A(n_770), .Y(n_798) );
O2A1O1Ixp33_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_779), .B(n_780), .C(n_781), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_777), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
BUFx2_ASAP7_75t_L g800 ( .A(n_778), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_786), .B1(n_789), .B2(n_791), .Y(n_781) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_782), .A2(n_831), .B1(n_833), .B2(n_836), .Y(n_830) );
INVx4_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_784), .B(n_785), .Y(n_783) );
AND2x4_ASAP7_75t_L g869 ( .A(n_785), .B(n_828), .Y(n_869) );
INVx6_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_788), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
OR2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
AOI211x1_ASAP7_75t_L g794 ( .A1(n_795), .A2(n_806), .B(n_807), .C(n_817), .Y(n_794) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NAND2x1_ASAP7_75t_SL g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g815 ( .A(n_801), .Y(n_815) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_811), .B1(n_815), .B2(n_816), .Y(n_807) );
INVx2_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
OR2x2_ASAP7_75t_L g831 ( .A(n_810), .B(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g865 ( .A(n_810), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_838), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_819), .A2(n_821), .B1(n_823), .B2(n_827), .C(n_830), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g827 ( .A(n_828), .B(n_829), .Y(n_827) );
NAND2xp5_ASAP7_75t_SL g857 ( .A(n_836), .B(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NAND3xp33_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .C(n_846), .Y(n_843) );
NOR2xp67_ASAP7_75t_L g847 ( .A(n_848), .B(n_861), .Y(n_847) );
OAI21xp33_ASAP7_75t_SL g848 ( .A1(n_849), .A2(n_852), .B(n_853), .Y(n_848) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g872 ( .A(n_858), .Y(n_872) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g863 ( .A(n_864), .B(n_866), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx4_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
NOR2x1_ASAP7_75t_L g870 ( .A(n_871), .B(n_872), .Y(n_870) );
OAI21xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_877), .B(n_880), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx1_ASAP7_75t_SL g894 ( .A(n_888), .Y(n_894) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g895 ( .A(n_896), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g898 ( .A1(n_899), .A2(n_901), .B(n_916), .Y(n_898) );
BUFx6f_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
OAI21xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_910), .B(n_913), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_905), .Y(n_904) );
NOR2xp67_ASAP7_75t_SL g914 ( .A(n_905), .B(n_915), .Y(n_914) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx2_ASAP7_75t_SL g906 ( .A(n_907), .Y(n_906) );
NOR2x1p5_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
NOR2xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_918), .Y(n_916) );
BUFx6f_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
CKINVDCx5p33_ASAP7_75t_R g920 ( .A(n_921), .Y(n_920) );
endmodule