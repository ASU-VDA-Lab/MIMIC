module fake_jpeg_19549_n_119 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_119);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_119;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

BUFx16f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_15),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_21),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_59),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_49),
.Y(n_74)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_53),
.B1(n_50),
.B2(n_51),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_73),
.B1(n_1),
.B2(n_3),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_70),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_53),
.B1(n_44),
.B2(n_48),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_88)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_0),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_40),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g87 ( 
.A(n_75),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_42),
.C(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_81),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_63),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_24),
.B1(n_36),
.B2(n_35),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_85),
.B1(n_5),
.B2(n_6),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_1),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_86),
.B(n_4),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_13),
.B1(n_16),
.B2(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_92),
.Y(n_100)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_104),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_91),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_97),
.B(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_97),
.C(n_78),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_109),
.B1(n_103),
.B2(n_89),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_87),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_110),
.B(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_113),
.A2(n_103),
.B1(n_93),
.B2(n_25),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_39),
.B1(n_23),
.B2(n_26),
.Y(n_115)
);

AOI21x1_ASAP7_75t_L g116 ( 
.A1(n_115),
.A2(n_19),
.B(n_27),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_29),
.B(n_30),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_117),
.A2(n_31),
.B(n_33),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_34),
.Y(n_119)
);


endmodule