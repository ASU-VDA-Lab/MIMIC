module fake_jpeg_25598_n_310 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_310);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_310;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_43),
.Y(n_55)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_28),
.B1(n_22),
.B2(n_17),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_34),
.B1(n_16),
.B2(n_33),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_30),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_62),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_57),
.B1(n_22),
.B2(n_17),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_88),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_39),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_72),
.C(n_90),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_22),
.B1(n_17),
.B2(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_66),
.B(n_75),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_46),
.A2(n_26),
.A3(n_41),
.B1(n_37),
.B2(n_39),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_76),
.B(n_92),
.C(n_62),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_39),
.Y(n_72)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_73),
.Y(n_103)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_79),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_50),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_32),
.B1(n_43),
.B2(n_40),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_93),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g94 ( 
.A(n_83),
.B(n_27),
.C(n_31),
.Y(n_94)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_84),
.B(n_23),
.Y(n_97)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g117 ( 
.A(n_85),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_44),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_86),
.A2(n_25),
.B1(n_23),
.B2(n_19),
.Y(n_111)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_34),
.C(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_37),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_122),
.B1(n_115),
.B2(n_93),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_123),
.B(n_105),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_97),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_81),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_99),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_92),
.A2(n_16),
.B1(n_40),
.B2(n_43),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_101),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_27),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_104),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_64),
.B(n_29),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_61),
.B1(n_74),
.B2(n_68),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_88),
.B1(n_72),
.B2(n_82),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_20),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_115),
.B(n_122),
.Y(n_130)
);

O2A1O1Ixp33_ASAP7_75t_L g119 ( 
.A1(n_66),
.A2(n_31),
.B(n_18),
.C(n_21),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_85),
.B1(n_80),
.B2(n_69),
.Y(n_132)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g123 ( 
.A(n_77),
.B(n_18),
.CI(n_23),
.CON(n_123),
.SN(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_125),
.Y(n_179)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_128),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_96),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_127),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_118),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_134),
.B1(n_138),
.B2(n_106),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_139),
.B(n_140),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_90),
.C(n_77),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_110),
.C(n_109),
.Y(n_170)
);

AO21x2_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_73),
.B(n_87),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_104),
.B1(n_109),
.B2(n_110),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_139),
.B1(n_149),
.B2(n_124),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_68),
.B1(n_91),
.B2(n_71),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_123),
.A2(n_71),
.B1(n_19),
.B2(n_25),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_95),
.A2(n_73),
.B1(n_11),
.B2(n_15),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_148),
.B1(n_120),
.B2(n_116),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_13),
.B(n_11),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_89),
.Y(n_144)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_144),
.Y(n_153)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_108),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_150),
.B(n_121),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_151),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_155),
.B1(n_137),
.B2(n_147),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_156),
.B(n_172),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_132),
.A2(n_123),
.B1(n_119),
.B2(n_108),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_169),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_119),
.B1(n_117),
.B2(n_98),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_101),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_162),
.B(n_165),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_117),
.B1(n_98),
.B2(n_100),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_94),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_164),
.A2(n_171),
.B1(n_175),
.B2(n_125),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_136),
.A2(n_100),
.B(n_103),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_145),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_167),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_168),
.B(n_180),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_99),
.B1(n_103),
.B2(n_120),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_180),
.C(n_1),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_0),
.B(n_1),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_173),
.A2(n_178),
.B(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_174),
.B(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_143),
.A2(n_21),
.B1(n_20),
.B2(n_25),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_127),
.B(n_21),
.C(n_20),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_134),
.A2(n_138),
.B1(n_126),
.B2(n_128),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_181),
.A2(n_133),
.B1(n_135),
.B2(n_144),
.Y(n_190)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_183),
.A2(n_191),
.B(n_194),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_196),
.B1(n_197),
.B2(n_173),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_167),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_179),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_190),
.A2(n_193),
.B1(n_195),
.B2(n_205),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_147),
.B(n_145),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_192),
.B(n_198),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_129),
.B1(n_19),
.B2(n_3),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_129),
.B1(n_14),
.B2(n_13),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_13),
.B1(n_12),
.B2(n_10),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_12),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_200),
.B(n_206),
.Y(n_212)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_204),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_162),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_165),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_10),
.C(n_3),
.Y(n_206)
);

AO22x2_ASAP7_75t_L g207 ( 
.A1(n_171),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_207),
.A2(n_153),
.B1(n_177),
.B2(n_174),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g208 ( 
.A(n_160),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_163),
.B(n_9),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_168),
.B(n_2),
.C(n_4),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_178),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_161),
.Y(n_211)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_213),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_187),
.A2(n_207),
.B1(n_211),
.B2(n_204),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_216),
.B1(n_227),
.B2(n_207),
.Y(n_244)
);

OAI22x1_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_162),
.B1(n_158),
.B2(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_222),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_203),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_221),
.B(n_202),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_228),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_153),
.B1(n_162),
.B2(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_231),
.Y(n_234)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_248),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_184),
.B1(n_190),
.B2(n_189),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_239),
.A2(n_245),
.B1(n_247),
.B2(n_219),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_200),
.C(n_206),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_159),
.C(n_188),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_212),
.B(n_226),
.C(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_243),
.B(n_214),
.Y(n_258)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_217),
.A2(n_195),
.B1(n_207),
.B2(n_205),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_246),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_222),
.A2(n_219),
.B1(n_233),
.B2(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_252),
.Y(n_259)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_247),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_264),
.Y(n_279)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_258),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_235),
.B1(n_245),
.B2(n_239),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_260),
.A2(n_263),
.B1(n_268),
.B2(n_152),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_230),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_262),
.B(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_224),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_183),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_265),
.B(n_266),
.Y(n_271)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_212),
.C(n_221),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_240),
.C(n_210),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_235),
.A2(n_208),
.B1(n_162),
.B2(n_203),
.Y(n_268)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_241),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_278),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_238),
.C(n_234),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_159),
.C(n_201),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_260),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_265),
.B(n_199),
.C(n_246),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_259),
.B1(n_261),
.B2(n_264),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_262),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_274),
.B(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_272),
.A2(n_256),
.B1(n_261),
.B2(n_266),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_285),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_271),
.A2(n_258),
.B(n_268),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_277),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_286),
.B(n_282),
.Y(n_297)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_275),
.B(n_273),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_254),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_160),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_287),
.A2(n_199),
.B1(n_166),
.B2(n_152),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_297),
.B(n_281),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_299),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_296),
.A2(n_269),
.B(n_254),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_300),
.B(n_301),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_303),
.A2(n_293),
.B(n_298),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_304),
.C(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_306),
.B(n_291),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_292),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g309 ( 
.A1(n_308),
.A2(n_302),
.A3(n_166),
.B1(n_6),
.B2(n_7),
.C(n_4),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_309),
.A2(n_5),
.B(n_6),
.Y(n_310)
);


endmodule