module real_aes_8521_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_555;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_728;
wire n_598;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_283;
wire n_252;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_1), .A2(n_144), .B(n_148), .C(n_229), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_2), .A2(n_178), .B(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g519 ( .A(n_3), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_4), .B(n_245), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g484 ( .A1(n_5), .A2(n_178), .B(n_485), .Y(n_484) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g219 ( .A(n_7), .Y(n_219) );
INVx1_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g466 ( .A(n_8), .B(n_41), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_9), .A2(n_177), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_10), .B(n_156), .Y(n_231) );
INVx1_ASAP7_75t_L g489 ( .A(n_11), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_12), .B(n_259), .Y(n_543) );
INVx1_ASAP7_75t_L g164 ( .A(n_13), .Y(n_164) );
INVx1_ASAP7_75t_L g555 ( .A(n_14), .Y(n_555) );
A2O1A1Ixp33_ASAP7_75t_L g240 ( .A1(n_15), .A2(n_154), .B(n_241), .C(n_243), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_16), .B(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_17), .B(n_507), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_18), .B(n_178), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_19), .B(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_20), .A2(n_259), .B(n_274), .C(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_21), .B(n_245), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_22), .B(n_156), .Y(n_201) );
A2O1A1Ixp33_ASAP7_75t_L g553 ( .A1(n_23), .A2(n_186), .B(n_243), .C(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_24), .B(n_156), .Y(n_155) );
CKINVDCx16_ASAP7_75t_R g195 ( .A(n_25), .Y(n_195) );
INVx1_ASAP7_75t_L g152 ( .A(n_26), .Y(n_152) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_27), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g227 ( .A(n_28), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_29), .B(n_156), .Y(n_520) );
OAI22xp5_ASAP7_75t_SL g752 ( .A1(n_30), .A2(n_31), .B1(n_753), .B2(n_754), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_30), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_31), .Y(n_753) );
INVx1_ASAP7_75t_L g184 ( .A(n_32), .Y(n_184) );
INVx1_ASAP7_75t_L g498 ( .A(n_33), .Y(n_498) );
INVx2_ASAP7_75t_L g142 ( .A(n_34), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g233 ( .A(n_35), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_36), .A2(n_259), .B(n_260), .C(n_262), .Y(n_258) );
INVxp67_ASAP7_75t_L g185 ( .A(n_37), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_38), .A2(n_148), .B(n_151), .C(n_159), .Y(n_147) );
CKINVDCx14_ASAP7_75t_R g257 ( .A(n_39), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_40), .A2(n_144), .B(n_148), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_41), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g497 ( .A(n_42), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_43), .A2(n_203), .B(n_217), .C(n_218), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_44), .B(n_156), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_45), .A2(n_750), .B1(n_756), .B2(n_757), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_45), .Y(n_756) );
AOI22xp5_ASAP7_75t_L g750 ( .A1(n_46), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_46), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g166 ( .A(n_47), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g180 ( .A(n_48), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_49), .B(n_460), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_50), .A2(n_464), .B1(n_470), .B2(n_758), .Y(n_469) );
INVx1_ASAP7_75t_L g272 ( .A(n_51), .Y(n_272) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_52), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_53), .B(n_178), .Y(n_545) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_54), .A2(n_148), .B1(n_276), .B2(n_496), .Y(n_495) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_55), .A2(n_71), .B1(n_128), .B2(n_129), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_55), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_56), .Y(n_516) );
CKINVDCx14_ASAP7_75t_R g215 ( .A(n_57), .Y(n_215) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_58), .A2(n_217), .B(n_262), .C(n_488), .Y(n_487) );
CKINVDCx20_ASAP7_75t_R g571 ( .A(n_59), .Y(n_571) );
INVx1_ASAP7_75t_L g486 ( .A(n_60), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_61), .A2(n_91), .B1(n_458), .B2(n_459), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_61), .Y(n_459) );
INVx1_ASAP7_75t_L g145 ( .A(n_62), .Y(n_145) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_63), .A2(n_105), .B1(n_119), .B2(n_760), .Y(n_104) );
INVx1_ASAP7_75t_L g163 ( .A(n_64), .Y(n_163) );
INVx1_ASAP7_75t_SL g261 ( .A(n_65), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_66), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_67), .B(n_245), .Y(n_278) );
INVx1_ASAP7_75t_L g198 ( .A(n_68), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_SL g506 ( .A1(n_69), .A2(n_262), .B(n_507), .C(n_508), .Y(n_506) );
INVxp67_ASAP7_75t_L g509 ( .A(n_70), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_71), .Y(n_129) );
INVx1_ASAP7_75t_L g118 ( .A(n_72), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_73), .A2(n_178), .B(n_214), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g207 ( .A(n_74), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_75), .A2(n_178), .B(n_238), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_76), .Y(n_501) );
INVx1_ASAP7_75t_L g565 ( .A(n_77), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_78), .A2(n_177), .B(n_179), .Y(n_176) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_79), .Y(n_146) );
INVx1_ASAP7_75t_L g239 ( .A(n_80), .Y(n_239) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_81), .A2(n_144), .B(n_148), .C(n_567), .Y(n_566) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_82), .A2(n_178), .B(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g242 ( .A(n_83), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_84), .B(n_153), .Y(n_532) );
INVx2_ASAP7_75t_L g161 ( .A(n_85), .Y(n_161) );
INVx1_ASAP7_75t_L g230 ( .A(n_86), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_87), .B(n_507), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_88), .A2(n_144), .B(n_148), .C(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g115 ( .A(n_89), .Y(n_115) );
OR2x2_ASAP7_75t_L g463 ( .A(n_89), .B(n_464), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_L g196 ( .A1(n_90), .A2(n_148), .B(n_197), .C(n_205), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_91), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_92), .B(n_160), .Y(n_490) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_93), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g540 ( .A1(n_94), .A2(n_144), .B(n_148), .C(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_95), .Y(n_547) );
INVx1_ASAP7_75t_L g505 ( .A(n_96), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_97), .Y(n_552) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_98), .B(n_153), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_99), .B(n_168), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_100), .B(n_168), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_101), .B(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g275 ( .A(n_102), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_103), .A2(n_178), .B(n_504), .Y(n_503) );
BUFx4f_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g762 ( .A(n_108), .Y(n_762) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_112), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
NAND3xp33_ASAP7_75t_SL g113 ( .A(n_114), .B(n_115), .C(n_116), .Y(n_113) );
AND2x2_ASAP7_75t_L g465 ( .A(n_114), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g472 ( .A(n_115), .Y(n_472) );
INVx1_ASAP7_75t_L g475 ( .A(n_115), .Y(n_475) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_115), .B(n_464), .Y(n_758) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
AO21x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_124), .B(n_468), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g759 ( .A(n_122), .Y(n_759) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OAI21xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_460), .B(n_467), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_127), .B1(n_130), .B2(n_131), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g534 ( .A(n_128), .B(n_167), .Y(n_534) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
XOR2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_457), .Y(n_131) );
INVx2_ASAP7_75t_L g473 ( .A(n_132), .Y(n_473) );
OR4x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_347), .C(n_394), .D(n_434), .Y(n_132) );
NAND3xp33_ASAP7_75t_SL g133 ( .A(n_134), .B(n_293), .C(n_322), .Y(n_133) );
AOI211xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_208), .B(n_246), .C(n_286), .Y(n_134) );
O2A1O1Ixp33_ASAP7_75t_L g322 ( .A1(n_135), .A2(n_306), .B(n_323), .C(n_327), .Y(n_322) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_137), .B(n_170), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g284 ( .A(n_137), .B(n_285), .Y(n_284) );
INVx3_ASAP7_75t_SL g289 ( .A(n_137), .Y(n_289) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_137), .Y(n_301) );
AND2x4_ASAP7_75t_L g305 ( .A(n_137), .B(n_253), .Y(n_305) );
AND2x2_ASAP7_75t_L g316 ( .A(n_137), .B(n_193), .Y(n_316) );
OR2x2_ASAP7_75t_L g340 ( .A(n_137), .B(n_249), .Y(n_340) );
AND2x2_ASAP7_75t_L g353 ( .A(n_137), .B(n_254), .Y(n_353) );
AND2x2_ASAP7_75t_L g393 ( .A(n_137), .B(n_379), .Y(n_393) );
AND2x2_ASAP7_75t_L g400 ( .A(n_137), .B(n_363), .Y(n_400) );
AND2x2_ASAP7_75t_L g430 ( .A(n_137), .B(n_171), .Y(n_430) );
OR2x6_ASAP7_75t_L g137 ( .A(n_138), .B(n_165), .Y(n_137) );
O2A1O1Ixp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_146), .B(n_147), .C(n_160), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g194 ( .A1(n_139), .A2(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g226 ( .A1(n_139), .A2(n_227), .B(n_228), .Y(n_226) );
OAI22xp33_ASAP7_75t_L g494 ( .A1(n_139), .A2(n_188), .B1(n_495), .B2(n_499), .Y(n_494) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_139), .A2(n_516), .B(n_517), .Y(n_515) );
OAI21xp5_ASAP7_75t_L g564 ( .A1(n_139), .A2(n_565), .B(n_566), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
AND2x4_ASAP7_75t_L g178 ( .A(n_140), .B(n_144), .Y(n_178) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g149 ( .A(n_142), .Y(n_149) );
INVx1_ASAP7_75t_L g277 ( .A(n_142), .Y(n_277) );
INVx1_ASAP7_75t_L g150 ( .A(n_143), .Y(n_150) );
INVx3_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_143), .Y(n_156) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_143), .Y(n_187) );
INVx1_ASAP7_75t_L g507 ( .A(n_143), .Y(n_507) );
BUFx3_ASAP7_75t_L g159 ( .A(n_144), .Y(n_159) );
INVx4_ASAP7_75t_SL g188 ( .A(n_144), .Y(n_188) );
INVx5_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
AND2x6_ASAP7_75t_L g148 ( .A(n_149), .B(n_150), .Y(n_148) );
BUFx3_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_149), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_153), .B(n_155), .C(n_157), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g183 ( .A1(n_153), .A2(n_184), .B1(n_185), .B2(n_186), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_153), .A2(n_519), .B(n_520), .C(n_521), .Y(n_518) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_154), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_154), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_154), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g217 ( .A(n_156), .Y(n_217) );
INVx4_ASAP7_75t_L g259 ( .A(n_156), .Y(n_259) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_158), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g191 ( .A(n_160), .Y(n_191) );
OA21x2_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B(n_220), .Y(n_212) );
INVx1_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_160), .A2(n_550), .B(n_556), .Y(n_549) );
AND2x2_ASAP7_75t_SL g160 ( .A(n_161), .B(n_162), .Y(n_160) );
AND2x2_ASAP7_75t_L g169 ( .A(n_161), .B(n_162), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
AO21x2_ASAP7_75t_L g193 ( .A1(n_167), .A2(n_194), .B(n_206), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_167), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g245 ( .A(n_167), .Y(n_245) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_168), .Y(n_236) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_168), .A2(n_503), .B(n_510), .Y(n_502) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g175 ( .A(n_169), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_170), .B(n_357), .Y(n_369) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_192), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_171), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g307 ( .A(n_171), .B(n_192), .Y(n_307) );
BUFx3_ASAP7_75t_L g315 ( .A(n_171), .Y(n_315) );
OR2x2_ASAP7_75t_L g336 ( .A(n_171), .B(n_211), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_171), .B(n_357), .Y(n_447) );
OA21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_176), .B(n_189), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_173), .A2(n_250), .B(n_251), .Y(n_249) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_173), .A2(n_564), .B(n_570), .Y(n_563) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_SL g528 ( .A1(n_174), .A2(n_529), .B(n_530), .Y(n_528) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_175), .A2(n_494), .B(n_500), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_175), .B(n_501), .Y(n_500) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_175), .A2(n_515), .B(n_522), .Y(n_514) );
INVx1_ASAP7_75t_L g250 ( .A(n_176), .Y(n_250) );
BUFx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_SL g179 ( .A1(n_180), .A2(n_181), .B(n_182), .C(n_188), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_SL g214 ( .A1(n_181), .A2(n_188), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g238 ( .A1(n_181), .A2(n_188), .B(n_239), .C(n_240), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_181), .A2(n_188), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_181), .A2(n_188), .B(n_272), .C(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_181), .A2(n_188), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_181), .A2(n_188), .B(n_505), .C(n_506), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_181), .A2(n_188), .B(n_552), .C(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_186), .B(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_186), .B(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_186), .B(n_555), .Y(n_554) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g200 ( .A(n_187), .Y(n_200) );
OAI22xp5_ASAP7_75t_SL g496 ( .A1(n_187), .A2(n_200), .B1(n_497), .B2(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g205 ( .A(n_188), .Y(n_205) );
INVx1_ASAP7_75t_L g251 ( .A(n_189), .Y(n_251) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_191), .B(n_207), .Y(n_206) );
AO21x2_ASAP7_75t_L g538 ( .A1(n_191), .A2(n_539), .B(n_546), .Y(n_538) );
AND2x2_ASAP7_75t_L g252 ( .A(n_192), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g300 ( .A(n_192), .Y(n_300) );
AND2x2_ASAP7_75t_L g363 ( .A(n_192), .B(n_254), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g365 ( .A1(n_192), .A2(n_366), .B1(n_368), .B2(n_370), .C(n_371), .Y(n_365) );
AND2x2_ASAP7_75t_L g379 ( .A(n_192), .B(n_249), .Y(n_379) );
AND2x2_ASAP7_75t_L g405 ( .A(n_192), .B(n_289), .Y(n_405) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
AND2x2_ASAP7_75t_L g285 ( .A(n_193), .B(n_254), .Y(n_285) );
BUFx2_ASAP7_75t_L g419 ( .A(n_193), .Y(n_419) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_201), .C(n_202), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_L g229 ( .A1(n_199), .A2(n_202), .B(n_230), .C(n_231), .Y(n_229) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_202), .A2(n_532), .B(n_533), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_202), .A2(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g243 ( .A(n_204), .Y(n_243) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
OAI32xp33_ASAP7_75t_L g385 ( .A1(n_209), .A2(n_346), .A3(n_360), .B1(n_386), .B2(n_387), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
AND2x2_ASAP7_75t_L g326 ( .A(n_210), .B(n_268), .Y(n_326) );
INVx1_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
OR2x2_ASAP7_75t_L g308 ( .A(n_211), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_211), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g380 ( .A(n_211), .B(n_268), .Y(n_380) );
AND2x2_ASAP7_75t_L g391 ( .A(n_211), .B(n_283), .Y(n_391) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_L g292 ( .A(n_212), .B(n_269), .Y(n_292) );
AND2x2_ASAP7_75t_L g296 ( .A(n_212), .B(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g331 ( .A(n_212), .B(n_282), .Y(n_331) );
AND2x2_ASAP7_75t_L g338 ( .A(n_212), .B(n_234), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g343 ( .A1(n_212), .A2(n_289), .B(n_300), .C(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g397 ( .A(n_212), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_212), .B(n_223), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_221), .B(n_280), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_221), .B(n_296), .Y(n_386) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
OR2x2_ASAP7_75t_L g291 ( .A(n_222), .B(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_234), .Y(n_222) );
AND2x2_ASAP7_75t_L g283 ( .A(n_223), .B(n_235), .Y(n_283) );
OR2x2_ASAP7_75t_L g298 ( .A(n_223), .B(n_235), .Y(n_298) );
AND2x2_ASAP7_75t_L g321 ( .A(n_223), .B(n_282), .Y(n_321) );
INVx1_ASAP7_75t_L g325 ( .A(n_223), .Y(n_325) );
AND2x2_ASAP7_75t_L g344 ( .A(n_223), .B(n_281), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g354 ( .A1(n_223), .A2(n_309), .B1(n_355), .B2(n_356), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_223), .B(n_397), .Y(n_421) );
AND2x2_ASAP7_75t_L g436 ( .A(n_223), .B(n_296), .Y(n_436) );
INVx4_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
BUFx3_ASAP7_75t_L g266 ( .A(n_224), .Y(n_266) );
AND2x2_ASAP7_75t_L g310 ( .A(n_224), .B(n_235), .Y(n_310) );
AND2x2_ASAP7_75t_L g312 ( .A(n_224), .B(n_268), .Y(n_312) );
AND3x2_ASAP7_75t_L g374 ( .A(n_224), .B(n_338), .C(n_375), .Y(n_374) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_225), .B(n_523), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g546 ( .A(n_225), .B(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_225), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g409 ( .A(n_234), .B(n_281), .Y(n_409) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g268 ( .A(n_235), .B(n_269), .Y(n_268) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_235), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_235), .B(n_280), .Y(n_342) );
NAND3xp33_ASAP7_75t_L g449 ( .A(n_235), .B(n_321), .C(n_397), .Y(n_449) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B(n_244), .Y(n_235) );
OA21x2_ASAP7_75t_L g254 ( .A1(n_236), .A2(n_255), .B(n_264), .Y(n_254) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_236), .A2(n_270), .B(n_278), .Y(n_269) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_245), .A2(n_484), .B(n_490), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_265), .B1(n_279), .B2(n_284), .Y(n_246) );
INVx1_ASAP7_75t_SL g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_252), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_249), .B(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g361 ( .A(n_249), .Y(n_361) );
OAI31xp33_ASAP7_75t_L g377 ( .A1(n_252), .A2(n_378), .A3(n_379), .B(n_380), .Y(n_377) );
AND2x2_ASAP7_75t_L g402 ( .A(n_252), .B(n_289), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_252), .B(n_315), .Y(n_448) );
AND2x2_ASAP7_75t_L g357 ( .A(n_253), .B(n_289), .Y(n_357) );
AND2x2_ASAP7_75t_L g418 ( .A(n_253), .B(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g288 ( .A(n_254), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g346 ( .A(n_254), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_259), .B(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_263), .Y(n_544) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
CKINVDCx16_ASAP7_75t_R g367 ( .A(n_266), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_267), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AOI221x1_ASAP7_75t_SL g334 ( .A1(n_268), .A2(n_335), .B1(n_337), .B2(n_339), .C(n_341), .Y(n_334) );
INVx2_ASAP7_75t_L g282 ( .A(n_269), .Y(n_282) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_269), .Y(n_376) );
INVx2_ASAP7_75t_L g521 ( .A(n_276), .Y(n_521) );
INVx3_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g364 ( .A(n_279), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_280), .B(n_297), .Y(n_389) );
INVx1_ASAP7_75t_SL g452 ( .A(n_280), .Y(n_452) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g370 ( .A(n_283), .B(n_296), .Y(n_370) );
INVx1_ASAP7_75t_L g438 ( .A(n_284), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_284), .B(n_367), .Y(n_451) );
INVx2_ASAP7_75t_SL g290 ( .A(n_285), .Y(n_290) );
AND2x2_ASAP7_75t_L g333 ( .A(n_285), .B(n_289), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_285), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_285), .B(n_360), .Y(n_387) );
AOI21xp33_ASAP7_75t_SL g286 ( .A1(n_287), .A2(n_290), .B(n_291), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_288), .B(n_360), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_288), .B(n_315), .Y(n_456) );
OR2x2_ASAP7_75t_L g328 ( .A(n_289), .B(n_307), .Y(n_328) );
AND2x2_ASAP7_75t_L g427 ( .A(n_289), .B(n_418), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g302 ( .A1(n_290), .A2(n_303), .B1(n_308), .B2(n_311), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_290), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g350 ( .A(n_292), .B(n_298), .Y(n_350) );
INVx1_ASAP7_75t_L g414 ( .A(n_292), .Y(n_414) );
AOI311xp33_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_299), .A3(n_301), .B(n_302), .C(n_313), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_297), .A2(n_429), .B1(n_441), .B2(n_444), .C(n_446), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_297), .B(n_452), .Y(n_454) );
INVx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g351 ( .A(n_299), .Y(n_351) );
AOI211xp5_ASAP7_75t_L g341 ( .A1(n_300), .A2(n_342), .B(n_343), .C(n_345), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_306), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_SL g410 ( .A1(n_304), .A2(n_306), .B(n_411), .C(n_412), .Y(n_410) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_305), .B(n_379), .Y(n_445) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
OAI221xp5_ASAP7_75t_L g327 ( .A1(n_308), .A2(n_328), .B1(n_329), .B2(n_332), .C(n_334), .Y(n_327) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g330 ( .A(n_310), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g413 ( .A(n_310), .B(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_317), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g371 ( .A1(n_314), .A2(n_372), .B(n_373), .C(n_377), .Y(n_371) );
NAND2xp5_ASAP7_75t_SL g314 ( .A(n_315), .B(n_316), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_315), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_315), .B(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g337 ( .A(n_321), .B(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_325), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g439 ( .A(n_328), .Y(n_439) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_331), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g366 ( .A(n_331), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_SL g443 ( .A(n_331), .Y(n_443) );
INVx1_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g384 ( .A(n_333), .B(n_360), .Y(n_384) );
INVx1_ASAP7_75t_SL g378 ( .A(n_340), .Y(n_378) );
INVx1_ASAP7_75t_L g355 ( .A(n_346), .Y(n_355) );
NAND3xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_365), .C(n_381), .Y(n_347) );
AOI322xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .A3(n_352), .B1(n_354), .B2(n_358), .C1(n_362), .C2(n_364), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g401 ( .A1(n_349), .A2(n_402), .B(n_403), .C(n_410), .Y(n_401) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g403 ( .A1(n_352), .A2(n_373), .B1(n_404), .B2(n_406), .Y(n_403) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g362 ( .A(n_360), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g399 ( .A(n_360), .B(n_400), .Y(n_399) );
AOI32xp33_ASAP7_75t_L g450 ( .A1(n_360), .A2(n_451), .A3(n_452), .B1(n_453), .B2(n_455), .Y(n_450) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g372 ( .A(n_363), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g415 ( .A1(n_363), .A2(n_416), .B1(n_420), .B2(n_422), .C(n_425), .Y(n_415) );
AND2x2_ASAP7_75t_L g429 ( .A(n_363), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g432 ( .A(n_367), .B(n_433), .Y(n_432) );
OR2x2_ASAP7_75t_L g442 ( .A(n_367), .B(n_443), .Y(n_442) );
INVxp67_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g433 ( .A(n_376), .B(n_397), .Y(n_433) );
AOI211xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B(n_385), .C(n_388), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI211xp5_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_398), .B(n_401), .C(n_415), .Y(n_394) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_409), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g424 ( .A(n_421), .Y(n_424) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AOI21xp33_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_431), .Y(n_425) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI211xp5_ASAP7_75t_SL g434 ( .A1(n_435), .A2(n_437), .B(n_440), .C(n_450), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_436), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_448), .B(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_467), .A2(n_469), .B(n_759), .Y(n_468) );
XNOR2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_749), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B1(n_474), .B2(n_476), .Y(n_471) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND3x1_ASAP7_75t_L g478 ( .A(n_479), .B(n_671), .C(n_716), .Y(n_478) );
NOR4xp25_ASAP7_75t_L g479 ( .A(n_480), .B(n_594), .C(n_635), .D(n_652), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_511), .B(n_525), .C(n_557), .Y(n_480) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_491), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_482), .B(n_512), .Y(n_511) );
NOR4xp25_ASAP7_75t_L g618 ( .A(n_482), .B(n_612), .C(n_619), .D(n_625), .Y(n_618) );
AND2x2_ASAP7_75t_L g691 ( .A(n_482), .B(n_580), .Y(n_691) );
AND2x2_ASAP7_75t_L g710 ( .A(n_482), .B(n_656), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_482), .B(n_705), .Y(n_719) );
AND2x2_ASAP7_75t_L g732 ( .A(n_482), .B(n_524), .Y(n_732) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g577 ( .A(n_483), .Y(n_577) );
AND2x2_ASAP7_75t_L g584 ( .A(n_483), .B(n_585), .Y(n_584) );
OR2x2_ASAP7_75t_L g634 ( .A(n_483), .B(n_492), .Y(n_634) );
AND2x2_ASAP7_75t_SL g645 ( .A(n_483), .B(n_580), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_483), .B(n_492), .Y(n_649) );
AND2x2_ASAP7_75t_L g658 ( .A(n_483), .B(n_583), .Y(n_658) );
BUFx2_ASAP7_75t_L g681 ( .A(n_483), .Y(n_681) );
AND2x2_ASAP7_75t_L g685 ( .A(n_483), .B(n_502), .Y(n_685) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_502), .Y(n_491) );
AND2x2_ASAP7_75t_L g524 ( .A(n_492), .B(n_502), .Y(n_524) );
BUFx2_ASAP7_75t_L g587 ( .A(n_492), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_492), .A2(n_620), .B1(n_622), .B2(n_623), .Y(n_619) );
OR2x2_ASAP7_75t_L g641 ( .A(n_492), .B(n_514), .Y(n_641) );
AND2x2_ASAP7_75t_L g705 ( .A(n_492), .B(n_583), .Y(n_705) );
INVx3_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g573 ( .A(n_493), .B(n_514), .Y(n_573) );
AND2x2_ASAP7_75t_L g580 ( .A(n_493), .B(n_502), .Y(n_580) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_493), .Y(n_622) );
OR2x2_ASAP7_75t_L g657 ( .A(n_493), .B(n_513), .Y(n_657) );
INVx1_ASAP7_75t_L g576 ( .A(n_502), .Y(n_576) );
INVx3_ASAP7_75t_L g585 ( .A(n_502), .Y(n_585) );
BUFx2_ASAP7_75t_L g609 ( .A(n_502), .Y(n_609) );
AND2x2_ASAP7_75t_L g642 ( .A(n_502), .B(n_577), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_511), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_513), .B(n_585), .Y(n_589) );
INVx1_ASAP7_75t_L g617 ( .A(n_513), .Y(n_617) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g583 ( .A(n_514), .Y(n_583) );
INVx1_ASAP7_75t_L g595 ( .A(n_524), .Y(n_595) );
NAND2x1_ASAP7_75t_SL g525 ( .A(n_526), .B(n_535), .Y(n_525) );
AND2x2_ASAP7_75t_L g593 ( .A(n_526), .B(n_548), .Y(n_593) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_526), .Y(n_667) );
AND2x2_ASAP7_75t_L g694 ( .A(n_526), .B(n_614), .Y(n_694) );
AND2x2_ASAP7_75t_L g702 ( .A(n_526), .B(n_664), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_526), .B(n_560), .Y(n_729) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g561 ( .A(n_527), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g578 ( .A(n_527), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g599 ( .A(n_527), .Y(n_599) );
INVx1_ASAP7_75t_L g605 ( .A(n_527), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_527), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g638 ( .A(n_527), .B(n_563), .Y(n_638) );
OR2x2_ASAP7_75t_L g676 ( .A(n_527), .B(n_631), .Y(n_676) );
AOI32xp33_ASAP7_75t_L g688 ( .A1(n_527), .A2(n_689), .A3(n_692), .B1(n_693), .B2(n_694), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_527), .B(n_664), .Y(n_728) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_527), .B(n_624), .Y(n_739) );
OR2x6_ASAP7_75t_L g527 ( .A(n_528), .B(n_534), .Y(n_527) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g650 ( .A(n_536), .B(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_548), .Y(n_536) );
INVx1_ASAP7_75t_L g612 ( .A(n_537), .Y(n_612) );
AND2x2_ASAP7_75t_L g614 ( .A(n_537), .B(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_537), .B(n_562), .Y(n_631) );
AND2x2_ASAP7_75t_L g664 ( .A(n_537), .B(n_640), .Y(n_664) );
AND2x2_ASAP7_75t_L g701 ( .A(n_537), .B(n_563), .Y(n_701) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g560 ( .A(n_538), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_538), .B(n_562), .Y(n_591) );
AND2x2_ASAP7_75t_L g598 ( .A(n_538), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g639 ( .A(n_538), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_545), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_543), .B(n_544), .Y(n_541) );
INVx2_ASAP7_75t_L g615 ( .A(n_548), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_548), .B(n_562), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_548), .B(n_606), .Y(n_687) );
INVx1_ASAP7_75t_L g709 ( .A(n_548), .Y(n_709) );
INVx1_ASAP7_75t_L g726 ( .A(n_548), .Y(n_726) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g579 ( .A(n_549), .B(n_562), .Y(n_579) );
AND2x2_ASAP7_75t_L g601 ( .A(n_549), .B(n_563), .Y(n_601) );
INVx1_ASAP7_75t_L g640 ( .A(n_549), .Y(n_640) );
AOI221x1_ASAP7_75t_SL g557 ( .A1(n_558), .A2(n_572), .B1(n_578), .B2(n_580), .C(n_581), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_558), .A2(n_645), .B1(n_712), .B2(n_713), .Y(n_711) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
AND2x2_ASAP7_75t_L g603 ( .A(n_559), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g698 ( .A(n_559), .B(n_578), .Y(n_698) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g654 ( .A(n_560), .B(n_579), .Y(n_654) );
INVx1_ASAP7_75t_L g666 ( .A(n_561), .Y(n_666) );
AND2x2_ASAP7_75t_L g677 ( .A(n_561), .B(n_664), .Y(n_677) );
AND2x2_ASAP7_75t_L g744 ( .A(n_561), .B(n_639), .Y(n_744) );
INVx2_ASAP7_75t_L g606 ( .A(n_562), .Y(n_606) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_573), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g696 ( .A(n_573), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_574), .B(n_657), .Y(n_660) );
INVx3_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AOI21xp5_ASAP7_75t_L g740 ( .A1(n_575), .A2(n_696), .B(n_741), .Y(n_740) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR2xp33_ASAP7_75t_SL g718 ( .A(n_578), .B(n_604), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_579), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g670 ( .A(n_579), .B(n_598), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_579), .B(n_605), .Y(n_747) );
AND2x2_ASAP7_75t_L g616 ( .A(n_580), .B(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g683 ( .A(n_580), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_590), .Y(n_581) );
NAND2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_583), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g632 ( .A(n_583), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g644 ( .A(n_583), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_583), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g668 ( .A(n_584), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_584), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_584), .B(n_587), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_587), .A2(n_626), .B(n_656), .C(n_658), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g673 ( .A1(n_587), .A2(n_674), .B1(n_677), .B2(n_678), .C(n_682), .Y(n_673) );
AND2x2_ASAP7_75t_L g669 ( .A(n_588), .B(n_622), .Y(n_669) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g629 ( .A(n_593), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g700 ( .A(n_593), .B(n_701), .Y(n_700) );
OAI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B(n_602), .C(n_627), .Y(n_594) );
NAND3xp33_ASAP7_75t_SL g713 ( .A(n_595), .B(n_714), .C(n_715), .Y(n_713) );
OR2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_600), .Y(n_596) );
OR2x2_ASAP7_75t_L g686 ( .A(n_597), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_607), .B1(n_610), .B2(n_616), .C(n_618), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_604), .B(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_604), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g626 ( .A(n_609), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_609), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_665) );
OR2x2_ASAP7_75t_L g746 ( .A(n_609), .B(n_657), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g610 ( .A(n_611), .B(n_613), .Y(n_610) );
INVxp67_ASAP7_75t_L g720 ( .A(n_612), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_614), .B(n_735), .Y(n_734) );
INVxp67_ASAP7_75t_L g621 ( .A(n_615), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_617), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_617), .B(n_664), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_617), .B(n_684), .Y(n_723) );
HB1xp67_ASAP7_75t_L g647 ( .A(n_621), .Y(n_647) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g737 ( .A(n_626), .B(n_657), .Y(n_737) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_632), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g715 ( .A(n_632), .Y(n_715) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OAI322xp33_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_641), .A3(n_642), .B1(n_643), .B2(n_646), .C1(n_648), .C2(n_650), .Y(n_635) );
OAI322xp33_ASAP7_75t_L g717 ( .A1(n_636), .A2(n_718), .A3(n_719), .B1(n_720), .B2(n_721), .C1(n_722), .C2(n_724), .Y(n_717) );
CKINVDCx16_ASAP7_75t_R g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
INVx4_ASAP7_75t_L g651 ( .A(n_638), .Y(n_651) );
AND2x2_ASAP7_75t_L g712 ( .A(n_638), .B(n_664), .Y(n_712) );
AND2x2_ASAP7_75t_L g725 ( .A(n_638), .B(n_726), .Y(n_725) );
CKINVDCx16_ASAP7_75t_R g736 ( .A(n_641), .Y(n_736) );
INVx1_ASAP7_75t_L g714 ( .A(n_642), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
OR2x2_ASAP7_75t_L g648 ( .A(n_644), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g731 ( .A(n_644), .B(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_644), .B(n_685), .Y(n_742) );
OR2x2_ASAP7_75t_L g675 ( .A(n_647), .B(n_676), .Y(n_675) );
INVxp33_ASAP7_75t_L g692 ( .A(n_647), .Y(n_692) );
OAI221xp5_ASAP7_75t_SL g652 ( .A1(n_651), .A2(n_653), .B1(n_655), .B2(n_659), .C(n_661), .Y(n_652) );
NOR2xp67_ASAP7_75t_L g708 ( .A(n_651), .B(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g735 ( .A(n_651), .Y(n_735) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx3_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g699 ( .A1(n_658), .A2(n_683), .A3(n_700), .B1(n_702), .B2(n_703), .C1(n_706), .C2(n_710), .Y(n_699) );
INVxp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B1(n_669), .B2(n_670), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_695), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_673), .B(n_688), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_676), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g678 ( .A(n_679), .Y(n_678) );
NAND2xp33_ASAP7_75t_SL g693 ( .A(n_679), .B(n_690), .Y(n_693) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
OAI322xp33_ASAP7_75t_L g733 ( .A1(n_681), .A2(n_734), .A3(n_736), .B1(n_737), .B2(n_738), .C1(n_740), .C2(n_743), .Y(n_733) );
AOI21xp33_ASAP7_75t_SL g682 ( .A1(n_683), .A2(n_684), .B(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_691), .B(n_739), .Y(n_748) );
OAI211xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_697), .B(n_699), .C(n_711), .Y(n_695) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NOR4xp25_ASAP7_75t_L g716 ( .A(n_717), .B(n_727), .C(n_733), .D(n_745), .Y(n_716) );
INVxp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
CKINVDCx14_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
OAI21xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_747), .B(n_748), .Y(n_745) );
CKINVDCx16_ASAP7_75t_R g757 ( .A(n_750), .Y(n_757) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
endmodule