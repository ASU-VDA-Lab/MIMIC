module fake_jpeg_21186_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_28),
.B(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_0),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_37),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_23),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_42),
.B(n_50),
.Y(n_61)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_14),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_35),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_28),
.B(n_14),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.C(n_35),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g49 ( 
.A1(n_28),
.A2(n_14),
.B1(n_20),
.B2(n_24),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_35),
.A3(n_34),
.B1(n_37),
.B2(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_13),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_53),
.B(n_63),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_69),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_33),
.B1(n_31),
.B2(n_34),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_56),
.A2(n_73),
.B1(n_41),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_65),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_48),
.A2(n_37),
.B1(n_31),
.B2(n_33),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_15),
.C(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_18),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_23),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_17),
.B1(n_13),
.B2(n_25),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_18),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_17),
.B1(n_37),
.B2(n_26),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_22),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_85),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_51),
.A2(n_66),
.B(n_57),
.C(n_68),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_78),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_84),
.B1(n_56),
.B2(n_52),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_41),
.B1(n_43),
.B2(n_27),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_89),
.B(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_93),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g94 ( 
.A(n_77),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_SL g101 ( 
.A1(n_94),
.A2(n_95),
.A3(n_96),
.B1(n_84),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_74),
.B(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_87),
.B(n_55),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_107),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_79),
.B(n_88),
.C(n_87),
.D(n_85),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_15),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_76),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_91),
.C(n_89),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_83),
.B(n_80),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_81),
.B(n_94),
.C(n_77),
.D(n_67),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_9),
.A3(n_11),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_112),
.C(n_114),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_100),
.A2(n_83),
.B1(n_73),
.B2(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_111),
.Y(n_116)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_52),
.C(n_58),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_113),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_103),
.B(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_117),
.B(n_118),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_102),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_116),
.A2(n_113),
.B1(n_109),
.B2(n_94),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_69),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_15),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_123),
.Y(n_125)
);

OAI21x1_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_116),
.B(n_64),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_120),
.A2(n_16),
.B(n_22),
.Y(n_124)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_126),
.A3(n_16),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_2),
.Y(n_128)
);

OAI21x1_ASAP7_75t_L g127 ( 
.A1(n_125),
.A2(n_122),
.B(n_3),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.C(n_5),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_129),
.Y(n_130)
);


endmodule