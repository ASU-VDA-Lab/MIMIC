module fake_jpeg_8599_n_259 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_37),
.B(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_40),
.A2(n_17),
.B1(n_31),
.B2(n_29),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_41),
.A2(n_56),
.B1(n_16),
.B2(n_21),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_43),
.A2(n_45),
.B1(n_50),
.B2(n_26),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_35),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_36),
.B(n_25),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_53),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_21),
.B1(n_19),
.B2(n_18),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_47),
.A2(n_18),
.B1(n_19),
.B2(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_17),
.B1(n_31),
.B2(n_22),
.Y(n_50)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_36),
.B(n_18),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_37),
.A2(n_24),
.B1(n_31),
.B2(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_36),
.B(n_25),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_57),
.B(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_60),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_59),
.B(n_85),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_57),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_32),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_61),
.A2(n_62),
.B1(n_74),
.B2(n_83),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_52),
.A2(n_26),
.B1(n_25),
.B2(n_19),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g109 ( 
.A(n_63),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_71),
.Y(n_92)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_68),
.B1(n_57),
.B2(n_77),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_75),
.B1(n_84),
.B2(n_43),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_28),
.B1(n_21),
.B2(n_23),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_49),
.A2(n_35),
.B1(n_16),
.B2(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_48),
.B(n_16),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_47),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_65),
.B1(n_73),
.B2(n_84),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_28),
.B1(n_21),
.B2(n_27),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_34),
.B(n_33),
.C(n_36),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_55),
.A2(n_28),
.B1(n_10),
.B2(n_2),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_56),
.B1(n_41),
.B2(n_50),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_87),
.A2(n_90),
.B1(n_110),
.B2(n_70),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_89),
.A2(n_11),
.B1(n_15),
.B2(n_2),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_72),
.A2(n_71),
.B1(n_81),
.B2(n_85),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_101),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_47),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_82),
.B(n_47),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_70),
.B1(n_67),
.B2(n_66),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_47),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_106),
.B(n_107),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_55),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_108),
.B(n_111),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_45),
.B(n_34),
.C(n_33),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g112 ( 
.A1(n_69),
.A2(n_21),
.A3(n_27),
.B1(n_55),
.B2(n_54),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_54),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_107),
.B(n_0),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_113),
.A2(n_134),
.B(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_114),
.B(n_118),
.Y(n_162)
);

BUFx10_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_58),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_63),
.B1(n_79),
.B2(n_27),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_119),
.A2(n_135),
.B1(n_104),
.B2(n_105),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_120),
.A2(n_139),
.B1(n_104),
.B2(n_109),
.Y(n_148)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_122),
.B(n_124),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_9),
.Y(n_124)
);

AO22x1_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_106),
.B1(n_101),
.B2(n_88),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_129),
.Y(n_155)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_8),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_0),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_94),
.B(n_11),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_89),
.A2(n_78),
.B(n_1),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_137),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_8),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_138),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_90),
.C(n_91),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_142),
.C(n_159),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_91),
.C(n_88),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_134),
.A2(n_111),
.B1(n_103),
.B2(n_109),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_144),
.A2(n_148),
.B1(n_150),
.B2(n_166),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_109),
.B1(n_105),
.B2(n_3),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_157),
.B(n_161),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_118),
.A2(n_93),
.B1(n_99),
.B2(n_3),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_137),
.B(n_115),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_121),
.B(n_1),
.Y(n_158)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_93),
.C(n_99),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_128),
.B(n_93),
.C(n_67),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_119),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_1),
.B(n_66),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_113),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_4),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_2),
.Y(n_164)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_153),
.B(n_114),
.Y(n_167)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_126),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_169),
.B(n_174),
.Y(n_194)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_164),
.C(n_151),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_178),
.Y(n_200)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_131),
.B(n_125),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_180),
.B(n_181),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_162),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_145),
.B(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_160),
.C(n_144),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_129),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_125),
.CI(n_122),
.CON(n_179),
.SN(n_179)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_179),
.B(n_182),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_156),
.B(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_120),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_183),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_186),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_165),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_115),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_149),
.B(n_6),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_170),
.A2(n_143),
.B1(n_150),
.B2(n_156),
.Y(n_189)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_189),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_146),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_190),
.B(n_179),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_203),
.C(n_205),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_148),
.B1(n_166),
.B2(n_152),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_192),
.A2(n_195),
.B1(n_202),
.B2(n_181),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_157),
.B1(n_165),
.B2(n_141),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_149),
.B1(n_141),
.B2(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_198),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_174),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_6),
.C(n_12),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_176),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_199),
.A2(n_177),
.B(n_169),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_213),
.B1(n_210),
.B2(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_194),
.B(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_177),
.B(n_173),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_190),
.B(n_178),
.C(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_198),
.Y(n_215)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_215),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_216),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_200),
.B(n_188),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_220),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_184),
.C(n_175),
.Y(n_219)
);

AOI321xp33_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_173),
.A3(n_184),
.B1(n_188),
.B2(n_182),
.C(n_185),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_212),
.A2(n_196),
.B1(n_204),
.B2(n_193),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_211),
.B1(n_209),
.B2(n_202),
.Y(n_236)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_199),
.B(n_193),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_227),
.A2(n_213),
.B(n_211),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_228),
.B(n_214),
.Y(n_238)
);

AO22x1_ASAP7_75t_L g230 ( 
.A1(n_212),
.A2(n_189),
.B1(n_192),
.B2(n_220),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_224),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_233),
.B(n_236),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_239),
.B1(n_227),
.B2(n_229),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_223),
.B(n_197),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_238),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_196),
.C(n_203),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_226),
.B(n_221),
.Y(n_244)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_222),
.B(n_230),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_246),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_239),
.C(n_234),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_235),
.A2(n_231),
.B1(n_186),
.B2(n_206),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_241),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_249),
.B(n_250),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_245),
.B(n_187),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_252),
.Y(n_253)
);

NAND4xp25_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_186),
.C(n_13),
.D(n_14),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_243),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_254),
.B(n_13),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_257),
.B(n_253),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_255),
.B(n_13),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_14),
.Y(n_259)
);


endmodule