module fake_jpeg_16390_n_374 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_374);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_374;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_7),
.Y(n_38)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_39),
.B(n_42),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_6),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_18),
.Y(n_68)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_41),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_46),
.B(n_48),
.Y(n_89)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_54),
.Y(n_110)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_28),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_60),
.B(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_23),
.B(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_65),
.B(n_26),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_41),
.A2(n_14),
.B1(n_33),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_67),
.A2(n_71),
.B1(n_79),
.B2(n_81),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_80),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_32),
.B1(n_19),
.B2(n_22),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_84),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_60),
.A2(n_18),
.B1(n_25),
.B2(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_40),
.B(n_64),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_18),
.B1(n_25),
.B2(n_12),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_39),
.A2(n_34),
.B1(n_23),
.B2(n_30),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_83),
.B(n_85),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_49),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_32),
.C(n_19),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_25),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_87),
.B(n_95),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_30),
.B1(n_28),
.B2(n_26),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_91),
.A2(n_101),
.B1(n_103),
.B2(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_46),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_104),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_17),
.B(n_31),
.C(n_27),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_100),
.B(n_0),
.C(n_1),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_53),
.A2(n_17),
.B(n_31),
.C(n_27),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_22),
.B1(n_32),
.B2(n_19),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_45),
.A2(n_32),
.B1(n_22),
.B2(n_31),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_52),
.B(n_22),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_63),
.A2(n_31),
.B1(n_27),
.B2(n_35),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_59),
.A2(n_27),
.B1(n_31),
.B2(n_9),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_5),
.B(n_12),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_10),
.B(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_51),
.A2(n_27),
.B1(n_8),
.B2(n_13),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_111),
.B1(n_4),
.B2(n_8),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_51),
.A2(n_55),
.B1(n_61),
.B2(n_56),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_52),
.B(n_35),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_0),
.Y(n_146)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_57),
.B1(n_10),
.B2(n_3),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_116),
.A2(n_122),
.B(n_136),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_80),
.B(n_57),
.CI(n_48),
.CON(n_117),
.SN(n_117)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_117),
.B(n_124),
.Y(n_202)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_92),
.A2(n_77),
.B1(n_90),
.B2(n_82),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_96),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_127),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_58),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g128 ( 
.A(n_83),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_128),
.B(n_131),
.Y(n_187)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_98),
.A2(n_61),
.B1(n_44),
.B2(n_35),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_130),
.A2(n_145),
.B1(n_157),
.B2(n_124),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_78),
.B(n_5),
.Y(n_131)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_133),
.Y(n_205)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_90),
.A2(n_5),
.B1(n_11),
.B2(n_3),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_137),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_138),
.B(n_140),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_8),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_104),
.A2(n_44),
.B1(n_35),
.B2(n_8),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_141),
.A2(n_155),
.B1(n_1),
.B2(n_85),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_147),
.B1(n_66),
.B2(n_69),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_94),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_143),
.B(n_159),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_SL g192 ( 
.A1(n_144),
.A2(n_132),
.B(n_146),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_68),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_138),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_66),
.A2(n_11),
.B1(n_1),
.B2(n_2),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_100),
.B(n_105),
.Y(n_178)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_107),
.Y(n_151)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_74),
.Y(n_152)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_81),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_155)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_70),
.A2(n_2),
.B(n_0),
.Y(n_156)
);

OR2x2_ASAP7_75t_SL g207 ( 
.A(n_156),
.B(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_94),
.Y(n_159)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_114),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_163),
.Y(n_197)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_97),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_76),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_164),
.B(n_143),
.Y(n_182)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_113),
.Y(n_165)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_165),
.Y(n_170)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_166),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_167),
.A2(n_168),
.B1(n_180),
.B2(n_181),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_174),
.B(n_183),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_132),
.B(n_112),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_185),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_178),
.A2(n_184),
.B(n_186),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_158),
.A2(n_82),
.B1(n_69),
.B2(n_86),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_115),
.B1(n_93),
.B2(n_71),
.Y(n_181)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

A2O1A1Ixp33_ASAP7_75t_SL g184 ( 
.A1(n_142),
.A2(n_111),
.B(n_93),
.C(n_88),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_118),
.B(n_76),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_93),
.B(n_72),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_72),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_195),
.B(n_164),
.C(n_153),
.D(n_166),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_128),
.A2(n_150),
.B1(n_117),
.B2(n_149),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_190),
.A2(n_198),
.B1(n_204),
.B2(n_206),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_192),
.A2(n_174),
.B1(n_207),
.B2(n_185),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_118),
.B(n_117),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_178),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_123),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_166),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_118),
.A2(n_139),
.B(n_162),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_160),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_126),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_148),
.A2(n_150),
.B1(n_141),
.B2(n_133),
.Y(n_198)
);

NOR2x1_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_151),
.Y(n_200)
);

NAND2x1p5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_120),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_121),
.A2(n_154),
.B1(n_129),
.B2(n_134),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_120),
.A2(n_119),
.B1(n_152),
.B2(n_161),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_165),
.C(n_166),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_171),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_213),
.B(n_222),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_214),
.B(n_250),
.Y(n_270)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_216),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_217),
.A2(n_227),
.B(n_245),
.Y(n_264)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_173),
.Y(n_218)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_218),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_221),
.Y(n_260)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_189),
.B(n_191),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_225),
.B(n_237),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_228),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_231),
.B(n_234),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_137),
.C(n_135),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_246),
.C(n_168),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_238),
.Y(n_269)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_170),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_236),
.A2(n_244),
.B1(n_247),
.B2(n_249),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_126),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_194),
.B(n_200),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_239),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_135),
.B1(n_137),
.B2(n_198),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_180),
.B1(n_184),
.B2(n_181),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_135),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_241),
.B(n_242),
.Y(n_281)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_212),
.A2(n_193),
.B1(n_202),
.B2(n_174),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_243),
.A2(n_242),
.B1(n_228),
.B2(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_176),
.B(n_188),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_201),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_182),
.B(n_187),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_227),
.B(n_215),
.Y(n_275)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_251),
.A2(n_211),
.B1(n_203),
.B2(n_179),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_186),
.B(n_184),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_SL g297 ( 
.A(n_253),
.B(n_267),
.C(n_279),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_197),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_254),
.B(n_257),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_261),
.A2(n_282),
.B1(n_283),
.B2(n_253),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_184),
.B1(n_208),
.B2(n_170),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_263),
.A2(n_266),
.B1(n_276),
.B2(n_278),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_229),
.A2(n_249),
.B1(n_252),
.B2(n_214),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_232),
.B(n_208),
.C(n_175),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_271),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_175),
.C(n_201),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_219),
.A2(n_184),
.B1(n_211),
.B2(n_210),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_251),
.B1(n_238),
.B2(n_236),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_205),
.C(n_196),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_275),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_245),
.B1(n_240),
.B2(n_243),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_223),
.A2(n_233),
.B1(n_215),
.B2(n_237),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_233),
.A2(n_210),
.B1(n_231),
.B2(n_218),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_221),
.B(n_224),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_282),
.B1(n_284),
.B2(n_260),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_216),
.B1(n_244),
.B2(n_226),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_288),
.A2(n_290),
.B1(n_304),
.B2(n_305),
.Y(n_317)
);

BUFx12_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_255),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_292),
.B(n_294),
.Y(n_328)
);

INVx13_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_293),
.A2(n_303),
.B1(n_306),
.B2(n_308),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_262),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_269),
.B(n_278),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_295),
.B(n_302),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_274),
.C(n_264),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_277),
.B(n_260),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_298),
.B(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_280),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_285),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_269),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_259),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_254),
.C(n_257),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_297),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_266),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_258),
.B1(n_284),
.B2(n_282),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_261),
.A2(n_263),
.B1(n_271),
.B2(n_276),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_310),
.A2(n_308),
.B1(n_290),
.B2(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_280),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_264),
.B(n_272),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_313),
.A2(n_320),
.B1(n_321),
.B2(n_323),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_270),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_315),
.B(n_323),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_326),
.C(n_289),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_318),
.A2(n_320),
.B1(n_322),
.B2(n_332),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_319),
.B(n_314),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_307),
.C(n_301),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_321),
.B(n_331),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_310),
.A2(n_295),
.B1(n_292),
.B2(n_301),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_299),
.B(n_291),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_291),
.B(n_296),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_329),
.B(n_315),
.Y(n_345)
);

NOR3xp33_ASAP7_75t_SL g331 ( 
.A(n_297),
.B(n_293),
.C(n_289),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_309),
.A2(n_303),
.B1(n_308),
.B2(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_334),
.B(n_336),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_335),
.B(n_344),
.C(n_343),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_317),
.A2(n_329),
.B1(n_324),
.B2(n_322),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_325),
.B(n_324),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_337),
.B(n_333),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_331),
.B(n_314),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_338),
.A2(n_346),
.B1(n_348),
.B2(n_347),
.Y(n_358)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_330),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_330),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_342),
.B(n_347),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_326),
.B(n_316),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_340),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_328),
.A2(n_318),
.B(n_319),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_350),
.C(n_355),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_344),
.C(n_343),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_351),
.B(n_352),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g352 ( 
.A1(n_346),
.A2(n_339),
.B(n_336),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_358),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_338),
.B(n_340),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_356),
.B(n_341),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_359),
.B(n_360),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_342),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_334),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_364),
.B(n_357),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_365),
.B(n_362),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_361),
.B(n_355),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_367),
.B(n_361),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_368),
.A2(n_369),
.B(n_366),
.C(n_367),
.Y(n_370)
);

AOI21x1_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_363),
.B(n_349),
.Y(n_371)
);

BUFx24_ASAP7_75t_SL g372 ( 
.A(n_371),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_350),
.C(n_363),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_373),
.B(n_353),
.Y(n_374)
);


endmodule