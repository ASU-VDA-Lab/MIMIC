module fake_aes_5813_n_33 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x6_ASAP7_75t_L g13 ( .A(n_1), .B(n_11), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_12), .Y(n_14) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_8), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_10), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_16), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_20), .A2(n_13), .B1(n_16), .B2(n_14), .Y(n_22) );
AOI22xp5_ASAP7_75t_L g23 ( .A1(n_20), .A2(n_15), .B1(n_13), .B2(n_2), .Y(n_23) );
OR2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_25), .B(n_19), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_25), .B(n_22), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_19), .B1(n_1), .B2(n_2), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_0), .A3(n_3), .B1(n_4), .B2(n_5), .C1(n_13), .C2(n_9), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
XNOR2xp5_ASAP7_75t_L g31 ( .A(n_29), .B(n_0), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
AOI322xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_31), .A3(n_4), .B1(n_5), .B2(n_3), .C1(n_13), .C2(n_7), .Y(n_33) );
endmodule