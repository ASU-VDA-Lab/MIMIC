module fake_jpeg_2886_n_157 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_25),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_43),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_52),
.Y(n_56)
);

CKINVDCx9p33_ASAP7_75t_R g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_45),
.C(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_2),
.Y(n_64)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_39),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_70),
.Y(n_82)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_51),
.B1(n_44),
.B2(n_47),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_53),
.B1(n_18),
.B2(n_19),
.Y(n_92)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_54),
.B(n_55),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_81),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_69),
.B(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_79),
.Y(n_96)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_66),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_80),
.B(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_39),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_66),
.A2(n_39),
.B1(n_44),
.B2(n_52),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_53),
.B(n_5),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_85),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_3),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_93),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_101),
.Y(n_110)
);

OR2x4_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_72),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_98),
.B(n_9),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_3),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_4),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_8),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_76),
.B(n_53),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_6),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_107),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_22),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_7),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_8),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_109),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_113),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_14),
.B(n_15),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_97),
.B(n_10),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_117),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_26),
.C(n_13),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_115),
.B(n_24),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_100),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_121),
.A2(n_103),
.B(n_29),
.Y(n_141)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_107),
.Y(n_124)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_16),
.CI(n_17),
.CON(n_127),
.SN(n_127)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_127),
.B(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_116),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_102),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_132),
.C(n_130),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_38),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_132),
.C(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_119),
.B1(n_137),
.B2(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_143),
.B(n_137),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_131),
.C(n_135),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_147),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_151),
.B(n_123),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_150),
.B(n_146),
.C(n_145),
.D(n_126),
.Y(n_153)
);

NOR2xp67_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_127),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_154),
.B(n_28),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_SL g156 ( 
.A1(n_155),
.A2(n_30),
.B(n_31),
.C(n_35),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_37),
.Y(n_157)
);


endmodule