module fake_jpeg_28522_n_148 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_148);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_148;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_12),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_1),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_1),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_2),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_44),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_57),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_57),
.B1(n_43),
.B2(n_48),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_50),
.B1(n_45),
.B2(n_47),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_49),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_58),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_88),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_45),
.B1(n_59),
.B2(n_50),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_86),
.A2(n_70),
.B1(n_4),
.B2(n_5),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_82),
.A2(n_47),
.B1(n_55),
.B2(n_54),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_94),
.B(n_96),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_52),
.B(n_53),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_95),
.B(n_97),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_81),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_80),
.B(n_2),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_99),
.B(n_100),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_18),
.B(n_40),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_118),
.B1(n_42),
.B2(n_33),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_107),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_5),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_24),
.B1(n_38),
.B2(n_37),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_6),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_17),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_112),
.B(n_85),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_7),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_7),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_8),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_122),
.B(n_125),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_108),
.A2(n_9),
.B(n_10),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_123),
.A2(n_128),
.B(n_131),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_102),
.A2(n_9),
.B(n_11),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_124),
.A2(n_103),
.B(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_19),
.B(n_29),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_112),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_110),
.B1(n_104),
.B2(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_122),
.B1(n_130),
.B2(n_135),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_136),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_142),
.A2(n_141),
.B(n_140),
.Y(n_143)
);

OAI31xp33_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_139),
.A3(n_120),
.B(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_129),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_124),
.B(n_138),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_137),
.C(n_101),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_32),
.B(n_34),
.Y(n_148)
);


endmodule