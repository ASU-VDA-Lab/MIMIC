module fake_netlist_1_1137_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
OR2x6_ASAP7_75t_L g3 ( .A(n_2), .B(n_0), .Y(n_3) );
INVx2_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
AOI21xp5_ASAP7_75t_L g5 ( .A1(n_3), .A2(n_0), .B(n_1), .Y(n_5) );
NOR2xp33_ASAP7_75t_SL g6 ( .A(n_3), .B(n_0), .Y(n_6) );
NOR2xp33_ASAP7_75t_L g7 ( .A(n_6), .B(n_3), .Y(n_7) );
INVxp33_ASAP7_75t_SL g8 ( .A(n_6), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_5), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_4), .Y(n_10) );
AOI321xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_8), .C(n_9), .Y(n_11) );
OAI211xp5_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_1), .B(n_2), .C(n_0), .Y(n_12) );
AOI211xp5_ASAP7_75t_L g13 ( .A1(n_12), .A2(n_0), .B(n_2), .C(n_1), .Y(n_13) );
NAND4xp75_ASAP7_75t_L g14 ( .A(n_11), .B(n_1), .C(n_2), .D(n_7), .Y(n_14) );
AOI22x1_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_11), .B1(n_1), .B2(n_2), .Y(n_15) );
NAND2xp33_ASAP7_75t_L g16 ( .A(n_15), .B(n_13), .Y(n_16) );
endmodule