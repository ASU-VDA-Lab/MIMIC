module fake_ariane_3349_n_1738 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1738);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1738;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1614;
wire n_1162;
wire n_536;
wire n_1377;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

BUFx3_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_93),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_47),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_87),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_70),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_50),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_62),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_34),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_19),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_152),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_2),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_3),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_24),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_17),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_54),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_94),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_26),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_48),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_30),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_18),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_117),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_40),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_72),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_98),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_55),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_0),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_21),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_150),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_33),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_4),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_146),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_115),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_38),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_18),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_7),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_105),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_131),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_55),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_107),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_90),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_85),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_45),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_83),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_114),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_49),
.Y(n_225)
);

CKINVDCx11_ASAP7_75t_R g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_40),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_151),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_15),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_103),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_59),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_33),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_12),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_15),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_38),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_22),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_13),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_80),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_58),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_43),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_5),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_45),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_20),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_141),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_63),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_116),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_48),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_52),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_148),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_99),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_61),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_68),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_20),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_135),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_5),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_75),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_74),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_69),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_134),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_73),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_129),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_11),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_122),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_3),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_10),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_143),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

BUFx10_ASAP7_75t_L g271 ( 
.A(n_56),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_35),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_46),
.Y(n_273)
);

BUFx10_ASAP7_75t_L g274 ( 
.A(n_110),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_9),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_6),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_10),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_127),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_30),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_104),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_46),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_121),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_57),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_35),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_64),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_37),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_139),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_21),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_19),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_43),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_56),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_89),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_24),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_37),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_133),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_92),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_153),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_14),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_27),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_11),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_31),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_140),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_130),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_41),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_13),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_58),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_17),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_138),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_172),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_297),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_172),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_226),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_256),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_203),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_185),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_185),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_269),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_188),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_160),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_188),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_189),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_186),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_159),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_189),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_265),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_197),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_196),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_197),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_256),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g336 ( 
.A(n_293),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_200),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_164),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_200),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_166),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_157),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_204),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_204),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_212),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_256),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_220),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_167),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_223),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_242),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_223),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_265),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_232),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_224),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_232),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_280),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_174),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_175),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_176),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_253),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_253),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_264),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_178),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_180),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_264),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_286),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_166),
.Y(n_367)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_192),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_270),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_166),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_191),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_184),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_270),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_192),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_279),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_279),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g377 ( 
.A(n_230),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_256),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_187),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_224),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_199),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_289),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_191),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_157),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_289),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_295),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_230),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_201),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_378),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_378),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_380),
.A2(n_234),
.B1(n_310),
.B2(n_309),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_378),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_378),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_368),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_313),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_368),
.B(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_313),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_210),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_315),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_354),
.B(n_340),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_325),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_376),
.B(n_240),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_341),
.B(n_230),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_318),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_322),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_321),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_320),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_328),
.A2(n_211),
.B1(n_202),
.B2(n_207),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_198),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_345),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_320),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_345),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_314),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_367),
.B(n_295),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

NOR2x1_ASAP7_75t_L g421 ( 
.A(n_323),
.B(n_157),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_329),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_326),
.B(n_237),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_345),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_333),
.Y(n_426)
);

INVxp33_ASAP7_75t_SL g427 ( 
.A(n_338),
.Y(n_427)
);

AND3x2_ASAP7_75t_L g428 ( 
.A(n_331),
.B(n_170),
.C(n_278),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_347),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_327),
.Y(n_432)
);

NOR2xp67_ASAP7_75t_L g433 ( 
.A(n_327),
.B(n_173),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_357),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_330),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_330),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_370),
.B(n_237),
.Y(n_437)
);

CKINVDCx11_ASAP7_75t_R g438 ( 
.A(n_316),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_336),
.A2(n_268),
.B1(n_222),
.B2(n_306),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_317),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_324),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_335),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_335),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_332),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_332),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_334),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_334),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_337),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g451 ( 
.A(n_358),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_339),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_359),
.B(n_298),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_377),
.B(n_298),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_363),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_387),
.B(n_237),
.Y(n_457)
);

OR2x6_ASAP7_75t_L g458 ( 
.A(n_451),
.B(n_413),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_431),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_451),
.B(n_376),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_403),
.B(n_372),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_404),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_379),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_447),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_381),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_403),
.B(n_388),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_389),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_447),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_455),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_430),
.B(n_371),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_447),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_390),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_406),
.B(n_384),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_449),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_397),
.B(n_407),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

OAI22x1_ASAP7_75t_L g485 ( 
.A1(n_439),
.A2(n_383),
.B1(n_213),
.B2(n_292),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_456),
.B(n_374),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_427),
.B(n_375),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_396),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_449),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_408),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_449),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_397),
.B(n_339),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_449),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_397),
.B(n_342),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_449),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_391),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_393),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g498 ( 
.A1(n_398),
.A2(n_386),
.B1(n_385),
.B2(n_382),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_393),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_419),
.B(n_342),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_395),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_450),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_395),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_450),
.Y(n_505)
);

BUFx10_ASAP7_75t_L g506 ( 
.A(n_423),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_440),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_392),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_L g509 ( 
.A1(n_421),
.A2(n_424),
.B1(n_407),
.B2(n_414),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_410),
.B(n_240),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_429),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_429),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_437),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_407),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_429),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_418),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_429),
.Y(n_518)
);

INVx4_ASAP7_75t_L g519 ( 
.A(n_450),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_454),
.B(n_343),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_425),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_SL g522 ( 
.A1(n_399),
.A2(n_346),
.B(n_343),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_407),
.B(n_346),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_421),
.A2(n_386),
.B1(n_385),
.B2(n_382),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_424),
.A2(n_373),
.B1(n_369),
.B2(n_365),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_399),
.B(n_348),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_438),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_414),
.B(n_348),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_440),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_400),
.B(n_349),
.Y(n_530)
);

AND3x2_ASAP7_75t_L g531 ( 
.A(n_437),
.B(n_278),
.C(n_209),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_440),
.Y(n_533)
);

CKINVDCx6p67_ASAP7_75t_R g534 ( 
.A(n_401),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_401),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_400),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_457),
.B(n_349),
.Y(n_537)
);

OR2x6_ASAP7_75t_L g538 ( 
.A(n_457),
.B(n_351),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_402),
.A2(n_250),
.B1(n_238),
.B2(n_236),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_445),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_446),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_424),
.B(n_351),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_446),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_446),
.Y(n_545)
);

AND2x4_ASAP7_75t_L g546 ( 
.A(n_424),
.B(n_353),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_442),
.Y(n_547)
);

OAI21xp33_ASAP7_75t_SL g548 ( 
.A1(n_402),
.A2(n_355),
.B(n_353),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_405),
.B(n_355),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_452),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_405),
.B(n_360),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx1_ASAP7_75t_SL g553 ( 
.A(n_428),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_442),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_411),
.B(n_360),
.Y(n_555)
);

AND3x1_ASAP7_75t_L g556 ( 
.A(n_411),
.B(n_209),
.C(n_198),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_452),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_442),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_443),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_412),
.B(n_361),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_429),
.Y(n_561)
);

INVx5_ASAP7_75t_L g562 ( 
.A(n_401),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_412),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g564 ( 
.A(n_416),
.B(n_361),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_443),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_416),
.B(n_420),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_420),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_443),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_429),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_422),
.B(n_432),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_422),
.B(n_362),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_432),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_444),
.Y(n_573)
);

NAND2xp33_ASAP7_75t_L g574 ( 
.A(n_435),
.B(n_362),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_425),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_435),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_425),
.Y(n_577)
);

BUFx4f_ASAP7_75t_L g578 ( 
.A(n_401),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_436),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_401),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_436),
.B(n_365),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_441),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_401),
.A2(n_373),
.B1(n_369),
.B2(n_278),
.Y(n_583)
);

AND3x2_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_239),
.C(n_216),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_401),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_441),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_448),
.B(n_239),
.C(n_216),
.Y(n_587)
);

BUFx8_ASAP7_75t_SL g588 ( 
.A(n_441),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_441),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_433),
.B(n_243),
.Y(n_590)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_433),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_444),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_444),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_444),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_394),
.Y(n_595)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_394),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_394),
.B(n_248),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_394),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_394),
.Y(n_601)
);

INVx11_ASAP7_75t_L g602 ( 
.A(n_409),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_409),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_409),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_475),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_475),
.B(n_483),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_556),
.B(n_210),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_501),
.B(n_182),
.Y(n_608)
);

AND2x4_ASAP7_75t_SL g609 ( 
.A(n_459),
.B(n_344),
.Y(n_609)
);

AOI22x1_ASAP7_75t_L g610 ( 
.A1(n_519),
.A2(n_244),
.B1(n_275),
.B2(n_291),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_556),
.B(n_210),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_520),
.B(n_182),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_483),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_467),
.B(n_572),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_572),
.B(n_272),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_507),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_507),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_519),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_576),
.B(n_272),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_513),
.B(n_225),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_472),
.B(n_227),
.Y(n_621)
);

INVx4_ASAP7_75t_L g622 ( 
.A(n_602),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_536),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_519),
.B(n_173),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_494),
.B(n_282),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_529),
.Y(n_626)
);

O2A1O1Ixp5_ASAP7_75t_L g627 ( 
.A1(n_570),
.A2(n_282),
.B(n_303),
.C(n_244),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_536),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_459),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_578),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_536),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_538),
.A2(n_274),
.B1(n_257),
.B2(n_240),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_472),
.B(n_231),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g634 ( 
.A(n_464),
.B(n_356),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_494),
.B(n_284),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_494),
.B(n_284),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_488),
.B(n_490),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_529),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_500),
.Y(n_639)
);

INVxp67_ASAP7_75t_SL g640 ( 
.A(n_514),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_472),
.B(n_235),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_538),
.A2(n_485),
.B1(n_509),
.B2(n_514),
.Y(n_642)
);

OAI221xp5_ASAP7_75t_L g643 ( 
.A1(n_498),
.A2(n_291),
.B1(n_275),
.B2(n_285),
.C(n_308),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_533),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_538),
.A2(n_251),
.B1(n_312),
.B2(n_252),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_538),
.A2(n_251),
.B1(n_254),
.B2(n_190),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_519),
.B(n_229),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_578),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_494),
.B(n_284),
.Y(n_649)
);

AO221x1_ASAP7_75t_L g650 ( 
.A1(n_485),
.A2(n_303),
.B1(n_267),
.B2(n_296),
.C(n_245),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_500),
.Y(n_651)
);

NAND2xp33_ASAP7_75t_L g652 ( 
.A(n_474),
.B(n_241),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_578),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_510),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_566),
.A2(n_417),
.B(n_415),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_591),
.B(n_249),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_538),
.A2(n_277),
.B1(n_276),
.B2(n_290),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_547),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_506),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_535),
.B(n_229),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_504),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g663 ( 
.A(n_459),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_504),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_563),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_546),
.B(n_549),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_563),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_546),
.B(n_285),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_459),
.B(n_243),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_461),
.B(n_273),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_567),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_560),
.B(n_296),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_469),
.B(n_288),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_528),
.B(n_294),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_537),
.B(n_304),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_581),
.B(n_304),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_492),
.B(n_308),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_506),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_525),
.B(n_301),
.Y(n_679)
);

NAND3xp33_ASAP7_75t_L g680 ( 
.A(n_463),
.B(n_302),
.C(n_229),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_535),
.B(n_169),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_SL g682 ( 
.A(n_486),
.B(n_366),
.C(n_161),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_567),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_506),
.B(n_243),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_579),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_L g686 ( 
.A(n_505),
.B(n_409),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_579),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_574),
.A2(n_233),
.B1(n_162),
.B2(n_163),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_535),
.B(n_169),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_158),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_503),
.B(n_258),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_480),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_505),
.Y(n_693)
);

INVx4_ASAP7_75t_L g694 ( 
.A(n_602),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_564),
.B(n_165),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_503),
.B(n_258),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_482),
.A2(n_193),
.B1(n_195),
.B2(n_218),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_503),
.B(n_258),
.Y(n_698)
);

INVxp33_ASAP7_75t_L g699 ( 
.A(n_487),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_564),
.B(n_168),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_462),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_460),
.B(n_271),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_524),
.B(n_171),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_517),
.B(n_271),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_517),
.B(n_177),
.Y(n_705)
);

INVx8_ASAP7_75t_L g706 ( 
.A(n_458),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_458),
.A2(n_179),
.B1(n_181),
.B2(n_183),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_458),
.B(n_271),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_532),
.A2(n_274),
.B1(n_257),
.B2(n_271),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_470),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_598),
.A2(n_417),
.B(n_415),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_517),
.B(n_194),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_535),
.B(n_193),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_547),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_516),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_473),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_580),
.B(n_409),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_473),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_526),
.B(n_205),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_532),
.A2(n_257),
.B1(n_274),
.B2(n_311),
.Y(n_720)
);

NAND2xp33_ASAP7_75t_L g721 ( 
.A(n_476),
.B(n_478),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_543),
.B(n_311),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_580),
.B(n_409),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_479),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_479),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_590),
.B(n_311),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_530),
.B(n_206),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_571),
.B(n_208),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_489),
.B(n_311),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_497),
.B(n_214),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_497),
.B(n_502),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_554),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_458),
.A2(n_502),
.B1(n_551),
.B2(n_555),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_489),
.B(n_0),
.Y(n_734)
);

BUFx3_ASAP7_75t_L g735 ( 
.A(n_603),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_558),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_489),
.B(n_1),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_458),
.A2(n_195),
.B1(n_218),
.B2(n_246),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_580),
.B(n_415),
.Y(n_739)
);

BUFx6f_ASAP7_75t_SL g740 ( 
.A(n_527),
.Y(n_740)
);

INVx4_ASAP7_75t_L g741 ( 
.A(n_580),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_540),
.B(n_215),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_540),
.B(n_217),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_558),
.Y(n_744)
);

NOR2xp67_ASAP7_75t_L g745 ( 
.A(n_522),
.B(n_219),
.Y(n_745)
);

OR2x2_ASAP7_75t_L g746 ( 
.A(n_553),
.B(n_1),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_541),
.B(n_221),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_508),
.B(n_257),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_541),
.B(n_228),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_559),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_522),
.B(n_247),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_SL g752 ( 
.A(n_548),
.B(n_255),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_559),
.Y(n_753)
);

OAI22xp5_ASAP7_75t_L g754 ( 
.A1(n_542),
.A2(n_195),
.B1(n_218),
.B2(n_246),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_601),
.A2(n_417),
.B(n_415),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_542),
.B(n_259),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_548),
.B(n_261),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_489),
.B(n_8),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_539),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_508),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_544),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_465),
.A2(n_417),
.B(n_415),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_544),
.B(n_283),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_545),
.A2(n_550),
.B(n_552),
.C(n_557),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_545),
.B(n_281),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_476),
.B(n_9),
.Y(n_766)
);

INVx1_ASAP7_75t_SL g767 ( 
.A(n_588),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_476),
.B(n_12),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_565),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_531),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_665),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_630),
.Y(n_772)
);

AND2x6_ASAP7_75t_SL g773 ( 
.A(n_740),
.B(n_748),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_629),
.B(n_585),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_667),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_692),
.B(n_476),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_607),
.A2(n_552),
.B1(n_557),
.B2(n_550),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_629),
.B(n_585),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_630),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_616),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_606),
.B(n_584),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_671),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_614),
.B(n_589),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_605),
.B(n_587),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_683),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_613),
.B(n_583),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_666),
.B(n_589),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_663),
.B(n_660),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_608),
.B(n_478),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_630),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_685),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_612),
.B(n_478),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_622),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_759),
.A2(n_478),
.B(n_495),
.C(n_468),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_611),
.A2(n_585),
.B1(n_495),
.B2(n_534),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_611),
.A2(n_495),
.B1(n_534),
.B2(n_465),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_687),
.Y(n_797)
);

NOR2x2_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_582),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_639),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_619),
.B(n_495),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_663),
.B(n_562),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_651),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_650),
.A2(n_565),
.B1(n_568),
.B2(n_499),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_701),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_740),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_662),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_655),
.B(n_596),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_741),
.B(n_604),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_616),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_664),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_634),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_693),
.Y(n_812)
);

NOR2x2_ASAP7_75t_L g813 ( 
.A(n_609),
.B(n_586),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_630),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_648),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_648),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_637),
.Y(n_817)
);

AO22x1_ASAP7_75t_L g818 ( 
.A1(n_708),
.A2(n_562),
.B1(n_260),
.B2(n_246),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_621),
.B(n_586),
.Y(n_819)
);

INVx5_ASAP7_75t_L g820 ( 
.A(n_648),
.Y(n_820)
);

NOR2x2_ASAP7_75t_L g821 ( 
.A(n_609),
.B(n_592),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_760),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_648),
.Y(n_823)
);

AND3x2_ASAP7_75t_SL g824 ( 
.A(n_706),
.B(n_592),
.C(n_274),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_699),
.B(n_466),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_617),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_746),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_721),
.A2(n_624),
.B(n_731),
.Y(n_828)
);

INVx3_ASAP7_75t_L g829 ( 
.A(n_654),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_617),
.Y(n_830)
);

NOR2x2_ASAP7_75t_L g831 ( 
.A(n_707),
.B(n_652),
.Y(n_831)
);

INVx2_ASAP7_75t_SL g832 ( 
.A(n_706),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_626),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_620),
.B(n_599),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_678),
.B(n_562),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_654),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_621),
.B(n_466),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_654),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_633),
.B(n_468),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_633),
.B(n_471),
.Y(n_840)
);

INVxp67_ASAP7_75t_L g841 ( 
.A(n_641),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_623),
.A2(n_493),
.B1(n_491),
.B2(n_481),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_625),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_741),
.B(n_604),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_641),
.A2(n_493),
.B1(n_491),
.B2(n_477),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_695),
.B(n_471),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_770),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_620),
.B(n_484),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_654),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_733),
.B(n_477),
.Y(n_850)
);

NOR3xp33_ASAP7_75t_SL g851 ( 
.A(n_682),
.B(n_300),
.C(n_262),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_767),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_626),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_618),
.B(n_604),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_638),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_657),
.B(n_674),
.Y(n_856)
);

NOR2x1_ASAP7_75t_L g857 ( 
.A(n_680),
.B(n_603),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_638),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_642),
.A2(n_568),
.B1(n_521),
.B2(n_575),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_644),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_761),
.Y(n_861)
);

INVx5_ASAP7_75t_L g862 ( 
.A(n_618),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_657),
.Y(n_863)
);

INVx2_ASAP7_75t_SL g864 ( 
.A(n_706),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_710),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_644),
.Y(n_866)
);

BUFx4f_ASAP7_75t_L g867 ( 
.A(n_675),
.Y(n_867)
);

OR2x6_ASAP7_75t_L g868 ( 
.A(n_622),
.B(n_481),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_SL g869 ( 
.A(n_645),
.B(n_287),
.C(n_266),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_675),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_653),
.Y(n_871)
);

BUFx4f_ASAP7_75t_L g872 ( 
.A(n_675),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_694),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_716),
.Y(n_874)
);

AND3x2_ASAP7_75t_SL g875 ( 
.A(n_738),
.B(n_484),
.C(n_496),
.Y(n_875)
);

INVxp67_ASAP7_75t_L g876 ( 
.A(n_674),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_694),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_670),
.B(n_511),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_670),
.B(n_511),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_735),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_673),
.B(n_511),
.Y(n_881)
);

INVx5_ASAP7_75t_L g882 ( 
.A(n_735),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_691),
.A2(n_593),
.B1(n_600),
.B2(n_594),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_653),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_718),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_702),
.B(n_673),
.Y(n_886)
);

BUFx8_ASAP7_75t_L g887 ( 
.A(n_628),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_724),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_631),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_R g890 ( 
.A(n_691),
.B(n_562),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_684),
.B(n_669),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_745),
.B(n_604),
.Y(n_892)
);

AND2x6_ASAP7_75t_SL g893 ( 
.A(n_726),
.B(n_600),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_734),
.A2(n_518),
.B(n_561),
.C(n_515),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_659),
.Y(n_895)
);

NAND2x1_ASAP7_75t_L g896 ( 
.A(n_725),
.B(n_511),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_658),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_700),
.B(n_496),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_659),
.Y(n_899)
);

NOR3xp33_ASAP7_75t_SL g900 ( 
.A(n_751),
.B(n_757),
.C(n_752),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_696),
.B(n_496),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_734),
.B(n_604),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_696),
.B(n_499),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_714),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_737),
.B(n_604),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_698),
.B(n_499),
.Y(n_906)
);

NOR3xp33_ASAP7_75t_SL g907 ( 
.A(n_737),
.B(n_758),
.C(n_766),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_668),
.B(n_562),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_640),
.A2(n_515),
.B1(n_569),
.B2(n_512),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_714),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_698),
.B(n_521),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_732),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_732),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_722),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_704),
.B(n_521),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_758),
.B(n_512),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_704),
.B(n_575),
.Y(n_917)
);

OR2x2_ASAP7_75t_SL g918 ( 
.A(n_679),
.B(n_594),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_646),
.B(n_263),
.C(n_299),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_672),
.B(n_575),
.Y(n_920)
);

INVx5_ASAP7_75t_L g921 ( 
.A(n_736),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_635),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_736),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_676),
.B(n_577),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_615),
.B(n_577),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_764),
.B(n_561),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_744),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_744),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_729),
.B(n_577),
.Y(n_929)
);

NOR3xp33_ASAP7_75t_SL g930 ( 
.A(n_766),
.B(n_305),
.C(n_307),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_647),
.A2(n_597),
.B(n_561),
.Y(n_931)
);

BUFx6f_ASAP7_75t_SL g932 ( 
.A(n_643),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_769),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_750),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_750),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_753),
.Y(n_936)
);

BUFx4f_ASAP7_75t_L g937 ( 
.A(n_753),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_729),
.B(n_569),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_769),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_677),
.B(n_569),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_722),
.B(n_561),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_636),
.B(n_573),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_649),
.B(n_562),
.Y(n_943)
);

BUFx8_ASAP7_75t_L g944 ( 
.A(n_726),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_632),
.A2(n_593),
.B1(n_597),
.B2(n_512),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_705),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_627),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_688),
.A2(n_719),
.B1(n_727),
.B2(n_728),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_610),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_690),
.B(n_518),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_703),
.B(n_573),
.Y(n_951)
);

AND3x1_ASAP7_75t_SL g952 ( 
.A(n_768),
.B(n_14),
.C(n_16),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_712),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_856),
.A2(n_768),
.B1(n_647),
.B2(n_624),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_856),
.B(n_709),
.Y(n_955)
);

OAI21x1_ASAP7_75t_L g956 ( 
.A1(n_828),
.A2(n_762),
.B(n_656),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_938),
.A2(n_739),
.B(n_717),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_929),
.A2(n_723),
.B(n_739),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_841),
.A2(n_730),
.B(n_765),
.C(n_756),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_771),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_931),
.A2(n_755),
.B(n_711),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_876),
.B(n_720),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_902),
.A2(n_905),
.B(n_839),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_914),
.B(n_742),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_863),
.B(n_897),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_907),
.A2(n_763),
.B(n_743),
.C(n_749),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_880),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_902),
.A2(n_723),
.B(n_686),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_775),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_SL g970 ( 
.A1(n_822),
.A2(n_697),
.B1(n_754),
.B2(n_260),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_805),
.Y(n_971)
);

AND2x2_ASAP7_75t_SL g972 ( 
.A(n_867),
.B(n_747),
.Y(n_972)
);

AOI22xp5_ASAP7_75t_L g973 ( 
.A1(n_932),
.A2(n_661),
.B1(n_689),
.B2(n_681),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_870),
.B(n_661),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_804),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_907),
.A2(n_713),
.B(n_689),
.C(n_681),
.Y(n_976)
);

AOI222xp33_ASAP7_75t_L g977 ( 
.A1(n_932),
.A2(n_260),
.B1(n_713),
.B2(n_603),
.C1(n_415),
.C2(n_417),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_817),
.B(n_573),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_867),
.B(n_595),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_782),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_905),
.A2(n_573),
.B(n_569),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_886),
.B(n_518),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_837),
.A2(n_518),
.B(n_515),
.Y(n_983)
);

NAND2x1_ASAP7_75t_L g984 ( 
.A(n_779),
.B(n_515),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_848),
.B(n_512),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_780),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_785),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_R g988 ( 
.A(n_930),
.B(n_66),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_SL g989 ( 
.A(n_869),
.B(n_16),
.C(n_22),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_850),
.A2(n_417),
.B1(n_25),
.B2(n_26),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_840),
.A2(n_879),
.B(n_878),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_880),
.Y(n_992)
);

AOI22xp33_ASAP7_75t_L g993 ( 
.A1(n_872),
.A2(n_595),
.B1(n_28),
.B2(n_29),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_878),
.A2(n_595),
.B(n_76),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_817),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_811),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_879),
.A2(n_67),
.B(n_149),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_872),
.B(n_774),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_834),
.A2(n_23),
.B(n_28),
.C(n_29),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_881),
.A2(n_903),
.B(n_901),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_919),
.A2(n_776),
.B(n_819),
.C(n_783),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_881),
.A2(n_77),
.B(n_144),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_786),
.B(n_32),
.Y(n_1003)
);

O2A1O1Ixp5_ASAP7_75t_L g1004 ( 
.A1(n_916),
.A2(n_32),
.B(n_34),
.C(n_36),
.Y(n_1004)
);

INVxp67_ASAP7_75t_L g1005 ( 
.A(n_811),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_804),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_L g1007 ( 
.A1(n_916),
.A2(n_36),
.B(n_39),
.C(n_41),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_791),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_797),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_799),
.Y(n_1010)
);

NAND2x1_ASAP7_75t_SL g1011 ( 
.A(n_781),
.B(n_39),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_843),
.B(n_42),
.Y(n_1012)
);

OAI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_894),
.A2(n_42),
.B(n_44),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_944),
.B(n_44),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_802),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_806),
.Y(n_1016)
);

O2A1O1Ixp5_ASAP7_75t_L g1017 ( 
.A1(n_892),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_847),
.B(n_51),
.Y(n_1018)
);

OA22x2_ASAP7_75t_L g1019 ( 
.A1(n_827),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_810),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_SL g1021 ( 
.A1(n_776),
.A2(n_53),
.B(n_60),
.C(n_65),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_906),
.A2(n_79),
.B(n_82),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_882),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_784),
.A2(n_84),
.B1(n_96),
.B2(n_97),
.Y(n_1024)
);

OAI22x1_ASAP7_75t_L g1025 ( 
.A1(n_891),
.A2(n_100),
.B1(n_101),
.B2(n_106),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_812),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_787),
.B(n_119),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_843),
.B(n_120),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_882),
.Y(n_1029)
);

INVx3_ASAP7_75t_SL g1030 ( 
.A(n_813),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_911),
.A2(n_126),
.B(n_128),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_944),
.B(n_142),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_894),
.A2(n_154),
.B(n_846),
.C(n_794),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_780),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_861),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_882),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_948),
.A2(n_949),
.B(n_877),
.C(n_873),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_798),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_915),
.A2(n_917),
.B(n_950),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_854),
.A2(n_898),
.B(n_792),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_854),
.A2(n_789),
.B(n_844),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_926),
.A2(n_800),
.B(n_922),
.C(n_940),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_772),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_808),
.A2(n_844),
.B(n_926),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_850),
.B(n_777),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_825),
.B(n_922),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_SL g1047 ( 
.A1(n_852),
.A2(n_831),
.B1(n_891),
.B2(n_864),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_930),
.A2(n_900),
.B(n_946),
.C(n_953),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_809),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_777),
.B(n_920),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_773),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_851),
.B(n_900),
.C(n_883),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_SL g1053 ( 
.A1(n_831),
.A2(n_832),
.B1(n_788),
.B2(n_825),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_946),
.A2(n_953),
.B(n_851),
.C(n_942),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_924),
.B(n_865),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_788),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_807),
.B(n_874),
.Y(n_1057)
);

AOI22x1_ASAP7_75t_L g1058 ( 
.A1(n_947),
.A2(n_877),
.B1(n_873),
.B2(n_941),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_807),
.B(n_885),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_887),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_888),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_845),
.A2(n_796),
.B1(n_868),
.B2(n_862),
.Y(n_1062)
);

AND2x6_ASAP7_75t_L g1063 ( 
.A(n_774),
.B(n_778),
.Y(n_1063)
);

INVx2_ASAP7_75t_SL g1064 ( 
.A(n_887),
.Y(n_1064)
);

BUFx10_ASAP7_75t_L g1065 ( 
.A(n_893),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_772),
.Y(n_1066)
);

NAND3xp33_ASAP7_75t_SL g1067 ( 
.A(n_952),
.B(n_890),
.C(n_803),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_809),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_868),
.A2(n_862),
.B1(n_795),
.B2(n_937),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_808),
.A2(n_892),
.B(n_909),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_772),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_951),
.A2(n_842),
.B(n_925),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_826),
.B(n_860),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_826),
.B(n_860),
.Y(n_1075)
);

AO32x1_ASAP7_75t_L g1076 ( 
.A1(n_952),
.A2(n_935),
.A3(n_939),
.B1(n_936),
.B2(n_904),
.Y(n_1076)
);

OA22x2_ASAP7_75t_L g1077 ( 
.A1(n_798),
.A2(n_945),
.B1(n_813),
.B2(n_821),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_937),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_830),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_801),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_830),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_889),
.B(n_918),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_833),
.Y(n_1083)
);

NOR3xp33_ASAP7_75t_SL g1084 ( 
.A(n_951),
.B(n_824),
.C(n_821),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_833),
.B(n_866),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_L g1086 ( 
.A1(n_868),
.A2(n_803),
.B(n_889),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_793),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_853),
.B(n_910),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_772),
.Y(n_1089)
);

BUFx6f_ASAP7_75t_L g1090 ( 
.A(n_814),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_801),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_896),
.A2(n_862),
.B(n_921),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_779),
.A2(n_790),
.B(n_838),
.C(n_815),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_857),
.A2(n_818),
.B(n_936),
.Y(n_1094)
);

AND2x6_ASAP7_75t_SL g1095 ( 
.A(n_835),
.B(n_824),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_862),
.A2(n_921),
.B(n_934),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1045),
.B(n_899),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_991),
.A2(n_921),
.B(n_820),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_SL g1099 ( 
.A(n_971),
.B(n_820),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_956),
.A2(n_866),
.B(n_927),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1000),
.A2(n_1039),
.B(n_1073),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_986),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1045),
.B(n_928),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_955),
.B(n_910),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_972),
.B(n_820),
.Y(n_1105)
);

AOI21x1_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_871),
.B(n_927),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_995),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_969),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1034),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_962),
.A2(n_908),
.B(n_790),
.C(n_815),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_961),
.A2(n_855),
.B(n_912),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_SL g1112 ( 
.A1(n_1037),
.A2(n_816),
.B(n_849),
.C(n_829),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_964),
.A2(n_836),
.B(n_816),
.C(n_849),
.Y(n_1113)
);

AOI21x1_ASAP7_75t_L g1114 ( 
.A1(n_1070),
.A2(n_871),
.B(n_913),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_975),
.Y(n_1115)
);

OAI22x1_ASAP7_75t_L g1116 ( 
.A1(n_1038),
.A2(n_965),
.B1(n_1030),
.B2(n_1082),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1040),
.A2(n_1058),
.B(n_1044),
.Y(n_1117)
);

CKINVDCx11_ASAP7_75t_R g1118 ( 
.A(n_1060),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1051),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_1041),
.A2(n_855),
.B(n_912),
.Y(n_1120)
);

OAI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_954),
.A2(n_859),
.B(n_943),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1094),
.A2(n_884),
.B(n_913),
.Y(n_1122)
);

AOI21xp33_ASAP7_75t_L g1123 ( 
.A1(n_990),
.A2(n_875),
.B(n_859),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_967),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1055),
.B(n_884),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_954),
.A2(n_994),
.B(n_1027),
.Y(n_1126)
);

AND2x2_ASAP7_75t_L g1127 ( 
.A(n_996),
.B(n_1005),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_1006),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_1027),
.A2(n_1001),
.B(n_966),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1050),
.A2(n_858),
.A3(n_875),
.B(n_933),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_1053),
.B(n_836),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_1062),
.A2(n_858),
.A3(n_933),
.B(n_921),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_958),
.A2(n_890),
.B(n_933),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_1087),
.Y(n_1134)
);

NOR4xp25_ASAP7_75t_L g1135 ( 
.A(n_990),
.B(n_895),
.C(n_829),
.D(n_838),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_1080),
.B(n_835),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1055),
.B(n_895),
.Y(n_1137)
);

AO31x2_ASAP7_75t_L g1138 ( 
.A1(n_1062),
.A2(n_933),
.A3(n_943),
.B(n_814),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_983),
.A2(n_814),
.B(n_823),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_981),
.A2(n_814),
.B(n_823),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_SL g1141 ( 
.A1(n_1013),
.A2(n_823),
.B(n_1048),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_1057),
.B(n_823),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_957),
.A2(n_1033),
.B(n_959),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1065),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_1059),
.B(n_967),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_998),
.B(n_1077),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_1003),
.B(n_1046),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_1074),
.A2(n_1088),
.A3(n_1075),
.B(n_1085),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_L g1149 ( 
.A(n_999),
.B(n_989),
.C(n_1013),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1091),
.B(n_1063),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_967),
.Y(n_1151)
);

INVxp67_ASAP7_75t_L g1152 ( 
.A(n_1018),
.Y(n_1152)
);

O2A1O1Ixp5_ASAP7_75t_L g1153 ( 
.A1(n_997),
.A2(n_1002),
.B(n_979),
.C(n_968),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_976),
.A2(n_1069),
.B(n_985),
.Y(n_1154)
);

NAND3xp33_ASAP7_75t_SL g1155 ( 
.A(n_1014),
.B(n_1054),
.C(n_993),
.Y(n_1155)
);

AOI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1096),
.A2(n_1092),
.B(n_985),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1049),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1042),
.A2(n_1067),
.B(n_982),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1022),
.A2(n_1031),
.B(n_984),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1052),
.A2(n_1028),
.B(n_1021),
.Y(n_1160)
);

NAND3xp33_ASAP7_75t_L g1161 ( 
.A(n_1084),
.B(n_1007),
.C(n_1004),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1063),
.B(n_980),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1093),
.A2(n_1076),
.B(n_1075),
.Y(n_1163)
);

OR2x2_ASAP7_75t_L g1164 ( 
.A(n_1047),
.B(n_1012),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1063),
.B(n_987),
.Y(n_1165)
);

BUFx3_ASAP7_75t_L g1166 ( 
.A(n_992),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1068),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1017),
.A2(n_973),
.B(n_978),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1008),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1064),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_992),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1063),
.B(n_1009),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1074),
.A2(n_1085),
.A3(n_1088),
.B(n_1079),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1010),
.B(n_1015),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1086),
.B(n_1032),
.Y(n_1175)
);

OR2x2_ASAP7_75t_L g1176 ( 
.A(n_1016),
.B(n_1035),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_974),
.A2(n_1020),
.B(n_1026),
.Y(n_1177)
);

INVx2_ASAP7_75t_SL g1178 ( 
.A(n_992),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_970),
.B(n_1065),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1072),
.A2(n_1083),
.B(n_1081),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1025),
.A2(n_1061),
.B(n_1077),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1091),
.B(n_1078),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_1023),
.Y(n_1183)
);

OAI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1019),
.A2(n_1024),
.B1(n_1029),
.B2(n_1036),
.Y(n_1184)
);

INVx4_ASAP7_75t_L g1185 ( 
.A(n_1023),
.Y(n_1185)
);

OA21x2_ASAP7_75t_L g1186 ( 
.A1(n_1076),
.A2(n_1011),
.B(n_977),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_977),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1023),
.A2(n_1036),
.B(n_1090),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1043),
.B(n_1090),
.Y(n_1189)
);

AO22x2_ASAP7_75t_L g1190 ( 
.A1(n_1095),
.A2(n_1019),
.B1(n_988),
.B2(n_1056),
.Y(n_1190)
);

INVx6_ASAP7_75t_L g1191 ( 
.A(n_1036),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_R g1192 ( 
.A(n_1043),
.B(n_1066),
.Y(n_1192)
);

AO31x2_ASAP7_75t_L g1193 ( 
.A1(n_1043),
.A2(n_1066),
.A3(n_1071),
.B(n_1089),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1071),
.A2(n_1089),
.B(n_1090),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1089),
.A2(n_956),
.B(n_961),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_995),
.B(n_606),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_955),
.B(n_605),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_960),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_972),
.B(n_856),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1037),
.A2(n_856),
.B(n_841),
.C(n_966),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_995),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_972),
.B(n_856),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1045),
.A2(n_856),
.B(n_1050),
.Y(n_1206)
);

NOR4xp25_ASAP7_75t_L g1207 ( 
.A(n_990),
.B(n_999),
.C(n_955),
.D(n_1013),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_960),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_986),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_955),
.A2(n_856),
.B(n_876),
.C(n_841),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_956),
.A2(n_961),
.B(n_1040),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_956),
.A2(n_961),
.B(n_1040),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_995),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_955),
.A2(n_856),
.B(n_876),
.C(n_841),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_975),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_SL g1218 ( 
.A1(n_964),
.A2(n_467),
.B(n_856),
.C(n_737),
.Y(n_1218)
);

NOR2xp33_ASAP7_75t_L g1219 ( 
.A(n_955),
.B(n_474),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1220)
);

CKINVDCx11_ASAP7_75t_R g1221 ( 
.A(n_1060),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1005),
.B(n_474),
.Y(n_1222)
);

O2A1O1Ixp5_ASAP7_75t_SL g1223 ( 
.A1(n_990),
.A2(n_892),
.B(n_905),
.C(n_902),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_SL g1224 ( 
.A(n_972),
.B(n_856),
.Y(n_1224)
);

AND2x4_ASAP7_75t_L g1225 ( 
.A(n_1080),
.B(n_1091),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_960),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_991),
.A2(n_907),
.B(n_856),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_1080),
.B(n_1091),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_971),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1045),
.B(n_1055),
.Y(n_1230)
);

INVx5_ASAP7_75t_L g1231 ( 
.A(n_1063),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_956),
.A2(n_961),
.B(n_1040),
.Y(n_1232)
);

O2A1O1Ixp5_ASAP7_75t_L g1233 ( 
.A1(n_955),
.A2(n_856),
.B(n_991),
.C(n_954),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_991),
.A2(n_907),
.B(n_856),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_960),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1080),
.B(n_1091),
.Y(n_1238)
);

OA21x2_ASAP7_75t_L g1239 ( 
.A1(n_963),
.A2(n_956),
.B(n_991),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1240)
);

O2A1O1Ixp5_ASAP7_75t_L g1241 ( 
.A1(n_955),
.A2(n_856),
.B(n_991),
.C(n_954),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_991),
.A2(n_1000),
.B(n_1039),
.Y(n_1242)
);

NAND3x1_ASAP7_75t_L g1243 ( 
.A(n_1014),
.B(n_1032),
.C(n_856),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1197),
.B(n_1219),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1126),
.A2(n_1101),
.B(n_1233),
.Y(n_1245)
);

OA21x2_ASAP7_75t_L g1246 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1241),
.A2(n_1209),
.B(n_1200),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1195),
.A2(n_1117),
.B(n_1114),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1174),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1159),
.A2(n_1236),
.B(n_1234),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1174),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1123),
.A2(n_1149),
.B1(n_1164),
.B2(n_1155),
.Y(n_1252)
);

INVx1_ASAP7_75t_SL g1253 ( 
.A(n_1134),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1123),
.A2(n_1175),
.B1(n_1190),
.B2(n_1198),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1240),
.A2(n_1242),
.B(n_1106),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1154),
.A2(n_1143),
.A3(n_1097),
.B(n_1103),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1156),
.A2(n_1100),
.B(n_1111),
.Y(n_1257)
);

AND2x4_ASAP7_75t_L g1258 ( 
.A(n_1231),
.B(n_1150),
.Y(n_1258)
);

OAI21x1_ASAP7_75t_L g1259 ( 
.A1(n_1120),
.A2(n_1139),
.B(n_1133),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1212),
.A2(n_1216),
.B(n_1235),
.Y(n_1260)
);

AND2x4_ASAP7_75t_L g1261 ( 
.A(n_1231),
.B(n_1150),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1108),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_1146),
.B(n_1206),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1121),
.A2(n_1227),
.B(n_1158),
.C(n_1218),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1122),
.A2(n_1153),
.B(n_1140),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1121),
.A2(n_1158),
.B(n_1168),
.C(n_1160),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1169),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1207),
.B(n_1202),
.C(n_1175),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1231),
.B(n_1194),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1243),
.A2(n_1179),
.B1(n_1190),
.B2(n_1131),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1196),
.B(n_1203),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1223),
.A2(n_1098),
.B(n_1239),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_1229),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1196),
.B(n_1203),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1211),
.B(n_1220),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1097),
.A2(n_1103),
.A3(n_1184),
.B(n_1220),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1199),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1183),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1208),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1184),
.A2(n_1211),
.A3(n_1230),
.B(n_1125),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1187),
.A2(n_1147),
.B1(n_1230),
.B2(n_1146),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1204),
.B(n_1127),
.Y(n_1282)
);

INVx5_ASAP7_75t_L g1283 ( 
.A(n_1183),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1141),
.A2(n_1180),
.B(n_1125),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1186),
.A2(n_1104),
.B1(n_1152),
.B2(n_1168),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1201),
.A2(n_1224),
.B(n_1205),
.C(n_1113),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1177),
.A2(n_1194),
.B(n_1188),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1142),
.B(n_1162),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1137),
.A2(n_1165),
.B(n_1172),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1132),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1226),
.Y(n_1291)
);

AO21x2_ASAP7_75t_L g1292 ( 
.A1(n_1135),
.A2(n_1207),
.B(n_1110),
.Y(n_1292)
);

OR2x2_ASAP7_75t_L g1293 ( 
.A(n_1237),
.B(n_1145),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1161),
.A2(n_1128),
.B1(n_1222),
.B2(n_1172),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1162),
.A2(n_1165),
.B(n_1189),
.Y(n_1295)
);

AOI222xp33_ASAP7_75t_L g1296 ( 
.A1(n_1116),
.A2(n_1170),
.B1(n_1136),
.B2(n_1221),
.C1(n_1118),
.C2(n_1238),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1102),
.A2(n_1157),
.B(n_1167),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1181),
.A2(n_1105),
.B(n_1109),
.Y(n_1298)
);

NOR2xp67_ASAP7_75t_L g1299 ( 
.A(n_1115),
.B(n_1217),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1210),
.A2(n_1186),
.B(n_1182),
.Y(n_1300)
);

CKINVDCx8_ASAP7_75t_R g1301 ( 
.A(n_1119),
.Y(n_1301)
);

AO21x2_ASAP7_75t_L g1302 ( 
.A1(n_1135),
.A2(n_1112),
.B(n_1192),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1136),
.A2(n_1238),
.B1(n_1228),
.B2(n_1225),
.Y(n_1303)
);

OA21x2_ASAP7_75t_L g1304 ( 
.A1(n_1130),
.A2(n_1148),
.B(n_1132),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1132),
.A2(n_1138),
.B(n_1193),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1130),
.A2(n_1178),
.A3(n_1124),
.B1(n_1185),
.B2(n_1138),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1183),
.A2(n_1228),
.B(n_1225),
.Y(n_1307)
);

OAI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1144),
.A2(n_1166),
.B1(n_1151),
.B2(n_1171),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1138),
.Y(n_1309)
);

OAI21xp33_ASAP7_75t_SL g1310 ( 
.A1(n_1185),
.A2(n_1099),
.B(n_1191),
.Y(n_1310)
);

BUFx6f_ASAP7_75t_L g1311 ( 
.A(n_1191),
.Y(n_1311)
);

OAI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1130),
.A2(n_856),
.B(n_1233),
.Y(n_1312)
);

INVxp67_ASAP7_75t_L g1313 ( 
.A(n_1107),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1197),
.B(n_995),
.Y(n_1314)
);

CKINVDCx6p67_ASAP7_75t_R g1315 ( 
.A(n_1118),
.Y(n_1315)
);

INVx6_ASAP7_75t_L g1316 ( 
.A(n_1231),
.Y(n_1316)
);

AO32x2_ASAP7_75t_L g1317 ( 
.A1(n_1184),
.A2(n_990),
.A3(n_1047),
.B1(n_1053),
.B2(n_954),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1219),
.A2(n_955),
.B1(n_856),
.B2(n_897),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1219),
.A2(n_856),
.B1(n_1216),
.B2(n_1212),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1176),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1123),
.A2(n_856),
.B1(n_955),
.B2(n_1019),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1233),
.A2(n_856),
.B(n_1241),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1123),
.A2(n_856),
.B1(n_955),
.B2(n_1019),
.Y(n_1324)
);

AOI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1129),
.A2(n_1143),
.B(n_1160),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1123),
.A2(n_856),
.B1(n_955),
.B2(n_1019),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1227),
.A2(n_1235),
.B(n_1141),
.Y(n_1328)
);

AO31x2_ASAP7_75t_L g1329 ( 
.A1(n_1163),
.A2(n_1126),
.A3(n_1209),
.B(n_1200),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1233),
.A2(n_856),
.B(n_1241),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1129),
.A2(n_1143),
.B(n_1160),
.Y(n_1331)
);

NOR2xp67_ASAP7_75t_L g1332 ( 
.A(n_1115),
.B(n_1217),
.Y(n_1332)
);

INVx2_ASAP7_75t_L g1333 ( 
.A(n_1173),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1197),
.B(n_995),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1335)
);

OA21x2_ASAP7_75t_L g1336 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1219),
.A2(n_955),
.B1(n_856),
.B2(n_897),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1107),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1176),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1219),
.A2(n_955),
.B1(n_856),
.B2(n_897),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1176),
.Y(n_1342)
);

BUFx3_ASAP7_75t_L g1343 ( 
.A(n_1151),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1176),
.Y(n_1344)
);

OR2x2_ASAP7_75t_L g1345 ( 
.A(n_1107),
.B(n_1215),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1219),
.A2(n_856),
.B1(n_1216),
.B2(n_1212),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1118),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1123),
.A2(n_856),
.B1(n_955),
.B2(n_1019),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_SL g1351 ( 
.A(n_1233),
.B(n_856),
.C(n_955),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1118),
.Y(n_1352)
);

OA21x2_ASAP7_75t_L g1353 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1197),
.B(n_995),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1107),
.B(n_1215),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1176),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1213),
.A2(n_1232),
.B(n_1214),
.Y(n_1359)
);

NAND2x1p5_ASAP7_75t_L g1360 ( 
.A(n_1231),
.B(n_1183),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1163),
.A2(n_1126),
.A3(n_1209),
.B(n_1200),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1318),
.A2(n_1337),
.B1(n_1341),
.B2(n_1320),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_L g1363 ( 
.A1(n_1346),
.A2(n_1351),
.B(n_1264),
.C(n_1260),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1252),
.A2(n_1268),
.B1(n_1327),
.B2(n_1348),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_SL g1365 ( 
.A1(n_1266),
.A2(n_1264),
.B(n_1351),
.Y(n_1365)
);

NOR2xp67_ASAP7_75t_L g1366 ( 
.A(n_1270),
.B(n_1283),
.Y(n_1366)
);

NOR2xp67_ASAP7_75t_L g1367 ( 
.A(n_1283),
.B(n_1310),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1334),
.B(n_1354),
.Y(n_1369)
);

BUFx12f_ASAP7_75t_L g1370 ( 
.A(n_1347),
.Y(n_1370)
);

INVxp67_ASAP7_75t_SL g1371 ( 
.A(n_1290),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1275),
.B(n_1249),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1288),
.B(n_1282),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1252),
.A2(n_1327),
.B1(n_1348),
.B2(n_1322),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1250),
.A2(n_1272),
.B(n_1255),
.Y(n_1375)
);

NOR2xp67_ASAP7_75t_L g1376 ( 
.A(n_1283),
.B(n_1313),
.Y(n_1376)
);

BUFx8_ASAP7_75t_SL g1377 ( 
.A(n_1273),
.Y(n_1377)
);

AOI211xp5_ASAP7_75t_L g1378 ( 
.A1(n_1266),
.A2(n_1294),
.B(n_1281),
.C(n_1312),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1322),
.A2(n_1324),
.B1(n_1254),
.B2(n_1323),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1324),
.A2(n_1254),
.B1(n_1330),
.B2(n_1338),
.Y(n_1380)
);

O2A1O1Ixp5_ASAP7_75t_L g1381 ( 
.A1(n_1325),
.A2(n_1331),
.B(n_1308),
.C(n_1281),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1251),
.B(n_1321),
.Y(n_1382)
);

OAI22x1_ASAP7_75t_L g1383 ( 
.A1(n_1340),
.A2(n_1342),
.B1(n_1344),
.B2(n_1358),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1313),
.B(n_1338),
.Y(n_1384)
);

OA22x2_ASAP7_75t_L g1385 ( 
.A1(n_1263),
.A2(n_1261),
.B1(n_1258),
.B2(n_1253),
.Y(n_1385)
);

OA21x2_ASAP7_75t_L g1386 ( 
.A1(n_1257),
.A2(n_1248),
.B(n_1265),
.Y(n_1386)
);

AOI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1286),
.A2(n_1302),
.B(n_1328),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1345),
.B(n_1355),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1262),
.B(n_1267),
.Y(n_1389)
);

OAI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1285),
.A2(n_1263),
.B1(n_1303),
.B2(n_1332),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1277),
.B(n_1279),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1291),
.B(n_1293),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1297),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1343),
.B(n_1280),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1308),
.B(n_1286),
.C(n_1299),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1360),
.A2(n_1258),
.B(n_1261),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1256),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_SL g1398 ( 
.A1(n_1258),
.A2(n_1261),
.B(n_1302),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1301),
.A2(n_1273),
.B1(n_1285),
.B2(n_1347),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1317),
.B(n_1303),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1297),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1269),
.B(n_1295),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1292),
.A2(n_1296),
.B(n_1278),
.C(n_1317),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1317),
.A2(n_1283),
.B1(n_1315),
.B2(n_1316),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1276),
.B(n_1292),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1317),
.B(n_1311),
.Y(n_1406)
);

OAI211xp5_ASAP7_75t_L g1407 ( 
.A1(n_1352),
.A2(n_1307),
.B(n_1289),
.C(n_1309),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1284),
.A2(n_1298),
.B(n_1287),
.C(n_1300),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_1276),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1306),
.B(n_1256),
.Y(n_1410)
);

A2O1A1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1333),
.A2(n_1259),
.B(n_1256),
.C(n_1361),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1306),
.B(n_1352),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1304),
.B(n_1361),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1329),
.A2(n_1361),
.B(n_1339),
.C(n_1349),
.Y(n_1414)
);

OAI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1246),
.A2(n_1336),
.B1(n_1357),
.B2(n_1353),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1329),
.B(n_1304),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1319),
.B(n_1350),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1336),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1326),
.B(n_1335),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1356),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1359),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1318),
.A2(n_1341),
.B1(n_1337),
.B2(n_1219),
.Y(n_1422)
);

INVx5_ASAP7_75t_L g1423 ( 
.A(n_1283),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1250),
.A2(n_1245),
.B(n_1247),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1244),
.B(n_1314),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1318),
.A2(n_1341),
.B1(n_1337),
.B2(n_1219),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1351),
.A2(n_1126),
.B(n_991),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1266),
.A2(n_856),
.B(n_955),
.C(n_1233),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1250),
.A2(n_1245),
.B(n_1247),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1434)
);

CKINVDCx6p67_ASAP7_75t_R g1435 ( 
.A(n_1347),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1271),
.B(n_1274),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1244),
.B(n_1314),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1416),
.B(n_1410),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1397),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1418),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1412),
.B(n_1405),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1389),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1391),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1417),
.Y(n_1445)
);

HB1xp67_ASAP7_75t_L g1446 ( 
.A(n_1384),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1394),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_L g1448 ( 
.A1(n_1432),
.A2(n_1363),
.B(n_1362),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1413),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1382),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_L g1451 ( 
.A1(n_1432),
.A2(n_1365),
.B(n_1431),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1370),
.Y(n_1452)
);

INVx2_ASAP7_75t_SL g1453 ( 
.A(n_1402),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1372),
.B(n_1368),
.Y(n_1454)
);

OAI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1364),
.A2(n_1365),
.B(n_1374),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1402),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1392),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1419),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1424),
.B(n_1425),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1388),
.B(n_1373),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1393),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1411),
.B(n_1426),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1411),
.B(n_1426),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1401),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1404),
.A2(n_1379),
.B(n_1422),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_L g1466 ( 
.A(n_1427),
.B(n_1428),
.Y(n_1466)
);

BUFx2_ASAP7_75t_L g1467 ( 
.A(n_1409),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1426),
.B(n_1433),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1409),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1433),
.Y(n_1470)
);

INVxp67_ASAP7_75t_L g1471 ( 
.A(n_1387),
.Y(n_1471)
);

BUFx2_ASAP7_75t_L g1472 ( 
.A(n_1409),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1396),
.B(n_1398),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1371),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1414),
.A2(n_1430),
.B(n_1381),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1406),
.B(n_1414),
.Y(n_1476)
);

NOR2x1_ASAP7_75t_L g1477 ( 
.A(n_1407),
.B(n_1376),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_SL g1478 ( 
.A(n_1367),
.B(n_1366),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1476),
.B(n_1438),
.Y(n_1479)
);

INVx3_ASAP7_75t_L g1480 ( 
.A(n_1445),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1461),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1476),
.B(n_1421),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1445),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1438),
.B(n_1460),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1420),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1438),
.B(n_1375),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1469),
.B(n_1375),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1464),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1469),
.B(n_1375),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1448),
.B(n_1399),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1441),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1469),
.B(n_1386),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1460),
.B(n_1415),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1447),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1456),
.B(n_1386),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1467),
.Y(n_1496)
);

NAND2x1p5_ASAP7_75t_L g1497 ( 
.A(n_1451),
.B(n_1423),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1439),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1458),
.B(n_1408),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1458),
.B(n_1408),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1449),
.B(n_1369),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1446),
.B(n_1380),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1447),
.B(n_1436),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_L g1505 ( 
.A(n_1448),
.B(n_1429),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1443),
.B(n_1434),
.Y(n_1506)
);

OAI21xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1479),
.A2(n_1451),
.B(n_1475),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_SL g1508 ( 
.A(n_1504),
.B(n_1455),
.Y(n_1508)
);

AOI221xp5_ASAP7_75t_L g1509 ( 
.A1(n_1490),
.A2(n_1455),
.B1(n_1475),
.B2(n_1465),
.C(n_1403),
.Y(n_1509)
);

AOI221xp5_ASAP7_75t_L g1510 ( 
.A1(n_1490),
.A2(n_1505),
.B1(n_1479),
.B2(n_1486),
.C(n_1506),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1481),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1481),
.Y(n_1512)
);

NOR4xp25_ASAP7_75t_SL g1513 ( 
.A(n_1483),
.B(n_1472),
.C(n_1474),
.D(n_1443),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1502),
.A2(n_1400),
.B1(n_1390),
.B2(n_1442),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1502),
.B(n_1459),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1498),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1479),
.B(n_1472),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1496),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1484),
.B(n_1493),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1502),
.A2(n_1442),
.B1(n_1385),
.B2(n_1395),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1498),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1494),
.B(n_1459),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1491),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1492),
.A2(n_1468),
.B(n_1470),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1496),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1488),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1505),
.A2(n_1378),
.B1(n_1385),
.B2(n_1442),
.Y(n_1527)
);

NAND4xp25_ASAP7_75t_L g1528 ( 
.A(n_1499),
.B(n_1463),
.C(n_1462),
.D(n_1471),
.Y(n_1528)
);

OAI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1503),
.A2(n_1457),
.B1(n_1477),
.B2(n_1454),
.C(n_1450),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1453),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1506),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1501),
.Y(n_1533)
);

OAI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1503),
.A2(n_1494),
.B1(n_1457),
.B2(n_1477),
.C(n_1454),
.Y(n_1534)
);

NAND4xp25_ASAP7_75t_L g1535 ( 
.A(n_1499),
.B(n_1462),
.C(n_1463),
.D(n_1468),
.Y(n_1535)
);

NAND4xp25_ASAP7_75t_L g1536 ( 
.A(n_1499),
.B(n_1462),
.C(n_1463),
.D(n_1468),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1486),
.A2(n_1444),
.B1(n_1450),
.B2(n_1466),
.C(n_1383),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1493),
.B(n_1474),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1500),
.A2(n_1473),
.B1(n_1440),
.B2(n_1478),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1523),
.A2(n_1492),
.B(n_1489),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1524),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1511),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1524),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1524),
.B(n_1486),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1512),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1524),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1518),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1507),
.B(n_1480),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1517),
.B(n_1492),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1507),
.Y(n_1551)
);

INVx4_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1516),
.Y(n_1553)
);

NOR3xp33_ASAP7_75t_SL g1554 ( 
.A(n_1509),
.B(n_1452),
.C(n_1435),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1515),
.B(n_1535),
.Y(n_1555)
);

OA21x2_ASAP7_75t_L g1556 ( 
.A1(n_1531),
.A2(n_1487),
.B(n_1489),
.Y(n_1556)
);

AND2x6_ASAP7_75t_SL g1557 ( 
.A(n_1522),
.B(n_1435),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_SL g1558 ( 
.A(n_1508),
.B(n_1497),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1517),
.B(n_1487),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1508),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1536),
.B(n_1488),
.Y(n_1561)
);

INVxp67_ASAP7_75t_SL g1562 ( 
.A(n_1521),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1518),
.Y(n_1563)
);

OA21x2_ASAP7_75t_L g1564 ( 
.A1(n_1526),
.A2(n_1489),
.B(n_1495),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1551),
.A2(n_1528),
.B1(n_1527),
.B2(n_1510),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1547),
.Y(n_1566)
);

INVx4_ASAP7_75t_L g1567 ( 
.A(n_1557),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1551),
.B(n_1519),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1561),
.B(n_1519),
.Y(n_1569)
);

NAND2x1_ASAP7_75t_L g1570 ( 
.A(n_1551),
.B(n_1525),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1547),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1555),
.B(n_1532),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1555),
.B(n_1532),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1555),
.B(n_1537),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1551),
.B(n_1533),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1561),
.B(n_1560),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1561),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1541),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1541),
.Y(n_1580)
);

NAND2xp33_ASAP7_75t_L g1581 ( 
.A(n_1554),
.B(n_1538),
.Y(n_1581)
);

NAND2x1p5_ASAP7_75t_L g1582 ( 
.A(n_1558),
.B(n_1423),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1560),
.B(n_1513),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1547),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1560),
.B(n_1539),
.Y(n_1585)
);

CKINVDCx16_ASAP7_75t_R g1586 ( 
.A(n_1560),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1547),
.A2(n_1514),
.B1(n_1520),
.B2(n_1529),
.Y(n_1587)
);

INVx1_ASAP7_75t_SL g1588 ( 
.A(n_1557),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1541),
.Y(n_1589)
);

AOI211xp5_ASAP7_75t_L g1590 ( 
.A1(n_1558),
.A2(n_1549),
.B(n_1545),
.C(n_1544),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1543),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1543),
.Y(n_1592)
);

INVx4_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1543),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1543),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1563),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1546),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1546),
.Y(n_1598)
);

AND2x4_ASAP7_75t_SL g1599 ( 
.A(n_1554),
.B(n_1548),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1553),
.B(n_1482),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1546),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1553),
.B(n_1485),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1547),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1547),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1550),
.B(n_1530),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1594),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1550),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1568),
.B(n_1553),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1578),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1574),
.A2(n_1547),
.B1(n_1544),
.B2(n_1542),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1578),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1565),
.B(n_1554),
.C(n_1558),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1586),
.A2(n_1547),
.B1(n_1542),
.B2(n_1544),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1586),
.B(n_1562),
.Y(n_1616)
);

AOI222xp33_ASAP7_75t_L g1617 ( 
.A1(n_1587),
.A2(n_1544),
.B1(n_1542),
.B2(n_1545),
.C1(n_1547),
.C2(n_1534),
.Y(n_1617)
);

NAND2xp33_ASAP7_75t_R g1618 ( 
.A(n_1583),
.B(n_1564),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1571),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1562),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1576),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1623)
);

INVx1_ASAP7_75t_SL g1624 ( 
.A(n_1588),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1572),
.B(n_1573),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1599),
.B(n_1550),
.Y(n_1626)
);

OAI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1585),
.A2(n_1542),
.B1(n_1544),
.B2(n_1556),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_1570),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1567),
.B(n_1559),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1569),
.B(n_1562),
.Y(n_1630)
);

NAND2x1p5_ASAP7_75t_L g1631 ( 
.A(n_1567),
.B(n_1423),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1569),
.B(n_1564),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1567),
.B(n_1370),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1581),
.A2(n_1544),
.B(n_1542),
.Y(n_1634)
);

AOI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1583),
.A2(n_1542),
.B1(n_1545),
.B2(n_1540),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1571),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1579),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1575),
.B(n_1564),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1579),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1590),
.A2(n_1549),
.B(n_1545),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1570),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1611),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1629),
.B(n_1567),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1633),
.B(n_1593),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1621),
.B(n_1606),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1629),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1616),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1628),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1624),
.B(n_1593),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1625),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

AO21x2_ASAP7_75t_L g1653 ( 
.A1(n_1627),
.A2(n_1605),
.B(n_1584),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1613),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1614),
.A2(n_1593),
.B1(n_1590),
.B2(n_1549),
.Y(n_1655)
);

INVx2_ASAP7_75t_SL g1656 ( 
.A(n_1628),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1628),
.Y(n_1657)
);

AOI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1618),
.A2(n_1545),
.B1(n_1593),
.B2(n_1540),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1630),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1617),
.A2(n_1556),
.B1(n_1540),
.B2(n_1564),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1609),
.B(n_1606),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1613),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1559),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1639),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1607),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1640),
.B(n_1596),
.Y(n_1667)
);

OAI321xp33_ASAP7_75t_L g1668 ( 
.A1(n_1658),
.A2(n_1612),
.A3(n_1635),
.B1(n_1615),
.B2(n_1634),
.C(n_1638),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1651),
.B(n_1607),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_SL g1670 ( 
.A1(n_1655),
.A2(n_1659),
.B(n_1660),
.C(n_1643),
.Y(n_1670)
);

OAI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1643),
.A2(n_1632),
.B1(n_1638),
.B2(n_1582),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1653),
.A2(n_1650),
.B1(n_1644),
.B2(n_1647),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1647),
.B(n_1620),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1650),
.B(n_1559),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_SL g1675 ( 
.A1(n_1653),
.A2(n_1632),
.B1(n_1622),
.B2(n_1626),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1642),
.Y(n_1676)
);

AOI21xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1650),
.A2(n_1653),
.B(n_1631),
.Y(n_1677)
);

AOI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1648),
.A2(n_1584),
.B1(n_1605),
.B2(n_1636),
.C(n_1608),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1644),
.B(n_1559),
.Y(n_1679)
);

AOI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1667),
.A2(n_1623),
.B1(n_1626),
.B2(n_1622),
.Y(n_1680)
);

O2A1O1Ixp33_ASAP7_75t_L g1681 ( 
.A1(n_1657),
.A2(n_1641),
.B(n_1631),
.C(n_1582),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1642),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1652),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1654),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1662),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1646),
.B(n_1559),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1674),
.B(n_1661),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1673),
.B(n_1663),
.Y(n_1688)
);

OAI321xp33_ASAP7_75t_L g1689 ( 
.A1(n_1670),
.A2(n_1667),
.A3(n_1649),
.B1(n_1656),
.B2(n_1666),
.C(n_1645),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1680),
.B(n_1672),
.Y(n_1690)
);

OAI31xp33_ASAP7_75t_SL g1691 ( 
.A1(n_1675),
.A2(n_1666),
.A3(n_1623),
.B(n_1665),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1679),
.B(n_1649),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1669),
.B(n_1664),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1678),
.A2(n_1665),
.B1(n_1664),
.B2(n_1584),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1683),
.B(n_1656),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1693),
.B(n_1690),
.Y(n_1697)
);

OAI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1691),
.A2(n_1677),
.B(n_1681),
.C(n_1678),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1692),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1694),
.A2(n_1695),
.B1(n_1686),
.B2(n_1688),
.Y(n_1700)
);

NOR3xp33_ASAP7_75t_SL g1701 ( 
.A(n_1689),
.B(n_1668),
.C(n_1684),
.Y(n_1701)
);

NAND5xp2_ASAP7_75t_L g1702 ( 
.A(n_1695),
.B(n_1631),
.C(n_1682),
.D(n_1685),
.E(n_1582),
.Y(n_1702)
);

NOR2xp33_ASAP7_75t_L g1703 ( 
.A(n_1694),
.B(n_1557),
.Y(n_1703)
);

AOI221xp5_ASAP7_75t_L g1704 ( 
.A1(n_1692),
.A2(n_1671),
.B1(n_1605),
.B2(n_1604),
.C(n_1566),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_SL g1705 ( 
.A(n_1696),
.B(n_1596),
.Y(n_1705)
);

OAI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1698),
.A2(n_1687),
.B(n_1619),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1563),
.Y(n_1707)
);

AO21x1_ASAP7_75t_L g1708 ( 
.A1(n_1700),
.A2(n_1636),
.B(n_1619),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1699),
.B(n_1600),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1701),
.A2(n_1703),
.B(n_1704),
.C(n_1702),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1707),
.B(n_1705),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1710),
.B(n_1608),
.C(n_1604),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1706),
.A2(n_1566),
.B(n_1602),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1709),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1708),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1706),
.B(n_1603),
.Y(n_1716)
);

AOI22xp33_ASAP7_75t_L g1717 ( 
.A1(n_1715),
.A2(n_1556),
.B1(n_1540),
.B2(n_1564),
.Y(n_1717)
);

INVx1_ASAP7_75t_SL g1718 ( 
.A(n_1714),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1711),
.Y(n_1719)
);

XOR2xp5_ASAP7_75t_L g1720 ( 
.A(n_1716),
.B(n_1377),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1712),
.Y(n_1721)
);

NOR3xp33_ASAP7_75t_L g1722 ( 
.A(n_1718),
.B(n_1713),
.C(n_1377),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1719),
.B(n_1580),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1720),
.A2(n_1552),
.B(n_1548),
.C(n_1549),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1723),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1720),
.B1(n_1721),
.B2(n_1722),
.Y(n_1726)
);

AO21x1_ASAP7_75t_L g1727 ( 
.A1(n_1726),
.A2(n_1724),
.B(n_1589),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1726),
.A2(n_1717),
.B1(n_1556),
.B2(n_1540),
.Y(n_1728)
);

NAND2xp33_ASAP7_75t_R g1729 ( 
.A(n_1727),
.B(n_1540),
.Y(n_1729)
);

NAND3xp33_ASAP7_75t_L g1730 ( 
.A(n_1728),
.B(n_1602),
.C(n_1601),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1729),
.Y(n_1731)
);

OAI22xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1730),
.A2(n_1540),
.B1(n_1556),
.B2(n_1564),
.Y(n_1732)
);

AOI22xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1731),
.A2(n_1592),
.B1(n_1598),
.B2(n_1597),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_SL g1734 ( 
.A(n_1733),
.B(n_1732),
.C(n_1601),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1734),
.B(n_1580),
.Y(n_1735)
);

AOI21xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1598),
.B(n_1597),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1736),
.A2(n_1595),
.B1(n_1592),
.B2(n_1591),
.C(n_1589),
.Y(n_1737)
);

AOI211xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1595),
.B(n_1591),
.C(n_1563),
.Y(n_1738)
);


endmodule