module fake_jpeg_9077_n_59 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_59);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_1),
.B(n_2),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_17),
.A2(n_6),
.B(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_7),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_35),
.A2(n_11),
.B1(n_12),
.B2(n_8),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_40),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_8),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_36),
.B1(n_32),
.B2(n_28),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_25),
.A2(n_30),
.B1(n_27),
.B2(n_20),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_22),
.B(n_21),
.C(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_26),
.A2(n_20),
.B1(n_23),
.B2(n_29),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_23),
.A2(n_29),
.B1(n_33),
.B2(n_18),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_49),
.A2(n_38),
.B1(n_45),
.B2(n_46),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_50),
.B(n_51),
.Y(n_52)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_53),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_44),
.C(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_44),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_54),
.C(n_47),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_56),
.B1(n_42),
.B2(n_48),
.Y(n_58)
);

AOI211xp5_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_33),
.B(n_45),
.C(n_19),
.Y(n_59)
);


endmodule