module fake_jpeg_9252_n_61 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_61);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_61;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_8),
.B(n_1),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_21),
.B(n_16),
.C(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_11),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_1),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_25),
.A2(n_13),
.B1(n_14),
.B2(n_8),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g26 ( 
.A(n_20),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_22),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_25),
.A2(n_21),
.B1(n_19),
.B2(n_15),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_32),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_24),
.B(n_26),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_34),
.B(n_17),
.Y(n_42)
);

AOI22x1_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_11),
.B1(n_2),
.B2(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_36),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_34),
.B1(n_17),
.B2(n_35),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_48),
.C(n_50),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_38),
.B1(n_28),
.B2(n_3),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_40),
.C(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_43),
.C(n_44),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_54),
.B(n_45),
.Y(n_56)
);

AO21x1_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_57),
.B(n_28),
.Y(n_58)
);

A2O1A1O1Ixp25_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_42),
.B(n_44),
.C(n_41),
.D(n_50),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_2),
.Y(n_59)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_38),
.C(n_28),
.Y(n_60)
);

BUFx24_ASAP7_75t_SL g61 ( 
.A(n_60),
.Y(n_61)
);


endmodule