module fake_jpeg_283_n_73 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_73);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_73;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx5_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_7),
.B(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_3),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_4),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_19),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_26),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_16),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_24),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_38),
.C(n_18),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_15),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_9),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_22),
.B1(n_28),
.B2(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_46),
.Y(n_53)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_50),
.B(n_33),
.C(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_55),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_39),
.C(n_31),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_43),
.C(n_49),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_20),
.B(n_25),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_54),
.A2(n_56),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_18),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_21),
.B(n_13),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_61),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_53),
.A2(n_47),
.B1(n_46),
.B2(n_44),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_21),
.B(n_43),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_58),
.B(n_61),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_64),
.B(n_12),
.Y(n_68)
);

BUFx24_ASAP7_75t_SL g65 ( 
.A(n_57),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_5),
.C(n_6),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_68),
.B(n_13),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_13),
.C(n_1),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_69),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_1),
.C(n_2),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_71),
.Y(n_73)
);


endmodule