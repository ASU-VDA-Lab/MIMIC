module fake_jpeg_2846_n_630 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_630);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_630;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_568;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_11),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_13),
.B(n_2),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_59),
.Y(n_139)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_60),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_61),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_62),
.B(n_66),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_63),
.Y(n_179)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_65),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_27),
.B(n_18),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_67),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_71),
.Y(n_149)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_69),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_70),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_27),
.B(n_19),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_72),
.Y(n_138)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_74),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_19),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_76),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_21),
.B(n_18),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_77),
.Y(n_143)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_35),
.Y(n_78)
);

INVx5_ASAP7_75t_SL g222 ( 
.A(n_78),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_79),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx8_ASAP7_75t_L g216 ( 
.A(n_80),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_83),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_34),
.B(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_88),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_42),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_85),
.B(n_91),
.Y(n_160)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_17),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_92),
.Y(n_195)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_93),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_45),
.B(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_126),
.Y(n_167)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_31),
.Y(n_97)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_98),
.B(n_99),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_38),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_100),
.Y(n_185)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_101),
.Y(n_157)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_105),
.Y(n_223)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_35),
.Y(n_106)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_38),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_113),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_39),
.Y(n_109)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_41),
.Y(n_111)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_111),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_41),
.Y(n_112)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_112),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_38),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_35),
.Y(n_114)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_114),
.Y(n_214)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_125),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_120),
.Y(n_224)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_37),
.Y(n_121)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_121),
.Y(n_226)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_37),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_122),
.B(n_123),
.Y(n_203)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_37),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_48),
.Y(n_124)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_50),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_48),
.B(n_1),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_24),
.A2(n_1),
.B(n_3),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_127),
.B(n_105),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_52),
.Y(n_129)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_52),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_129),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_66),
.A2(n_52),
.B1(n_56),
.B2(n_24),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_71),
.A2(n_46),
.B1(n_56),
.B2(n_40),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_74),
.B1(n_94),
.B2(n_92),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_64),
.A2(n_57),
.B1(n_53),
.B2(n_25),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_128),
.A2(n_23),
.B1(n_28),
.B2(n_51),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_140),
.A2(n_176),
.B1(n_192),
.B2(n_198),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_82),
.A2(n_57),
.B1(n_53),
.B2(n_25),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_142),
.A2(n_144),
.B1(n_148),
.B2(n_171),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_95),
.A2(n_40),
.B1(n_51),
.B2(n_46),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_83),
.A2(n_54),
.B1(n_28),
.B2(n_23),
.Y(n_147)
);

OA22x2_ASAP7_75t_L g260 ( 
.A1(n_147),
.A2(n_150),
.B1(n_151),
.B2(n_155),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_58),
.A2(n_37),
.B1(n_28),
.B2(n_23),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_86),
.A2(n_43),
.B1(n_3),
.B2(n_5),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_43),
.B1(n_3),
.B2(n_5),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_102),
.A2(n_43),
.B1(n_5),
.B2(n_7),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g282 ( 
.A(n_170),
.B(n_182),
.C(n_195),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_59),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_171)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_60),
.Y(n_175)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_63),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_70),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_181),
.A2(n_197),
.B1(n_202),
.B2(n_210),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_106),
.B(n_10),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_184),
.B(n_204),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_114),
.B(n_10),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_186),
.B(n_190),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_12),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_79),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_81),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_104),
.A2(n_16),
.B1(n_112),
.B2(n_111),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_65),
.Y(n_199)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_199),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_110),
.A2(n_16),
.B1(n_116),
.B2(n_109),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_122),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_121),
.Y(n_205)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_205),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_107),
.B(n_16),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_206),
.B(n_157),
.Y(n_248)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_69),
.Y(n_207)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_207),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_67),
.B(n_72),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_208),
.B(n_223),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_77),
.A2(n_97),
.B1(n_115),
.B2(n_103),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_123),
.A2(n_80),
.B1(n_78),
.B2(n_87),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_213),
.A2(n_225),
.B1(n_223),
.B2(n_182),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_L g297 ( 
.A1(n_215),
.A2(n_154),
.B(n_193),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_78),
.A2(n_90),
.B1(n_93),
.B2(n_119),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_218),
.A2(n_61),
.B1(n_225),
.B2(n_202),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_80),
.A2(n_44),
.B1(n_86),
.B2(n_23),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_216),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_228),
.B(n_229),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_231),
.A2(n_299),
.B1(n_307),
.B2(n_309),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_149),
.B(n_61),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_232),
.B(n_233),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_173),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_235),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_172),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_236),
.Y(n_330)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_238),
.Y(n_357)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_161),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_152),
.Y(n_241)
);

O2A1O1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_215),
.A2(n_140),
.B(n_151),
.C(n_176),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_242),
.A2(n_266),
.B(n_284),
.Y(n_341)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_156),
.B(n_169),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_243),
.Y(n_314)
);

OAI21xp33_ASAP7_75t_SL g329 ( 
.A1(n_245),
.A2(n_279),
.B(n_306),
.Y(n_329)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_145),
.A2(n_131),
.B(n_167),
.Y(n_246)
);

NOR3xp33_ASAP7_75t_SL g334 ( 
.A(n_246),
.B(n_257),
.C(n_281),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_158),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_247),
.B(n_270),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_248),
.B(n_250),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_194),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_251),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_172),
.Y(n_250)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_166),
.Y(n_252)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_164),
.B(n_203),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_253),
.B(n_276),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_139),
.Y(n_254)
);

INVx13_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_255),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_162),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_256),
.B(n_259),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_165),
.B(n_134),
.C(n_146),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_289),
.C(n_294),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_188),
.Y(n_259)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_189),
.Y(n_261)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_179),
.Y(n_263)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_264),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_265),
.B(n_267),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_L g266 ( 
.A1(n_151),
.A2(n_222),
.B(n_192),
.C(n_168),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_160),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_152),
.B(n_220),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_269),
.B(n_271),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_185),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_220),
.B(n_221),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g272 ( 
.A(n_216),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_272),
.B(n_277),
.Y(n_343)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_273),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_181),
.A2(n_191),
.B1(n_212),
.B2(n_209),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_275),
.B1(n_298),
.B2(n_231),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_174),
.A2(n_178),
.B1(n_195),
.B2(n_201),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_159),
.B(n_221),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_143),
.B(n_159),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_143),
.A2(n_138),
.B1(n_177),
.B2(n_141),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_187),
.B(n_138),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_280),
.B(n_301),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_282),
.B(n_288),
.Y(n_346)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_141),
.Y(n_283)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

NAND2x1_ASAP7_75t_SL g284 ( 
.A(n_196),
.B(n_217),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_179),
.Y(n_285)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_163),
.Y(n_286)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_286),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_177),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_163),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_219),
.B(n_196),
.C(n_193),
.Y(n_289)
);

BUFx12_ASAP7_75t_L g290 ( 
.A(n_154),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_290),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_178),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_291),
.Y(n_320)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_201),
.Y(n_292)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_292),
.Y(n_354)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_211),
.Y(n_293)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_183),
.B(n_211),
.Y(n_294)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_183),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_296),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_297),
.A2(n_284),
.B(n_294),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_154),
.A2(n_215),
.B1(n_135),
.B2(n_202),
.Y(n_298)
);

BUFx12f_ASAP7_75t_L g299 ( 
.A(n_180),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_180),
.B(n_157),
.C(n_153),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_253),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_200),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_200),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_303),
.B(n_250),
.Y(n_348)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_304),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_136),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_305),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g306 ( 
.A1(n_213),
.A2(n_28),
.B1(n_23),
.B2(n_148),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_207),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_200),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_237),
.A2(n_308),
.B1(n_262),
.B2(n_302),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_311),
.A2(n_324),
.B1(n_328),
.B2(n_238),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_244),
.B(n_247),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_313),
.B(n_355),
.Y(n_392)
);

AOI32xp33_ASAP7_75t_L g327 ( 
.A1(n_297),
.A2(n_242),
.A3(n_298),
.B1(n_260),
.B2(n_230),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_327),
.B(n_346),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_237),
.A2(n_266),
.B1(n_260),
.B2(n_274),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_241),
.C(n_236),
.Y(n_368)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_351),
.C(n_345),
.Y(n_362)
);

A2O1A1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_253),
.A2(n_300),
.B(n_270),
.C(n_260),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_335),
.B(n_353),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_276),
.A2(n_275),
.B1(n_240),
.B2(n_283),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_348),
.Y(n_405)
);

NOR3xp33_ASAP7_75t_SL g351 ( 
.A(n_260),
.B(n_258),
.C(n_278),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_294),
.A2(n_243),
.B1(n_289),
.B2(n_292),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_353),
.A2(n_272),
.B1(n_290),
.B2(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_243),
.B(n_304),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_261),
.B(n_268),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_352),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_372),
.Y(n_416)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_356),
.Y(n_363)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_313),
.B(n_295),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_365),
.B(n_374),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_276),
.C(n_264),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_366),
.B(n_368),
.C(n_377),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_325),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_367),
.B(n_369),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_355),
.Y(n_370)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_324),
.A2(n_293),
.B1(n_286),
.B2(n_296),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_371),
.A2(n_384),
.B1(n_398),
.B2(n_329),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_347),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_341),
.A2(n_255),
.B(n_239),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_373),
.A2(n_348),
.B(n_330),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_316),
.B(n_273),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_349),
.Y(n_375)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_375),
.Y(n_433)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_376),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_252),
.C(n_287),
.Y(n_377)
);

AND2x2_ASAP7_75t_SL g378 ( 
.A(n_358),
.B(n_227),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_378),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_350),
.B(n_309),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_379),
.B(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_380),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_315),
.B(n_263),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_382),
.A2(n_340),
.B1(n_320),
.B2(n_344),
.Y(n_413)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_311),
.A2(n_305),
.B1(n_234),
.B2(n_235),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_322),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_386),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_338),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_387),
.A2(n_395),
.B(n_402),
.Y(n_426)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_357),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_390),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_341),
.A2(n_254),
.B1(n_285),
.B2(n_299),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_394),
.B1(n_323),
.B2(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_359),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_359),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_393),
.Y(n_422)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_318),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_328),
.A2(n_299),
.B1(n_272),
.B2(n_227),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g395 ( 
.A(n_334),
.B(n_335),
.CI(n_361),
.CON(n_395),
.SN(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_397),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_343),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_350),
.B(n_290),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_400),
.Y(n_434)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

OA21x2_ASAP7_75t_L g401 ( 
.A1(n_327),
.A2(n_351),
.B(n_358),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_401),
.B(n_403),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_340),
.A2(n_314),
.B1(n_358),
.B2(n_310),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_350),
.B(n_310),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_404),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_406),
.Y(n_412)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_407),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_333),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_410),
.B(n_424),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_413),
.A2(n_370),
.B1(n_405),
.B2(n_398),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_401),
.A2(n_373),
.B(n_405),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_415),
.A2(n_425),
.B(n_442),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_382),
.A2(n_394),
.B1(n_363),
.B2(n_392),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_419),
.A2(n_436),
.B1(n_444),
.B2(n_445),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_420),
.B(n_428),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_406),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_421),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_392),
.B(n_339),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_384),
.A2(n_320),
.B1(n_344),
.B2(n_360),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_369),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_372),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_339),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g467 ( 
.A(n_439),
.B(n_378),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_366),
.B(n_331),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_443),
.C(n_378),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_401),
.A2(n_317),
.B(n_330),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_377),
.B(n_317),
.C(n_312),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_371),
.A2(n_342),
.B1(n_319),
.B2(n_357),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_401),
.A2(n_319),
.B1(n_342),
.B2(n_321),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_448),
.A2(n_473),
.B1(n_430),
.B2(n_429),
.Y(n_490)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_422),
.Y(n_449)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_449),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_435),
.B(n_368),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_450),
.B(n_458),
.C(n_471),
.Y(n_489)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_422),
.Y(n_451)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_451),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_432),
.A2(n_405),
.B1(n_364),
.B2(n_397),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_453),
.A2(n_460),
.B(n_462),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g456 ( 
.A(n_418),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_456),
.B(n_459),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_427),
.B(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_457),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_431),
.B(n_367),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_442),
.A2(n_364),
.B(n_395),
.Y(n_460)
);

XNOR2x2_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_395),
.Y(n_462)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_407),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_465),
.B(n_466),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_412),
.B(n_421),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_467),
.B(n_447),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_437),
.A2(n_379),
.B(n_399),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_468),
.A2(n_452),
.B(n_460),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_411),
.B(n_385),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_470),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_431),
.B(n_312),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_435),
.B(n_375),
.C(n_391),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_438),
.B(n_404),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_474),
.Y(n_487)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_423),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_412),
.B(n_400),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_433),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_475),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_417),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_477),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_396),
.Y(n_477)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_482),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_411),
.B(n_337),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_480),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_441),
.B(n_380),
.C(n_390),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_483),
.C(n_415),
.Y(n_491)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_423),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_383),
.C(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_490),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_491),
.B(n_453),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_493),
.A2(n_452),
.B(n_468),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_426),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_504),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_483),
.C(n_458),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_506),
.C(n_507),
.Y(n_525)
);

XOR2x2_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_426),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_476),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_455),
.A2(n_424),
.B1(n_429),
.B2(n_445),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_501),
.B(n_508),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_478),
.B(n_428),
.Y(n_503)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_503),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_461),
.B(n_420),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_439),
.C(n_432),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_461),
.B(n_434),
.C(n_425),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_455),
.A2(n_436),
.B1(n_419),
.B2(n_413),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_455),
.A2(n_410),
.B1(n_434),
.B2(n_414),
.Y(n_509)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_472),
.Y(n_510)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

O2A1O1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_466),
.A2(n_417),
.B(n_446),
.C(n_447),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_474),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_469),
.A2(n_416),
.B1(n_414),
.B2(n_409),
.Y(n_512)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_513),
.B(n_454),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_462),
.B(n_440),
.C(n_337),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_515),
.C(n_448),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_440),
.C(n_409),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_526),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_505),
.B(n_482),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_520),
.B(n_522),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_511),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_523),
.A2(n_493),
.B(n_516),
.Y(n_546)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_529),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_489),
.B(n_449),
.C(n_451),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_537),
.C(n_507),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_465),
.Y(n_531)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_531),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_532),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_491),
.B(n_457),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_533),
.B(n_534),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_489),
.B(n_463),
.Y(n_534)
);

NOR3xp33_ASAP7_75t_SL g563 ( 
.A(n_535),
.B(n_488),
.C(n_500),
.Y(n_563)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_517),
.Y(n_536)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_536),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_495),
.B(n_494),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_492),
.B(n_477),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_545),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_486),
.B(n_388),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_541),
.B(n_542),
.Y(n_562)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_500),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_499),
.B(n_497),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_543),
.A2(n_544),
.B1(n_497),
.B2(n_488),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_498),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g569 ( 
.A1(n_546),
.A2(n_558),
.B(n_529),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g571 ( 
.A(n_547),
.B(n_525),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_515),
.C(n_514),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_550),
.B(n_557),
.Y(n_576)
);

INVx13_ASAP7_75t_L g551 ( 
.A(n_536),
.Y(n_551)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_551),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_518),
.B(n_509),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_517),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_555),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_539),
.B(n_492),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_556),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_537),
.B(n_506),
.C(n_504),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_SL g558 ( 
.A1(n_523),
.A2(n_516),
.B(n_498),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_561),
.A2(n_563),
.B1(n_540),
.B2(n_518),
.Y(n_578)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_530),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_526),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_525),
.B(n_513),
.C(n_485),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_567),
.B(n_557),
.C(n_547),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_564),
.B(n_533),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_568),
.B(n_571),
.Y(n_593)
);

OR2x2_ASAP7_75t_L g597 ( 
.A(n_569),
.B(n_578),
.Y(n_597)
);

XOR2xp5_ASAP7_75t_L g570 ( 
.A(n_560),
.B(n_524),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_570),
.B(n_572),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_558),
.A2(n_539),
.B(n_527),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_575),
.A2(n_579),
.B(n_554),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_553),
.A2(n_527),
.B1(n_528),
.B2(n_508),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_580),
.A2(n_581),
.B1(n_585),
.B2(n_552),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_548),
.A2(n_549),
.B1(n_521),
.B2(n_562),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_565),
.B(n_524),
.C(n_519),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_583),
.B(n_567),
.C(n_560),
.Y(n_590)
);

MAJx2_ASAP7_75t_L g584 ( 
.A(n_550),
.B(n_496),
.C(n_545),
.Y(n_584)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_554),
.Y(n_598)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_553),
.A2(n_528),
.B1(n_501),
.B2(n_454),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_574),
.A2(n_549),
.B1(n_552),
.B2(n_559),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_586),
.B(n_588),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_587),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_576),
.B(n_571),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_572),
.B(n_565),
.Y(n_589)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_589),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_590),
.B(n_592),
.Y(n_611)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_591),
.B(n_594),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_570),
.B(n_583),
.C(n_575),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_559),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_SL g605 ( 
.A1(n_595),
.A2(n_487),
.B(n_556),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_598),
.B(n_599),
.C(n_600),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_569),
.B(n_546),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_580),
.B(n_566),
.Y(n_600)
);

A2O1A1Ixp33_ASAP7_75t_L g602 ( 
.A1(n_599),
.A2(n_484),
.B(n_577),
.C(n_555),
.Y(n_602)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_602),
.A2(n_606),
.B(n_596),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g613 ( 
.A(n_605),
.B(n_502),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_600),
.A2(n_577),
.B(n_563),
.Y(n_606)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_597),
.A2(n_585),
.B1(n_484),
.B2(n_566),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_607),
.B(n_592),
.Y(n_614)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_597),
.A2(n_487),
.B(n_538),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_608),
.A2(n_598),
.B(n_593),
.Y(n_612)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_612),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_613),
.B(n_614),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_609),
.B(n_611),
.C(n_604),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_615),
.B(n_616),
.Y(n_621)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_610),
.B(n_596),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_617),
.B(n_618),
.C(n_610),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_603),
.B(n_590),
.Y(n_618)
);

MAJx2_ASAP7_75t_L g625 ( 
.A(n_619),
.B(n_584),
.C(n_464),
.Y(n_625)
);

AO221x1_ASAP7_75t_L g622 ( 
.A1(n_613),
.A2(n_601),
.B1(n_606),
.B2(n_608),
.C(n_551),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_622),
.A2(n_602),
.B(n_607),
.Y(n_624)
);

OAI21xp5_ASAP7_75t_L g626 ( 
.A1(n_624),
.A2(n_625),
.B(n_620),
.Y(n_626)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_626),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g627 ( 
.A1(n_624),
.A2(n_623),
.B1(n_621),
.B2(n_475),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_628),
.B(n_627),
.Y(n_629)
);

XNOR2xp5_ASAP7_75t_L g630 ( 
.A(n_629),
.B(n_479),
.Y(n_630)
);


endmodule