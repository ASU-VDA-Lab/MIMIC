module real_jpeg_15612_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_202;
wire n_128;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_324;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx1_ASAP7_75t_L g151 ( 
.A(n_0),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_0),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_0),
.Y(n_165)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_2),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_2),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_2),
.A2(n_113),
.B1(n_175),
.B2(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_2),
.A2(n_113),
.B1(n_447),
.B2(n_449),
.Y(n_446)
);

AOI22xp33_ASAP7_75t_SL g457 ( 
.A1(n_2),
.A2(n_113),
.B1(n_458),
.B2(n_460),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_3),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_137),
.B1(n_178),
.B2(n_235),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_3),
.A2(n_178),
.B1(n_203),
.B2(n_347),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_3),
.A2(n_178),
.B1(n_385),
.B2(n_390),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_4),
.A2(n_216),
.B1(n_218),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_5),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g214 ( 
.A(n_5),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_6),
.Y(n_167)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_6),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g209 ( 
.A(n_6),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_7),
.A2(n_137),
.B1(n_141),
.B2(n_142),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_7),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_7),
.A2(n_141),
.B1(n_179),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_7),
.A2(n_141),
.B1(n_362),
.B2(n_365),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_7),
.A2(n_141),
.B1(n_434),
.B2(n_437),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_8),
.B(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_8),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_8),
.A2(n_273),
.B(n_340),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_8),
.A2(n_370),
.A3(n_373),
.B1(n_376),
.B2(n_381),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_8),
.B(n_261),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_8),
.A2(n_90),
.B1(n_474),
.B2(n_480),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_8),
.A2(n_336),
.B1(n_499),
.B2(n_503),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_9),
.A2(n_293),
.B1(n_294),
.B2(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_9),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_9),
.A2(n_296),
.B1(n_309),
.B2(n_314),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_9),
.A2(n_296),
.B1(n_425),
.B2(n_429),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_9),
.A2(n_296),
.B1(n_475),
.B2(n_477),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_10),
.A2(n_69),
.B1(n_73),
.B2(n_74),
.Y(n_68)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_10),
.A2(n_73),
.B1(n_240),
.B2(n_245),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_10),
.A2(n_73),
.B1(n_281),
.B2(n_285),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_78),
.B1(n_84),
.B2(n_89),
.Y(n_77)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_89),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_12),
.A2(n_95),
.B1(n_99),
.B2(n_103),
.Y(n_94)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_12),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_12),
.A2(n_103),
.B1(n_203),
.B2(n_205),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_13),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_13),
.Y(n_130)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_13),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_14),
.Y(n_155)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_15),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g330 ( 
.A(n_15),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_16),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_16),
.A2(n_61),
.B1(n_185),
.B2(n_189),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_16),
.A2(n_61),
.B1(n_324),
.B2(n_327),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_17),
.Y(n_112)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_17),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_17),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_299),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_297),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_250),
.Y(n_21)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_22),
.B(n_250),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_191),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_109),
.C(n_144),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_25),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_76),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g525 ( 
.A1(n_26),
.A2(n_27),
.B1(n_76),
.B2(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_55),
.B1(n_66),
.B2(n_68),
.Y(n_27)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_28),
.B(n_68),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_28),
.A2(n_66),
.B1(n_421),
.B2(n_424),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_28),
.A2(n_66),
.B1(n_424),
.B2(n_446),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_28),
.A2(n_66),
.B1(n_361),
.B2(n_446),
.Y(n_508)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_41),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_34),
.Y(n_439)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_35),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_35),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_36),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_38),
.Y(n_389)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B1(n_50),
.B2(n_52),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_44),
.Y(n_375)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_45),
.Y(n_409)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_49),
.Y(n_413)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_51),
.Y(n_405)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_53),
.Y(n_197)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_55),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g364 ( 
.A(n_60),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_60),
.Y(n_430)
);

INVx4_ASAP7_75t_L g448 ( 
.A(n_60),
.Y(n_448)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_64),
.Y(n_423)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_65),
.Y(n_350)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_65),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_66),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_67),
.A2(n_194),
.B1(n_195),
.B2(n_202),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_67),
.A2(n_194),
.B1(n_346),
.B2(n_351),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_67),
.A2(n_194),
.B1(n_346),
.B2(n_360),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_67),
.B(n_336),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_76),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_90),
.B1(n_94),
.B2(n_104),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_77),
.A2(n_90),
.B1(n_279),
.B2(n_287),
.Y(n_278)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_82),
.Y(n_436)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_83),
.Y(n_418)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_83),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_87),
.Y(n_217)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_88),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_90),
.A2(n_212),
.B(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_90),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_90),
.A2(n_433),
.B1(n_440),
.B2(n_441),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_90),
.A2(n_287),
.B1(n_457),
.B2(n_474),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_92),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_94),
.Y(n_228)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_98),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_102),
.Y(n_286)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_107),
.Y(n_483)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_108),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_109),
.B(n_144),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B1(n_136),
.B2(n_143),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_110),
.A2(n_115),
.B1(n_143),
.B2(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_111),
.Y(n_142)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_115),
.A2(n_136),
.B1(n_143),
.B2(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_115),
.A2(n_143),
.B1(n_292),
.B2(n_339),
.Y(n_338)
);

AO21x2_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_124),
.B(n_129),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_122),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_124),
.A2(n_264),
.B1(n_272),
.B2(n_274),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_125),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

AO22x2_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_132),
.Y(n_372)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_134),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2x1_ASAP7_75t_R g335 ( 
.A(n_143),
.B(n_336),
.Y(n_335)
);

OAI22x1_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_173),
.B1(n_183),
.B2(n_184),
.Y(n_144)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_145),
.A2(n_183),
.B1(n_184),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_145),
.A2(n_183),
.B1(n_308),
.B2(n_318),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_145),
.A2(n_183),
.B1(n_318),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_145),
.A2(n_183),
.B1(n_308),
.B2(n_498),
.Y(n_497)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_146),
.A2(n_174),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_156),
.B(n_162),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_153),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_153),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_155),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_155),
.Y(n_506)
);

INVxp33_ASAP7_75t_L g381 ( 
.A(n_156),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_161),
.Y(n_260)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_161),
.Y(n_317)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_161),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_166),
.B1(n_168),
.B2(n_170),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_167),
.Y(n_204)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_222),
.B1(n_248),
.B2(n_249),
.Y(n_191)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_210),
.B1(n_211),
.B2(n_221),
.Y(n_192)
);

INVxp33_ASAP7_75t_SL g221 ( 
.A(n_193),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVxp67_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_201),
.Y(n_366)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_201),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_212),
.Y(n_230)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_214),
.Y(n_289)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_214),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_232),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_225),
.B(n_227),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_225),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_254),
.Y(n_253)
);

AOI22x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_229),
.A2(n_280),
.B1(n_323),
.B2(n_331),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_229),
.A2(n_323),
.B1(n_384),
.B2(n_392),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_229),
.A2(n_456),
.B1(n_463),
.B2(n_464),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx6_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_244),
.Y(n_313)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.C(n_255),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_251),
.B(n_253),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_255),
.B(n_520),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.C(n_290),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_256),
.A2(n_290),
.B1(n_291),
.B2(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_256),
.Y(n_524)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_257),
.Y(n_353)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2x1_ASAP7_75t_L g522 ( 
.A(n_262),
.B(n_523),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_278),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_278),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_518),
.B(n_532),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_395),
.B(n_517),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_354),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_303),
.B(n_354),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_337),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_305),
.B(n_306),
.C(n_337),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_321),
.C(n_335),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_307),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_321),
.A2(n_322),
.B1(n_335),
.B2(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_330),
.Y(n_459)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_330),
.Y(n_462)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_330),
.Y(n_479)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_SL g472 ( 
.A(n_332),
.B(n_336),
.Y(n_472)
);

INVx6_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_335),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_336),
.B(n_377),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_336),
.B(n_407),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_SL g421 ( 
.A1(n_336),
.A2(n_406),
.B(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_344),
.Y(n_337)
);

MAJx2_ASAP7_75t_L g527 ( 
.A(n_338),
.B(n_345),
.C(n_352),
.Y(n_527)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_352),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_359),
.C(n_367),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_355),
.A2(n_356),
.B1(n_513),
.B2(n_514),
.Y(n_512)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_359),
.A2(n_367),
.B1(n_368),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_359),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx6_ASAP7_75t_L g402 ( 
.A(n_366),
.Y(n_402)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_382),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_369),
.A2(n_382),
.B1(n_383),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_384),
.Y(n_441)
);

OAI32xp33_ASAP7_75t_L g400 ( 
.A1(n_385),
.A2(n_401),
.A3(n_403),
.B1(n_406),
.B2(n_410),
.Y(n_400)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx6_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx6_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_394),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_510),
.B(n_516),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_490),
.B(n_509),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_453),
.B(n_489),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_431),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g489 ( 
.A(n_399),
.B(n_431),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_419),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_400),
.A2(n_419),
.B1(n_420),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_400),
.Y(n_466)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx5_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_414),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_442),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_432),
.B(n_444),
.C(n_452),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_433),
.Y(n_464)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_445),
.B2(n_452),
.Y(n_442)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_443),
.Y(n_452)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_467),
.B(n_488),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_465),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_455),
.B(n_465),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_484),
.B(n_487),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_473),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx4_ASAP7_75t_SL g482 ( 
.A(n_483),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_486),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_492),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_493),
.B(n_496),
.C(n_508),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_496),
.A2(n_497),
.B1(n_507),
.B2(n_508),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_512),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_511),
.B(n_512),
.Y(n_516)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_521),
.B(n_528),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_519),
.B(n_521),
.C(n_534),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.C(n_527),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g529 ( 
.A(n_522),
.B(n_530),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_525),
.B(n_527),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_529),
.B(n_531),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);


endmodule