module fake_jpeg_12969_n_185 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_185);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_1),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_25),
.B(n_1),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_46),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_10),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_25),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_26),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_47),
.B(n_49),
.Y(n_79)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_23),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_57),
.B(n_61),
.Y(n_90)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_37),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_31),
.B(n_19),
.C(n_18),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_19),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_32),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_39),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g71 ( 
.A(n_69),
.Y(n_71)
);

AND2x6_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_13),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_85),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_65),
.A2(n_40),
.B1(n_41),
.B2(n_39),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_74),
.A2(n_89),
.B1(n_30),
.B2(n_24),
.Y(n_101)
);

AO221x1_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_31),
.B1(n_37),
.B2(n_16),
.C(n_20),
.Y(n_75)
);

HAxp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_20),
.CON(n_109),
.SN(n_109)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_77),
.B(n_92),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_16),
.B(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_17),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_41),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_58),
.B1(n_51),
.B2(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_93),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_30),
.B1(n_24),
.B2(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_98),
.A2(n_109),
.B(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_90),
.A2(n_56),
.B1(n_55),
.B2(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_102),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_105),
.B1(n_113),
.B2(n_92),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_73),
.B(n_21),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_85),
.A2(n_55),
.B1(n_63),
.B2(n_60),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_60),
.B1(n_67),
.B2(n_30),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_52),
.B1(n_29),
.B2(n_22),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_79),
.B(n_22),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_70),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_80),
.A2(n_24),
.B1(n_29),
.B2(n_27),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_122),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_83),
.C(n_77),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_116),
.B(n_119),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_118),
.B1(n_99),
.B2(n_71),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_107),
.A2(n_72),
.B1(n_93),
.B2(n_87),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_86),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_78),
.C(n_82),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_76),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_100),
.C(n_103),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_111),
.A2(n_81),
.B(n_71),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_98),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_136),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_134),
.A2(n_125),
.B1(n_124),
.B2(n_120),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_129),
.B(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_138),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_140),
.B(n_143),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_144),
.B(n_146),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_127),
.B1(n_117),
.B2(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_78),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_155),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_132),
.B(n_151),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_141),
.B(n_119),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_154),
.C(n_155),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_128),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_101),
.Y(n_155)
);

OAI322xp33_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_127),
.A3(n_84),
.B1(n_124),
.B2(n_105),
.C1(n_20),
.C2(n_33),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_84),
.C(n_138),
.Y(n_163)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_152),
.B(n_144),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_154),
.Y(n_160)
);

OAI21x1_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_162),
.B(n_163),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g167 ( 
.A1(n_164),
.A2(n_165),
.B(n_137),
.C(n_145),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_136),
.B(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_133),
.Y(n_171)
);

OAI31xp33_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_147),
.A3(n_163),
.B(n_161),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_134),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_171),
.B(n_161),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_173),
.A2(n_174),
.B(n_175),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_156),
.B(n_135),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_133),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_172),
.A3(n_169),
.B1(n_91),
.B2(n_12),
.C1(n_14),
.C2(n_9),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_181),
.B(n_175),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_177),
.A2(n_11),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_110),
.C2(n_108),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_108),
.A3(n_3),
.B1(n_4),
.B2(n_7),
.C1(n_8),
.C2(n_2),
.Y(n_181)
);

OAI221xp5_ASAP7_75t_L g184 ( 
.A1(n_182),
.A2(n_178),
.B1(n_4),
.B2(n_7),
.C(n_3),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_183),
.Y(n_185)
);


endmodule