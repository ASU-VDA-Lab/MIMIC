module fake_jpeg_29930_n_106 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_44),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_36),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_43),
.B(n_40),
.C(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_29),
.B1(n_39),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_66)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_50),
.A2(n_31),
.B(n_2),
.C(n_3),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_47),
.A2(n_31),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_60),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_61),
.A2(n_49),
.B1(n_41),
.B2(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_69),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_70),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_8),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_10),
.Y(n_74)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_27),
.B1(n_14),
.B2(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_81),
.A2(n_83),
.B1(n_85),
.B2(n_77),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_63),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_82),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_69),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_83)
);

NAND2x1_ASAP7_75t_SL g84 ( 
.A(n_67),
.B(n_45),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

XNOR2x1_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_63),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_85),
.B1(n_82),
.B2(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_94),
.Y(n_95)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_92),
.Y(n_100)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_101),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_96),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

OAI311xp33_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_95),
.A3(n_89),
.B1(n_87),
.C1(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_81),
.Y(n_106)
);


endmodule