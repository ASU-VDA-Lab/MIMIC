module fake_jpeg_14121_n_650 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_650);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_650;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_398;
wire n_583;
wire n_56;
wire n_240;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_6),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_7),
.Y(n_53)
);

INVx11_ASAP7_75t_SL g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_62),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_17),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_65),
.B(n_125),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_69),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_70),
.Y(n_155)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_72),
.Y(n_184)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_73),
.Y(n_181)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_75),
.B(n_104),
.Y(n_148)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_77),
.B(n_82),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_79),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_80),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_39),
.B(n_0),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_83),
.Y(n_149)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_86),
.Y(n_211)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_88),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_89),
.Y(n_199)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_92),
.Y(n_151)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_93),
.Y(n_146)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_95),
.B(n_98),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g174 ( 
.A(n_96),
.Y(n_174)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_97),
.Y(n_169)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_100),
.Y(n_193)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx8_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_26),
.B(n_0),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_102),
.B(n_106),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_103),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_39),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_0),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_105),
.B(n_117),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_43),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_43),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_109),
.B(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_23),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_28),
.Y(n_166)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_25),
.Y(n_111)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_40),
.Y(n_115)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_115),
.Y(n_167)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_1),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_118),
.B(n_122),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_44),
.Y(n_120)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_19),
.B(n_60),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_24),
.Y(n_123)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_19),
.B(n_2),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_126),
.Y(n_187)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_25),
.Y(n_127)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_33),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_58),
.Y(n_182)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_36),
.Y(n_130)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_130),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_132),
.B(n_147),
.Y(n_236)
);

INVx13_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_74),
.B(n_60),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_138),
.B(n_150),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_115),
.A2(n_58),
.B1(n_41),
.B2(n_27),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_143),
.A2(n_161),
.B1(n_113),
.B2(n_108),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_79),
.B(n_32),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_32),
.B(n_30),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_156),
.A2(n_45),
.B(n_22),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_158),
.B(n_172),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_89),
.A2(n_48),
.B1(n_41),
.B2(n_27),
.Y(n_161)
);

INVx4_ASAP7_75t_SL g163 ( 
.A(n_71),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_163),
.B(n_164),
.Y(n_267)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_103),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_51),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_91),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_178),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_123),
.B(n_33),
.Y(n_179)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_179),
.B(n_29),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_182),
.B(n_212),
.Y(n_237)
);

BUFx4f_ASAP7_75t_SL g191 ( 
.A(n_72),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

BUFx12_ASAP7_75t_L g194 ( 
.A(n_88),
.Y(n_194)
);

CKINVDCx12_ASAP7_75t_R g240 ( 
.A(n_194),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_101),
.B(n_30),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_196),
.B(n_201),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_94),
.B(n_35),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_84),
.Y(n_203)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_120),
.A2(n_28),
.B1(n_24),
.B2(n_27),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_81),
.B1(n_80),
.B2(n_78),
.Y(n_232)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_126),
.Y(n_209)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_93),
.B(n_35),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_213),
.B(n_55),
.Y(n_272)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_66),
.Y(n_214)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_69),
.B(n_22),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_52),
.Y(n_277)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_199),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_220),
.Y(n_303)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_140),
.Y(n_221)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_221),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g222 ( 
.A(n_134),
.B(n_51),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_222),
.B(n_245),
.Y(n_321)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_223),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_224),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_226),
.A2(n_232),
.B1(n_281),
.B2(n_159),
.Y(n_348)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_227),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_133),
.Y(n_228)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_228),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_229),
.B(n_263),
.Y(n_344)
);

AOI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_166),
.A2(n_28),
.B(n_24),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_215),
.C(n_157),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_208),
.A2(n_107),
.B1(n_99),
.B2(n_86),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_231),
.A2(n_241),
.B1(n_280),
.B2(n_263),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_133),
.Y(n_234)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_177),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_284),
.Y(n_298)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_239),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_41),
.B1(n_48),
.B2(n_58),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_151),
.Y(n_244)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_244),
.Y(n_316)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_56),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_145),
.Y(n_246)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_146),
.Y(n_247)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_247),
.Y(n_310)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_185),
.Y(n_249)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_249),
.Y(n_317)
);

NAND2x1_ASAP7_75t_SL g250 ( 
.A(n_139),
.B(n_38),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_250),
.Y(n_353)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_202),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_251),
.Y(n_294)
);

CKINVDCx12_ASAP7_75t_R g252 ( 
.A(n_178),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_252),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_155),
.A2(n_48),
.B1(n_56),
.B2(n_38),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_253),
.A2(n_283),
.B1(n_292),
.B2(n_155),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_131),
.Y(n_254)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_254),
.Y(n_331)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_145),
.Y(n_255)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_255),
.Y(n_330)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_178),
.Y(n_259)
);

BUFx8_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_289),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_142),
.B(n_53),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_261),
.B(n_271),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_144),
.Y(n_262)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

AND2x2_ASAP7_75t_SL g263 ( 
.A(n_180),
.B(n_2),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g264 ( 
.A(n_204),
.B(n_42),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_264),
.B(n_286),
.Y(n_322)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_164),
.Y(n_265)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_265),
.Y(n_326)
);

INVx6_ASAP7_75t_L g266 ( 
.A(n_146),
.Y(n_266)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_266),
.Y(n_342)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_152),
.Y(n_268)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_210),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_277),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_136),
.Y(n_270)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_270),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_148),
.B(n_53),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_272),
.Y(n_334)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_163),
.Y(n_273)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_273),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_204),
.B(n_55),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_274),
.B(n_285),
.Y(n_319)
);

INVx5_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

INVx11_ASAP7_75t_L g309 ( 
.A(n_275),
.Y(n_309)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_184),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_276),
.Y(n_339)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_137),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_278),
.B(n_282),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_279),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_179),
.A2(n_52),
.B1(n_45),
.B2(n_49),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_L g281 ( 
.A1(n_143),
.A2(n_42),
.B1(n_49),
.B2(n_8),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

INVx8_ASAP7_75t_L g283 ( 
.A(n_144),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_177),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_195),
.B(n_4),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_141),
.B(n_4),
.Y(n_286)
);

INVx5_ASAP7_75t_L g287 ( 
.A(n_159),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_287),
.B(n_290),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_207),
.B(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_288),
.B(n_291),
.Y(n_343)
);

OR2x2_ASAP7_75t_SL g289 ( 
.A(n_170),
.B(n_149),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_175),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_154),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_153),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_281),
.A2(n_165),
.B1(n_193),
.B2(n_200),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_293),
.B(n_301),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_232),
.A2(n_171),
.B1(n_187),
.B2(n_188),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_304),
.A2(n_315),
.B1(n_345),
.B2(n_348),
.Y(n_355)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_242),
.B(n_174),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_306),
.B(n_325),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_307),
.A2(n_258),
.B(n_254),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_257),
.B(n_165),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_318),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_264),
.A2(n_215),
.B1(n_167),
.B2(n_157),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_237),
.B(n_173),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_235),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g394 ( 
.A1(n_327),
.A2(n_136),
.B1(n_258),
.B2(n_224),
.Y(n_394)
);

AO22x1_ASAP7_75t_SL g329 ( 
.A1(n_231),
.A2(n_189),
.B1(n_190),
.B2(n_193),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_335),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_267),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_333),
.B(n_337),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_222),
.B(n_200),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_236),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_289),
.B(n_192),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_341),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_279),
.B(n_192),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_253),
.A2(n_167),
.B1(n_188),
.B2(n_211),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_267),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_352),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_250),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_245),
.B(n_255),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g401 ( 
.A1(n_354),
.A2(n_390),
.B(n_372),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g356 ( 
.A(n_294),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_356),
.B(n_366),
.Y(n_404)
);

INVx13_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_358),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g359 ( 
.A(n_306),
.B(n_259),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_359),
.B(n_380),
.Y(n_437)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_301),
.A2(n_353),
.B1(n_336),
.B2(n_329),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_360),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_407)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_363),
.Y(n_421)
);

CKINVDCx11_ASAP7_75t_R g364 ( 
.A(n_340),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_364),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_343),
.Y(n_366)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_367),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_335),
.A2(n_307),
.B1(n_336),
.B2(n_329),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_293),
.A2(n_168),
.B1(n_227),
.B2(n_217),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_293),
.A2(n_168),
.B1(n_160),
.B2(n_176),
.Y(n_370)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_297),
.B(n_273),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_371),
.A2(n_391),
.B(n_392),
.Y(n_432)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_298),
.Y(n_373)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_344),
.B(n_225),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_376),
.C(n_238),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_341),
.B(n_233),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_381),
.Y(n_422)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx13_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_378),
.Y(n_423)
);

FAx1_ASAP7_75t_SL g380 ( 
.A(n_344),
.B(n_259),
.CI(n_219),
.CON(n_380),
.SN(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_332),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_318),
.B(n_243),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_387),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_304),
.A2(n_248),
.B1(n_283),
.B2(n_266),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_383),
.A2(n_310),
.B1(n_342),
.B2(n_349),
.Y(n_406)
);

INVx13_ASAP7_75t_L g384 ( 
.A(n_300),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_384),
.A2(n_394),
.B1(n_270),
.B2(n_218),
.Y(n_420)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_313),
.Y(n_385)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_385),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_322),
.A2(n_211),
.B1(n_176),
.B2(n_162),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_388),
.B1(n_342),
.B2(n_310),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_276),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_347),
.A2(n_293),
.B1(n_319),
.B2(n_334),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_328),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_L g431 ( 
.A1(n_389),
.A2(n_316),
.B1(n_323),
.B2(n_218),
.Y(n_431)
);

CKINVDCx14_ASAP7_75t_R g391 ( 
.A(n_321),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_311),
.B(n_265),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_330),
.Y(n_393)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_393),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_347),
.B(n_247),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_399),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_331),
.B(n_246),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_349),
.Y(n_408)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_330),
.Y(n_398)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_398),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_295),
.B(n_282),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_313),
.Y(n_400)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_400),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_401),
.Y(n_472)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_388),
.B(n_317),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_403),
.A2(n_395),
.B(n_387),
.C(n_364),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_406),
.A2(n_417),
.B1(n_428),
.B2(n_369),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_408),
.B(n_412),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_374),
.B(n_296),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_414),
.C(n_354),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_357),
.B(n_305),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_338),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g442 ( 
.A(n_415),
.B(n_427),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_365),
.A2(n_326),
.B(n_346),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_416),
.A2(n_426),
.B(n_397),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_362),
.A2(n_160),
.B1(n_162),
.B2(n_153),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_385),
.Y(n_424)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_365),
.A2(n_326),
.B(n_346),
.Y(n_426)
);

OAI22x1_ASAP7_75t_SL g428 ( 
.A1(n_355),
.A2(n_303),
.B1(n_314),
.B2(n_300),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_400),
.Y(n_430)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_430),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_383),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_395),
.A2(n_314),
.B1(n_312),
.B2(n_323),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_434),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_366),
.B(n_197),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_435),
.B(n_368),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_381),
.B(n_350),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_439),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_362),
.B(n_350),
.Y(n_439)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_441),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_444),
.A2(n_476),
.B1(n_407),
.B2(n_412),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_415),
.B(n_379),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g499 ( 
.A(n_447),
.Y(n_499)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_438),
.Y(n_450)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

INVx13_ASAP7_75t_L g451 ( 
.A(n_419),
.Y(n_451)
);

INVxp67_ASAP7_75t_SL g490 ( 
.A(n_451),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_371),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g488 ( 
.A(n_453),
.B(n_457),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_422),
.B(n_373),
.Y(n_454)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_454),
.Y(n_480)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_419),
.Y(n_455)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_455),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_456),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_392),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_416),
.B(n_395),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_459),
.B(n_461),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_376),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_410),
.C(n_414),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_396),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_462),
.B(n_464),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_422),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_463),
.B(n_474),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_423),
.B(n_403),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g465 ( 
.A(n_401),
.B(n_382),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_465),
.B(n_466),
.Y(n_510)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_408),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_419),
.Y(n_467)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_467),
.Y(n_483)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_468),
.Y(n_498)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_469),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_426),
.B(n_355),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_470),
.A2(n_477),
.B(n_429),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_404),
.B(n_375),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_471),
.B(n_411),
.Y(n_511)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_409),
.Y(n_473)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_473),
.Y(n_507)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_439),
.B(n_399),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_475),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_428),
.A2(n_370),
.B1(n_359),
.B2(n_386),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_489),
.C(n_494),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_436),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_481),
.Y(n_529)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_484),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_487),
.A2(n_458),
.B(n_448),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_460),
.B(n_435),
.C(n_433),
.Y(n_489)
);

INVx6_ASAP7_75t_L g491 ( 
.A(n_451),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_491),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_465),
.B(n_437),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_492),
.B(n_497),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_433),
.C(n_429),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_454),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_442),
.B(n_436),
.C(n_407),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_500),
.B(n_502),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_417),
.B1(n_406),
.B2(n_440),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_501),
.A2(n_476),
.B1(n_444),
.B2(n_477),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_459),
.B(n_408),
.C(n_397),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_471),
.B(n_425),
.Y(n_504)
);

CKINVDCx14_ASAP7_75t_R g527 ( 
.A(n_504),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_461),
.B(n_425),
.C(n_440),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_506),
.B(n_448),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_472),
.A2(n_411),
.B1(n_421),
.B2(n_380),
.Y(n_509)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_509),
.Y(n_515)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_511),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_513),
.A2(n_526),
.B1(n_532),
.B2(n_537),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_491),
.Y(n_516)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_463),
.Y(n_518)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_518),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_470),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_519),
.B(n_540),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_499),
.B(n_472),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_520),
.B(n_525),
.Y(n_548)
);

AND2x2_ASAP7_75t_SL g547 ( 
.A(n_521),
.B(n_487),
.Y(n_547)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_495),
.Y(n_522)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_522),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_488),
.A2(n_452),
.B1(n_450),
.B2(n_443),
.Y(n_524)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_524),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_480),
.B(n_443),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_503),
.A2(n_475),
.B1(n_452),
.B2(n_456),
.Y(n_526)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_495),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_530),
.B(n_531),
.Y(n_552)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_498),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_501),
.A2(n_448),
.B1(n_445),
.B2(n_469),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_533),
.B(n_541),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_486),
.B(n_468),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_535),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_496),
.B(n_363),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_478),
.B(n_500),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_536),
.B(n_542),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_479),
.A2(n_445),
.B1(n_446),
.B2(n_474),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_510),
.A2(n_446),
.B1(n_473),
.B2(n_455),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_538),
.A2(n_479),
.B1(n_483),
.B2(n_482),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_493),
.B(n_380),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_494),
.B(n_506),
.Y(n_541)
);

XNOR2x2_ASAP7_75t_SL g542 ( 
.A(n_481),
.B(n_377),
.Y(n_542)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_517),
.B(n_502),
.C(n_489),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_545),
.B(n_549),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_SL g546 ( 
.A1(n_539),
.A2(n_485),
.B(n_481),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_546),
.B(n_551),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_547),
.A2(n_523),
.B(n_367),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_517),
.B(n_485),
.C(n_482),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_514),
.A2(n_515),
.B1(n_512),
.B2(n_528),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_554),
.B(n_555),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_541),
.B(n_483),
.C(n_507),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_507),
.C(n_508),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_558),
.B(n_560),
.C(n_561),
.Y(n_572)
);

OAI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_512),
.A2(n_508),
.B1(n_505),
.B2(n_498),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_559),
.B(n_562),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_533),
.B(n_505),
.C(n_421),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_519),
.B(n_467),
.C(n_398),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_523),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_540),
.B(n_490),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_384),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_521),
.B(n_393),
.C(n_361),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_358),
.C(n_324),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_567),
.B(n_529),
.Y(n_568)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_568),
.Y(n_593)
);

AO221x1_ASAP7_75t_L g570 ( 
.A1(n_566),
.A2(n_550),
.B1(n_527),
.B2(n_553),
.C(n_564),
.Y(n_570)
);

CKINVDCx14_ASAP7_75t_R g589 ( 
.A(n_570),
.Y(n_589)
);

BUFx12_ASAP7_75t_L g571 ( 
.A(n_560),
.Y(n_571)
);

CKINVDCx14_ASAP7_75t_R g604 ( 
.A(n_571),
.Y(n_604)
);

CKINVDCx16_ASAP7_75t_R g573 ( 
.A(n_548),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_573),
.B(n_577),
.Y(n_603)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_552),
.A2(n_518),
.B(n_522),
.C(n_525),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_L g590 ( 
.A1(n_574),
.A2(n_556),
.B(n_561),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_547),
.A2(n_513),
.B1(n_532),
.B2(n_526),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_579),
.Y(n_596)
);

AOI321xp33_ASAP7_75t_L g577 ( 
.A1(n_547),
.A2(n_534),
.A3(n_542),
.B1(n_537),
.B2(n_449),
.C(n_378),
.Y(n_577)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_578),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_SL g579 ( 
.A(n_544),
.B(n_449),
.Y(n_579)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_580),
.A2(n_219),
.B(n_299),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_549),
.B(n_324),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_582),
.B(n_587),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_586),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g597 ( 
.A(n_584),
.B(n_588),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_556),
.A2(n_557),
.B1(n_558),
.B2(n_555),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_562),
.B(n_320),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_551),
.B(n_240),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g612 ( 
.A1(n_590),
.A2(n_594),
.B1(n_577),
.B2(n_571),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g594 ( 
.A1(n_585),
.A2(n_545),
.B1(n_563),
.B2(n_565),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_575),
.B(n_563),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_598),
.B(n_600),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_576),
.A2(n_544),
.B(n_320),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g609 ( 
.A1(n_599),
.A2(n_580),
.B(n_583),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_569),
.B(n_312),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_572),
.B(n_581),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_601),
.B(n_234),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_568),
.B(n_292),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_602),
.B(n_262),
.Y(n_615)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_299),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_174),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_606),
.A2(n_220),
.B1(n_275),
.B2(n_287),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_603),
.A2(n_592),
.B1(n_593),
.B2(n_568),
.Y(n_607)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_607),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_595),
.B(n_578),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_610),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_609),
.B(n_614),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_605),
.B(n_571),
.C(n_584),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_612),
.A2(n_596),
.B1(n_593),
.B2(n_597),
.Y(n_621)
);

AOI221xp5_ASAP7_75t_L g613 ( 
.A1(n_604),
.A2(n_574),
.B1(n_579),
.B2(n_588),
.C(n_299),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_613),
.B(n_616),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_591),
.Y(n_626)
);

BUFx24_ASAP7_75t_SL g617 ( 
.A(n_592),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_617),
.B(n_620),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g623 ( 
.A(n_618),
.B(n_597),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_590),
.B(n_228),
.C(n_191),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_619),
.B(n_606),
.C(n_596),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_589),
.B(n_4),
.Y(n_620)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_621),
.Y(n_632)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_623),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_626),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_611),
.B(n_591),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_628),
.B(n_630),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g629 ( 
.A1(n_612),
.A2(n_599),
.B(n_602),
.Y(n_629)
);

AOI21x1_ASAP7_75t_L g633 ( 
.A1(n_629),
.A2(n_619),
.B(n_610),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_633),
.A2(n_635),
.B(n_631),
.Y(n_639)
);

XOR2xp5_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_594),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_634),
.A2(n_622),
.B(n_623),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_625),
.A2(n_614),
.B1(n_135),
.B2(n_194),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_639),
.B(n_640),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_636),
.A2(n_630),
.B(n_622),
.Y(n_640)
);

AOI322xp5_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_642),
.A3(n_638),
.B1(n_637),
.B2(n_632),
.C1(n_635),
.C2(n_7),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_634),
.A2(n_624),
.B(n_9),
.Y(n_642)
);

OAI311xp33_ASAP7_75t_L g646 ( 
.A1(n_644),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.C1(n_13),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_643),
.B(n_9),
.C(n_10),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_645),
.A2(n_646),
.B(n_13),
.Y(n_647)
);

OAI21xp5_ASAP7_75t_SL g648 ( 
.A1(n_647),
.A2(n_10),
.B(n_11),
.Y(n_648)
);

XNOR2xp5_ASAP7_75t_L g649 ( 
.A(n_648),
.B(n_11),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_649),
.B(n_13),
.Y(n_650)
);


endmodule