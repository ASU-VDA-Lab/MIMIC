module real_aes_11601_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_488;
wire n_501;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1481;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_0), .Y(n_1117) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_1), .A2(n_496), .B1(n_499), .B2(n_508), .C(n_511), .Y(n_495) );
AOI21xp33_ASAP7_75t_L g566 ( .A1(n_1), .A2(n_567), .B(n_569), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g686 ( .A1(n_2), .A2(n_87), .B1(n_678), .B2(n_679), .Y(n_686) );
INVxp67_ASAP7_75t_SL g715 ( .A(n_2), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_3), .A2(n_73), .B1(n_1295), .B2(n_1307), .Y(n_1306) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_4), .Y(n_296) );
AND2x2_ASAP7_75t_L g386 ( .A(n_4), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g441 ( .A(n_4), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_4), .B(n_219), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_5), .A2(n_22), .B1(n_678), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_5), .A2(n_220), .B1(n_707), .B2(n_784), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_6), .Y(n_827) );
INVx1_ASAP7_75t_L g423 ( .A(n_7), .Y(n_423) );
AOI221xp5_ASAP7_75t_L g1050 ( .A1(n_8), .A2(n_175), .B1(n_322), .B2(n_642), .C(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1088 ( .A(n_8), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1107 ( .A1(n_9), .A2(n_1108), .B(n_1109), .C(n_1145), .Y(n_1107) );
OAI221xp5_ASAP7_75t_L g883 ( .A1(n_10), .A2(n_462), .B1(n_816), .B2(n_884), .C(n_890), .Y(n_883) );
INVx1_ASAP7_75t_L g906 ( .A(n_10), .Y(n_906) );
INVx1_ASAP7_75t_L g432 ( .A(n_11), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g1130 ( .A(n_12), .Y(n_1130) );
INVx1_ASAP7_75t_L g1587 ( .A(n_13), .Y(n_1587) );
OAI221xp5_ASAP7_75t_L g1603 ( .A1(n_13), .A2(n_462), .B1(n_816), .B2(n_1604), .C(n_1605), .Y(n_1603) );
OAI221xp5_ASAP7_75t_L g516 ( .A1(n_14), .A2(n_25), .B1(n_517), .B2(n_520), .C(n_521), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_14), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g878 ( .A1(n_15), .A2(n_62), .B1(n_437), .B2(n_522), .C(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g911 ( .A(n_15), .Y(n_911) );
INVx1_ASAP7_75t_L g873 ( .A(n_16), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_16), .A2(n_65), .B1(n_698), .B2(n_708), .Y(n_908) );
AO22x2_ASAP7_75t_L g915 ( .A1(n_17), .A2(n_916), .B1(n_971), .B2(n_972), .Y(n_915) );
CKINVDCx14_ASAP7_75t_R g971 ( .A(n_17), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_18), .A2(n_93), .B1(n_1054), .B2(n_1184), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_18), .A2(n_38), .B1(n_385), .B2(n_446), .Y(n_1211) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_19), .A2(n_83), .B1(n_1291), .B2(n_1295), .Y(n_1336) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_20), .Y(n_828) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_21), .A2(n_271), .B1(n_987), .B2(n_988), .C(n_990), .Y(n_986) );
INVx1_ASAP7_75t_L g1015 ( .A(n_21), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g779 ( .A1(n_22), .A2(n_99), .B1(n_630), .B2(n_780), .C(n_782), .Y(n_779) );
INVx1_ASAP7_75t_L g1612 ( .A(n_23), .Y(n_1612) );
OAI22xp33_ASAP7_75t_L g1622 ( .A1(n_23), .A2(n_34), .B1(n_1214), .B2(n_1216), .Y(n_1622) );
AOI221xp5_ASAP7_75t_L g1227 ( .A1(n_24), .A2(n_245), .B1(n_957), .B2(n_988), .C(n_1070), .Y(n_1227) );
INVx1_ASAP7_75t_L g1253 ( .A(n_24), .Y(n_1253) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_25), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g891 ( .A(n_26), .Y(n_891) );
INVx1_ASAP7_75t_L g805 ( .A(n_27), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_27), .A2(n_247), .B1(n_321), .B2(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g317 ( .A(n_28), .Y(n_317) );
OR2x2_ASAP7_75t_L g476 ( .A(n_28), .B(n_365), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g611 ( .A1(n_29), .A2(n_209), .B1(n_612), .B2(n_613), .C(n_615), .Y(n_611) );
INVx1_ASAP7_75t_L g625 ( .A(n_29), .Y(n_625) );
AO22x1_ASAP7_75t_L g868 ( .A1(n_30), .A2(n_869), .B1(n_913), .B2(n_914), .Y(n_868) );
INVx1_ASAP7_75t_L g914 ( .A(n_30), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1180 ( .A1(n_31), .A2(n_71), .B1(n_945), .B2(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1203 ( .A(n_31), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1206 ( .A1(n_32), .A2(n_171), .B1(n_437), .B2(n_758), .C(n_1207), .Y(n_1206) );
OAI22xp5_ASAP7_75t_L g1218 ( .A1(n_32), .A2(n_244), .B1(n_486), .B2(n_1219), .Y(n_1218) );
AOI22xp5_ASAP7_75t_L g1335 ( .A1(n_33), .A2(n_144), .B1(n_1279), .B2(n_1287), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g1614 ( .A1(n_34), .A2(n_142), .B1(n_530), .B2(n_1212), .C(n_1615), .Y(n_1614) );
OAI221xp5_ASAP7_75t_L g1118 ( .A1(n_35), .A2(n_229), .B1(n_1119), .B2(n_1120), .C(n_1121), .Y(n_1118) );
INVx1_ASAP7_75t_L g1158 ( .A(n_35), .Y(n_1158) );
BUFx2_ASAP7_75t_L g319 ( .A(n_36), .Y(n_319) );
BUFx2_ASAP7_75t_L g353 ( .A(n_36), .Y(n_353) );
INVx1_ASAP7_75t_L g367 ( .A(n_36), .Y(n_367) );
OR2x2_ASAP7_75t_L g519 ( .A(n_36), .B(n_448), .Y(n_519) );
AOI22xp33_ASAP7_75t_SL g762 ( .A1(n_37), .A2(n_169), .B1(n_682), .B2(n_683), .Y(n_762) );
INVxp33_ASAP7_75t_SL g789 ( .A(n_37), .Y(n_789) );
OAI222xp33_ASAP7_75t_L g1213 ( .A1(n_38), .A2(n_171), .B1(n_178), .B2(n_692), .C1(n_1214), .C2(n_1216), .Y(n_1213) );
INVx1_ASAP7_75t_L g1102 ( .A(n_39), .Y(n_1102) );
INVx1_ASAP7_75t_L g1327 ( .A(n_40), .Y(n_1327) );
INVx1_ASAP7_75t_L g919 ( .A(n_41), .Y(n_919) );
AOI21xp33_ASAP7_75t_L g961 ( .A1(n_41), .A2(n_698), .B(n_782), .Y(n_961) );
INVx1_ASAP7_75t_L g591 ( .A(n_42), .Y(n_591) );
INVxp33_ASAP7_75t_SL g753 ( .A(n_43), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_43), .A2(n_226), .B1(n_326), .B2(n_346), .C(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_44), .A2(n_185), .B1(n_449), .B2(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g557 ( .A(n_44), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g823 ( .A(n_45), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_46), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1230 ( .A1(n_47), .A2(n_76), .B1(n_994), .B2(n_1231), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_47), .A2(n_76), .B1(n_521), .B2(n_1018), .C(n_1019), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_48), .A2(n_205), .B1(n_678), .B2(n_679), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g716 ( .A1(n_48), .A2(n_263), .B1(n_346), .B2(n_717), .C(n_720), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_49), .A2(n_96), .B1(n_467), .B2(n_513), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_49), .A2(n_96), .B1(n_538), .B2(n_542), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g1598 ( .A1(n_50), .A2(n_64), .B1(n_358), .B2(n_370), .Y(n_1598) );
INVx1_ASAP7_75t_L g1619 ( .A(n_50), .Y(n_1619) );
INVx1_ASAP7_75t_L g1384 ( .A(n_51), .Y(n_1384) );
OAI221xp5_ASAP7_75t_L g962 ( .A1(n_52), .A2(n_236), .B1(n_963), .B2(n_964), .C(n_966), .Y(n_962) );
INVx1_ASAP7_75t_L g969 ( .A(n_52), .Y(n_969) );
INVx1_ASAP7_75t_L g889 ( .A(n_53), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_53), .A2(n_162), .B1(n_322), .B2(n_708), .Y(n_904) );
INVx1_ASAP7_75t_L g601 ( .A(n_54), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_55), .A2(n_180), .B1(n_834), .B2(n_881), .Y(n_880) );
OAI22xp5_ASAP7_75t_SL g897 ( .A1(n_55), .A2(n_180), .B1(n_358), .B2(n_370), .Y(n_897) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_56), .Y(n_368) );
INVx1_ASAP7_75t_L g1191 ( .A(n_57), .Y(n_1191) );
OAI221xp5_ASAP7_75t_L g1209 ( .A1(n_57), .A2(n_94), .B1(n_834), .B2(n_881), .C(n_1210), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_58), .A2(n_1107), .B1(n_1170), .B2(n_1171), .Y(n_1106) );
INVx1_ASAP7_75t_L g1171 ( .A(n_58), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_59), .A2(n_110), .B1(n_1279), .B2(n_1287), .Y(n_1278) );
INVx1_ASAP7_75t_L g502 ( .A(n_60), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_60), .A2(n_554), .B(n_555), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_61), .A2(n_101), .B1(n_682), .B2(n_683), .Y(n_685) );
INVxp33_ASAP7_75t_SL g729 ( .A(n_61), .Y(n_729) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_62), .A2(n_121), .B1(n_478), .B2(n_486), .Y(n_912) );
INVx1_ASAP7_75t_L g1591 ( .A(n_63), .Y(n_1591) );
OAI211xp5_ASAP7_75t_L g1610 ( .A1(n_63), .A2(n_392), .B(n_1611), .C(n_1616), .Y(n_1610) );
INVx1_ASAP7_75t_L g1617 ( .A(n_64), .Y(n_1617) );
INVx1_ASAP7_75t_L g874 ( .A(n_65), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g1527 ( .A1(n_66), .A2(n_123), .B1(n_1528), .B2(n_1529), .Y(n_1527) );
AOI221xp5_ASAP7_75t_L g1552 ( .A1(n_66), .A2(n_150), .B1(n_555), .B2(n_1553), .C(n_1555), .Y(n_1552) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_67), .Y(n_1066) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_68), .A2(n_217), .B1(n_346), .B2(n_347), .Y(n_345) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_68), .A2(n_278), .B1(n_382), .B2(n_392), .Y(n_381) );
AO22x2_ASAP7_75t_L g794 ( .A1(n_69), .A2(n_795), .B1(n_796), .B2(n_865), .Y(n_794) );
INVx1_ASAP7_75t_L g865 ( .A(n_69), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_70), .Y(n_830) );
INVx1_ASAP7_75t_L g1201 ( .A(n_71), .Y(n_1201) );
INVx1_ASAP7_75t_L g1116 ( .A(n_72), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1164 ( .A1(n_72), .A2(n_145), .B1(n_854), .B2(n_1165), .C(n_1167), .Y(n_1164) );
CKINVDCx5p33_ASAP7_75t_R g375 ( .A(n_74), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_75), .A2(n_124), .B1(n_1279), .B2(n_1287), .Y(n_1309) );
INVxp33_ASAP7_75t_SL g1520 ( .A(n_77), .Y(n_1520) );
AOI22xp33_ASAP7_75t_SL g1547 ( .A1(n_77), .A2(n_221), .B1(n_322), .B2(n_708), .Y(n_1547) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_78), .A2(n_211), .B1(n_799), .B2(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g857 ( .A1(n_78), .A2(n_211), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_79), .A2(n_272), .B1(n_561), .B2(n_1241), .Y(n_1240) );
INVx1_ASAP7_75t_L g1258 ( .A(n_79), .Y(n_1258) );
AOI221xp5_ASAP7_75t_L g596 ( .A1(n_80), .A2(n_149), .B1(n_425), .B2(n_597), .C(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_80), .A2(n_97), .B1(n_636), .B2(n_637), .Y(n_635) );
CKINVDCx5p33_ASAP7_75t_R g821 ( .A(n_81), .Y(n_821) );
INVx1_ASAP7_75t_L g1139 ( .A(n_82), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_82), .A2(n_257), .B1(n_542), .B2(n_545), .Y(n_1168) );
INVxp67_ASAP7_75t_SL g1518 ( .A(n_84), .Y(n_1518) );
OAI221xp5_ASAP7_75t_L g1544 ( .A1(n_84), .A2(n_224), .B1(n_964), .B2(n_994), .C(n_1545), .Y(n_1544) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_85), .A2(n_255), .B1(n_540), .B2(n_849), .Y(n_991) );
INVx1_ASAP7_75t_L g1016 ( .A(n_85), .Y(n_1016) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_86), .Y(n_505) );
INVxp33_ASAP7_75t_L g727 ( .A(n_87), .Y(n_727) );
INVx1_ASAP7_75t_L g600 ( .A(n_88), .Y(n_600) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_88), .A2(n_149), .B1(n_630), .B2(n_631), .C(n_633), .Y(n_629) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_89), .Y(n_832) );
INVx1_ASAP7_75t_L g1596 ( .A(n_90), .Y(n_1596) );
OAI22xp5_ASAP7_75t_L g1602 ( .A1(n_90), .A2(n_164), .B1(n_799), .B2(n_800), .Y(n_1602) );
INVx1_ASAP7_75t_L g316 ( .A(n_91), .Y(n_316) );
INVx1_ASAP7_75t_L g365 ( .A(n_91), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_92), .A2(n_266), .B1(n_644), .B2(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1094 ( .A(n_92), .Y(n_1094) );
INVx1_ASAP7_75t_L g1208 ( .A(n_93), .Y(n_1208) );
INVx1_ASAP7_75t_L g1190 ( .A(n_94), .Y(n_1190) );
INVx1_ASAP7_75t_L g616 ( .A(n_95), .Y(n_616) );
OAI221xp5_ASAP7_75t_L g620 ( .A1(n_95), .A2(n_209), .B1(n_621), .B2(n_623), .C(n_624), .Y(n_620) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_97), .Y(n_599) );
INVxp67_ASAP7_75t_SL g658 ( .A(n_98), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g699 ( .A1(n_98), .A2(n_235), .B1(n_700), .B2(n_702), .Y(n_699) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_99), .A2(n_220), .B1(n_682), .B2(n_760), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g818 ( .A1(n_100), .A2(n_392), .B1(n_819), .B2(n_824), .C(n_829), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g853 ( .A1(n_100), .A2(n_138), .B1(n_854), .B2(n_856), .Y(n_853) );
INVxp67_ASAP7_75t_SL g696 ( .A(n_101), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g531 ( .A1(n_102), .A2(n_170), .B1(n_532), .B2(n_535), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_102), .A2(n_228), .B1(n_323), .B2(n_561), .Y(n_565) );
INVx1_ASAP7_75t_L g608 ( .A(n_103), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_103), .A2(n_160), .B1(n_569), .B2(n_641), .C(n_642), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g1305 ( .A1(n_104), .A2(n_128), .B1(n_1279), .B2(n_1287), .Y(n_1305) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_105), .A2(n_228), .B1(n_525), .B2(n_528), .Y(n_524) );
INVx1_ASAP7_75t_L g563 ( .A(n_105), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_106), .A2(n_223), .B1(n_1279), .B2(n_1287), .Y(n_1298) );
INVxp33_ASAP7_75t_SL g1524 ( .A(n_107), .Y(n_1524) );
AOI21xp33_ASAP7_75t_L g1548 ( .A1(n_107), .A2(n_777), .B(n_1549), .Y(n_1548) );
AOI22xp5_ASAP7_75t_L g1290 ( .A1(n_108), .A2(n_146), .B1(n_1291), .B2(n_1295), .Y(n_1290) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_109), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_111), .A2(n_738), .B1(n_739), .B2(n_793), .Y(n_737) );
INVx1_ASAP7_75t_L g793 ( .A(n_111), .Y(n_793) );
INVx1_ASAP7_75t_L g1315 ( .A(n_112), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_112), .A2(n_1566), .B1(n_1568), .B2(n_1623), .Y(n_1565) );
XNOR2xp5_ASAP7_75t_L g1570 ( .A(n_112), .B(n_1571), .Y(n_1570) );
OAI21xp33_ASAP7_75t_L g582 ( .A1(n_113), .A2(n_583), .B(n_618), .Y(n_582) );
INVx1_ASAP7_75t_L g652 ( .A(n_113), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g1182 ( .A1(n_114), .A2(n_188), .B1(n_719), .B2(n_987), .Y(n_1182) );
AOI21xp33_ASAP7_75t_L g1199 ( .A1(n_114), .A2(n_449), .B(n_509), .Y(n_1199) );
INVx1_ASAP7_75t_L g617 ( .A(n_115), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_116), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g997 ( .A1(n_117), .A2(n_238), .B1(n_555), .B2(n_988), .C(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1028 ( .A(n_117), .Y(n_1028) );
INVx1_ASAP7_75t_L g1144 ( .A(n_118), .Y(n_1144) );
OAI211xp5_ASAP7_75t_SL g1146 ( .A1(n_118), .A2(n_1147), .B(n_1148), .C(n_1154), .Y(n_1146) );
INVx1_ASAP7_75t_L g752 ( .A(n_119), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_120), .A2(n_155), .B1(n_679), .B2(n_1537), .Y(n_1536) );
INVxp33_ASAP7_75t_SL g1559 ( .A(n_120), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_121), .A2(n_139), .B1(n_612), .B2(n_877), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_122), .A2(n_143), .B1(n_678), .B2(n_764), .Y(n_763) );
INVxp33_ASAP7_75t_L g788 ( .A(n_122), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_123), .A2(n_125), .B1(n_326), .B2(n_1557), .Y(n_1556) );
AOI22xp33_ASAP7_75t_L g1531 ( .A1(n_125), .A2(n_150), .B1(n_1532), .B2(n_1533), .Y(n_1531) );
INVx1_ASAP7_75t_L g814 ( .A(n_126), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_126), .A2(n_148), .B1(n_851), .B2(n_852), .Y(n_850) );
INVx1_ASAP7_75t_L g288 ( .A(n_127), .Y(n_288) );
AO22x1_ASAP7_75t_SL g1312 ( .A1(n_129), .A2(n_231), .B1(n_1279), .B2(n_1287), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g1007 ( .A(n_130), .Y(n_1007) );
CKINVDCx5p33_ASAP7_75t_R g1244 ( .A(n_131), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g929 ( .A(n_132), .Y(n_929) );
OA22x2_ASAP7_75t_L g981 ( .A1(n_133), .A2(n_982), .B1(n_1040), .B2(n_1041), .Y(n_981) );
INVx1_ASAP7_75t_L g1041 ( .A(n_133), .Y(n_1041) );
INVx1_ASAP7_75t_L g1268 ( .A(n_134), .Y(n_1268) );
AO221x2_ASAP7_75t_L g1321 ( .A1(n_135), .A2(n_274), .B1(n_1307), .B2(n_1322), .C(n_1323), .Y(n_1321) );
INVxp67_ASAP7_75t_SL g744 ( .A(n_136), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_136), .A2(n_281), .B1(n_700), .B2(n_702), .Y(n_771) );
OAI221xp5_ASAP7_75t_SL g604 ( .A1(n_137), .A2(n_254), .B1(n_605), .B2(n_606), .C(n_607), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_137), .A2(n_254), .B1(n_322), .B2(n_644), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_138), .A2(n_462), .B1(n_802), .B2(n_808), .C(n_816), .Y(n_801) );
INVx1_ASAP7_75t_L g910 ( .A(n_139), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g1228 ( .A1(n_140), .A2(n_215), .B1(n_1065), .B2(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1250 ( .A(n_140), .Y(n_1250) );
AOI22xp33_ASAP7_75t_L g1535 ( .A1(n_141), .A2(n_197), .B1(n_1532), .B2(n_1533), .Y(n_1535) );
INVxp67_ASAP7_75t_SL g1543 ( .A(n_141), .Y(n_1543) );
OAI22xp33_ASAP7_75t_L g1621 ( .A1(n_142), .A2(n_172), .B1(n_486), .B2(n_1219), .Y(n_1621) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_143), .Y(n_786) );
XOR2xp5_ASAP7_75t_L g492 ( .A(n_144), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g1114 ( .A(n_145), .Y(n_1114) );
INVx1_ASAP7_75t_L g1522 ( .A(n_147), .Y(n_1522) );
INVx1_ASAP7_75t_L g811 ( .A(n_148), .Y(n_811) );
INVx1_ASAP7_75t_L g750 ( .A(n_151), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g1072 ( .A(n_152), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g1577 ( .A(n_153), .Y(n_1577) );
CKINVDCx5p33_ASAP7_75t_R g935 ( .A(n_154), .Y(n_935) );
INVxp67_ASAP7_75t_SL g1551 ( .A(n_155), .Y(n_1551) );
CKINVDCx5p33_ASAP7_75t_R g1006 ( .A(n_156), .Y(n_1006) );
AOI221xp5_ASAP7_75t_L g1069 ( .A1(n_157), .A2(n_279), .B1(n_642), .B2(n_957), .C(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g1077 ( .A(n_157), .Y(n_1077) );
XNOR2xp5_ASAP7_75t_L g1175 ( .A(n_158), .B(n_1176), .Y(n_1175) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_159), .A2(n_265), .B1(n_321), .B2(n_326), .Y(n_320) );
INVx1_ASAP7_75t_L g405 ( .A(n_159), .Y(n_405) );
INVx1_ASAP7_75t_L g610 ( .A(n_160), .Y(n_610) );
INVx1_ASAP7_75t_L g1060 ( .A(n_161), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1080 ( .A1(n_161), .A2(n_251), .B1(n_520), .B2(n_1081), .C(n_1083), .Y(n_1080) );
INVx1_ASAP7_75t_L g887 ( .A(n_162), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g1243 ( .A(n_163), .Y(n_1243) );
INVx1_ASAP7_75t_L g1594 ( .A(n_164), .Y(n_1594) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_165), .A2(n_268), .B1(n_1291), .B2(n_1295), .Y(n_1299) );
INVx1_ASAP7_75t_L g920 ( .A(n_166), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g960 ( .A1(n_166), .A2(n_214), .B1(n_708), .B2(n_785), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g1511 ( .A1(n_167), .A2(n_1512), .B1(n_1513), .B2(n_1561), .Y(n_1511) );
CKINVDCx5p33_ASAP7_75t_R g1512 ( .A(n_167), .Y(n_1512) );
CKINVDCx5p33_ASAP7_75t_R g1234 ( .A(n_168), .Y(n_1234) );
INVxp67_ASAP7_75t_SL g770 ( .A(n_169), .Y(n_770) );
INVx1_ASAP7_75t_L g571 ( .A(n_170), .Y(n_571) );
INVx1_ASAP7_75t_L g1613 ( .A(n_172), .Y(n_1613) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_173), .Y(n_1049) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_174), .Y(n_693) );
INVx1_ASAP7_75t_L g1091 ( .A(n_175), .Y(n_1091) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_176), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_177), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1205 ( .A1(n_178), .A2(n_244), .B1(n_597), .B2(n_877), .Y(n_1205) );
CKINVDCx5p33_ASAP7_75t_R g1579 ( .A(n_179), .Y(n_1579) );
AOI22xp33_ASAP7_75t_SL g1185 ( .A1(n_181), .A2(n_194), .B1(n_327), .B2(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1194 ( .A(n_181), .Y(n_1194) );
INVxp67_ASAP7_75t_SL g1134 ( .A(n_182), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_182), .A2(n_212), .B1(n_630), .B2(n_780), .C(n_1153), .Y(n_1152) );
XOR2x2_ASAP7_75t_L g653 ( .A(n_183), .B(n_654), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_184), .A2(n_278), .B1(n_333), .B2(n_339), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g461 ( .A1(n_184), .A2(n_217), .B1(n_462), .B2(n_465), .Y(n_461) );
INVx1_ASAP7_75t_L g552 ( .A(n_185), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g938 ( .A1(n_186), .A2(n_207), .B1(n_939), .B2(n_940), .Y(n_938) );
INVx1_ASAP7_75t_L g951 ( .A(n_186), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g941 ( .A1(n_187), .A2(n_232), .B1(n_532), .B2(n_535), .Y(n_941) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_187), .A2(n_207), .B1(n_698), .B2(n_708), .Y(n_954) );
INVx1_ASAP7_75t_L g1198 ( .A(n_188), .Y(n_1198) );
AOI221xp5_ASAP7_75t_L g1235 ( .A1(n_189), .A2(n_248), .B1(n_1236), .B2(n_1238), .C(n_1239), .Y(n_1235) );
INVx1_ASAP7_75t_L g1261 ( .A(n_189), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_190), .A2(n_258), .B1(n_1295), .B2(n_1307), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g930 ( .A(n_191), .Y(n_930) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_192), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_192), .B(n_288), .Y(n_1286) );
AND3x2_ASAP7_75t_L g1292 ( .A(n_192), .B(n_288), .C(n_1283), .Y(n_1292) );
OA332x1_ASAP7_75t_L g917 ( .A1(n_193), .A2(n_496), .A3(n_508), .B1(n_918), .B2(n_923), .B3(n_927), .C1(n_931), .C2(n_936), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g955 ( .A1(n_193), .A2(n_956), .B(n_957), .Y(n_955) );
INVx1_ASAP7_75t_L g1195 ( .A(n_194), .Y(n_1195) );
INVx2_ASAP7_75t_L g301 ( .A(n_195), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_196), .A2(n_260), .B1(n_987), .B2(n_1000), .Y(n_999) );
INVx1_ASAP7_75t_L g1024 ( .A(n_196), .Y(n_1024) );
INVxp33_ASAP7_75t_SL g1560 ( .A(n_197), .Y(n_1560) );
INVx1_ASAP7_75t_L g1582 ( .A(n_198), .Y(n_1582) );
AOI21xp33_ASAP7_75t_L g1607 ( .A1(n_198), .A2(n_509), .B(n_1608), .Y(n_1607) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_199), .Y(n_1003) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_200), .Y(n_669) );
OAI211xp5_ASAP7_75t_L g871 ( .A1(n_201), .A2(n_392), .B(n_872), .C(n_875), .Y(n_871) );
INVx1_ASAP7_75t_L g907 ( .A(n_201), .Y(n_907) );
INVx1_ASAP7_75t_L g587 ( .A(n_202), .Y(n_587) );
INVxp33_ASAP7_75t_SL g671 ( .A(n_203), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_203), .A2(n_249), .B1(n_705), .B2(n_707), .C(n_709), .Y(n_704) );
INVx1_ASAP7_75t_L g1317 ( .A(n_204), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_205), .A2(n_225), .B1(n_644), .B2(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g1283 ( .A(n_206), .Y(n_1283) );
INVx1_ASAP7_75t_L g1600 ( .A(n_208), .Y(n_1600) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_210), .A2(n_275), .B1(n_449), .B2(n_507), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_210), .A2(n_275), .B1(n_545), .B2(n_547), .Y(n_544) );
INVxp67_ASAP7_75t_SL g1126 ( .A(n_212), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_213), .A2(n_259), .B1(n_333), .B2(n_339), .Y(n_332) );
INVx1_ASAP7_75t_L g417 ( .A(n_213), .Y(n_417) );
INVx1_ASAP7_75t_L g924 ( .A(n_214), .Y(n_924) );
INVx1_ASAP7_75t_L g1254 ( .A(n_215), .Y(n_1254) );
CKINVDCx5p33_ASAP7_75t_R g1226 ( .A(n_216), .Y(n_1226) );
CKINVDCx20_ASAP7_75t_R g1324 ( .A(n_218), .Y(n_1324) );
INVx1_ASAP7_75t_L g303 ( .A(n_219), .Y(n_303) );
INVx2_ASAP7_75t_L g387 ( .A(n_219), .Y(n_387) );
INVxp33_ASAP7_75t_SL g1525 ( .A(n_221), .Y(n_1525) );
INVx1_ASAP7_75t_L g895 ( .A(n_222), .Y(n_895) );
INVxp67_ASAP7_75t_SL g1517 ( .A(n_224), .Y(n_1517) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_225), .A2(n_263), .B1(n_682), .B2(n_683), .Y(n_681) );
INVxp33_ASAP7_75t_SL g748 ( .A(n_226), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g1379 ( .A1(n_227), .A2(n_230), .B1(n_1380), .B2(n_1381), .C(n_1382), .Y(n_1379) );
INVx1_ASAP7_75t_L g1160 ( .A(n_229), .Y(n_1160) );
INVx1_ASAP7_75t_L g967 ( .A(n_232), .Y(n_967) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_233), .Y(n_1057) );
INVx1_ASAP7_75t_L g452 ( .A(n_234), .Y(n_452) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_235), .Y(n_661) );
INVx1_ASAP7_75t_L g970 ( .A(n_236), .Y(n_970) );
XOR2xp5_ASAP7_75t_L g308 ( .A(n_237), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g1025 ( .A(n_238), .Y(n_1025) );
CKINVDCx5p33_ASAP7_75t_R g992 ( .A(n_239), .Y(n_992) );
INVx1_ASAP7_75t_L g666 ( .A(n_240), .Y(n_666) );
INVx1_ASAP7_75t_L g428 ( .A(n_241), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g1058 ( .A(n_242), .Y(n_1058) );
INVx1_ASAP7_75t_L g1132 ( .A(n_243), .Y(n_1132) );
INVx1_ASAP7_75t_L g1251 ( .A(n_245), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g993 ( .A1(n_246), .A2(n_253), .B1(n_994), .B2(n_995), .Y(n_993) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_246), .A2(n_253), .B1(n_1018), .B2(n_1019), .C(n_1020), .Y(n_1017) );
INVx1_ASAP7_75t_L g807 ( .A(n_247), .Y(n_807) );
INVx1_ASAP7_75t_L g1259 ( .A(n_248), .Y(n_1259) );
INVxp33_ASAP7_75t_SL g663 ( .A(n_249), .Y(n_663) );
INVx1_ASAP7_75t_L g1284 ( .A(n_250), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_250), .B(n_1282), .Y(n_1289) );
INVx1_ASAP7_75t_L g1061 ( .A(n_251), .Y(n_1061) );
INVx1_ASAP7_75t_L g1073 ( .A(n_252), .Y(n_1073) );
INVx1_ASAP7_75t_L g1012 ( .A(n_255), .Y(n_1012) );
INVx1_ASAP7_75t_L g1136 ( .A(n_256), .Y(n_1136) );
OAI211xp5_ASAP7_75t_L g1155 ( .A1(n_256), .A2(n_1156), .B(n_1157), .C(n_1161), .Y(n_1155) );
INVx1_ASAP7_75t_L g1141 ( .A(n_257), .Y(n_1141) );
INVx1_ASAP7_75t_L g413 ( .A(n_259), .Y(n_413) );
INVx1_ASAP7_75t_L g1030 ( .A(n_260), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g892 ( .A(n_261), .Y(n_892) );
INVx2_ASAP7_75t_L g300 ( .A(n_262), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g1068 ( .A(n_264), .Y(n_1068) );
INVx1_ASAP7_75t_L g399 ( .A(n_265), .Y(n_399) );
INVx1_ASAP7_75t_L g1086 ( .A(n_266), .Y(n_1086) );
CKINVDCx5p33_ASAP7_75t_R g925 ( .A(n_267), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g1584 ( .A(n_269), .Y(n_1584) );
CKINVDCx5p33_ASAP7_75t_R g1112 ( .A(n_270), .Y(n_1112) );
INVx1_ASAP7_75t_L g1013 ( .A(n_271), .Y(n_1013) );
INVx1_ASAP7_75t_L g1263 ( .A(n_272), .Y(n_1263) );
INVx1_ASAP7_75t_L g1245 ( .A(n_273), .Y(n_1245) );
BUFx3_ASAP7_75t_L g325 ( .A(n_276), .Y(n_325) );
INVx1_ASAP7_75t_L g331 ( .A(n_276), .Y(n_331) );
INVx1_ASAP7_75t_L g324 ( .A(n_277), .Y(n_324) );
BUFx3_ASAP7_75t_L g330 ( .A(n_277), .Y(n_330) );
INVx1_ASAP7_75t_L g1079 ( .A(n_279), .Y(n_1079) );
INVx1_ASAP7_75t_L g1540 ( .A(n_280), .Y(n_1540) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_281), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_304), .B(n_1271), .Y(n_282) );
HB1xp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_291), .Y(n_285) );
AND2x4_ASAP7_75t_L g1567 ( .A(n_286), .B(n_292), .Y(n_1567) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_287), .B(n_289), .Y(n_286) );
INVx1_ASAP7_75t_SL g1564 ( .A(n_287), .Y(n_1564) );
NAND2xp5_ASAP7_75t_L g1627 ( .A(n_287), .B(n_289), .Y(n_1627) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g1563 ( .A(n_289), .B(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_293), .B(n_297), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g420 ( .A(n_295), .B(n_303), .Y(n_420) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g509 ( .A(n_296), .B(n_510), .Y(n_509) );
OR2x6_ASAP7_75t_L g297 ( .A(n_298), .B(n_302), .Y(n_297) );
BUFx2_ASAP7_75t_L g416 ( .A(n_298), .Y(n_416) );
INVx1_ASAP7_75t_L g434 ( .A(n_298), .Y(n_434) );
OR2x2_ASAP7_75t_L g535 ( .A(n_298), .B(n_519), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g598 ( .A1(n_298), .A2(n_430), .B1(n_599), .B2(n_600), .Y(n_598) );
OAI22xp33_ASAP7_75t_L g615 ( .A1(n_298), .A2(n_430), .B1(n_616), .B2(n_617), .Y(n_615) );
INVx2_ASAP7_75t_SL g813 ( .A(n_298), .Y(n_813) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_298), .Y(n_928) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x4_ASAP7_75t_L g390 ( .A(n_300), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_300), .Y(n_396) );
INVx2_ASAP7_75t_L g404 ( .A(n_300), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_300), .Y(n_412) );
AND2x2_ASAP7_75t_L g451 ( .A(n_300), .B(n_301), .Y(n_451) );
INVx2_ASAP7_75t_L g391 ( .A(n_301), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_301), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g411 ( .A(n_301), .Y(n_411) );
INVx1_ASAP7_75t_L g458 ( .A(n_301), .Y(n_458) );
INVx1_ASAP7_75t_L g469 ( .A(n_301), .Y(n_469) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_975), .B1(n_976), .B2(n_1270), .Y(n_304) );
INVx2_ASAP7_75t_L g1270 ( .A(n_305), .Y(n_1270) );
XNOR2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_735), .Y(n_305) );
AO22x2_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_653), .B1(n_733), .B2(n_734), .Y(n_306) );
INVx1_ASAP7_75t_L g733 ( .A(n_307), .Y(n_733) );
XNOR2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_491), .Y(n_307) );
NAND4xp75_ASAP7_75t_L g309 ( .A(n_310), .B(n_380), .C(n_472), .D(n_481), .Y(n_309) );
AND2x2_ASAP7_75t_SL g310 ( .A(n_311), .B(n_356), .Y(n_310) );
AOI33xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_320), .A3(n_332), .B1(n_344), .B2(n_345), .B3(n_350), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_313), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_313), .Y(n_847) );
OR2x6_ASAP7_75t_L g313 ( .A(n_314), .B(n_318), .Y(n_313) );
INVx1_ASAP7_75t_L g1052 ( .A(n_314), .Y(n_1052) );
OR2x2_ASAP7_75t_L g1574 ( .A(n_314), .B(n_318), .Y(n_1574) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g555 ( .A(n_315), .Y(n_555) );
BUFx3_ASAP7_75t_L g634 ( .A(n_315), .Y(n_634) );
INVx1_ASAP7_75t_L g782 ( .A(n_315), .Y(n_782) );
INVx1_ASAP7_75t_L g900 ( .A(n_315), .Y(n_900) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x4_ASAP7_75t_L g354 ( .A(n_316), .B(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_317), .Y(n_355) );
AND2x2_ASAP7_75t_L g515 ( .A(n_318), .B(n_438), .Y(n_515) );
AND2x4_ASAP7_75t_L g595 ( .A(n_318), .B(n_420), .Y(n_595) );
INVx2_ASAP7_75t_L g648 ( .A(n_318), .Y(n_648) );
AND2x4_ASAP7_75t_L g676 ( .A(n_318), .B(n_420), .Y(n_676) );
BUFx2_ASAP7_75t_L g792 ( .A(n_318), .Y(n_792) );
OR2x2_ASAP7_75t_L g899 ( .A(n_318), .B(n_900), .Y(n_899) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
BUFx2_ASAP7_75t_L g471 ( .A(n_319), .Y(n_471) );
OR2x6_ASAP7_75t_L g508 ( .A(n_319), .B(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx3_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
INVx1_ASAP7_75t_L g706 ( .A(n_322), .Y(n_706) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_SL g484 ( .A(n_323), .Y(n_484) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_323), .Y(n_540) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_323), .Y(n_554) );
BUFx6f_ASAP7_75t_L g698 ( .A(n_323), .Y(n_698) );
BUFx2_ASAP7_75t_L g998 ( .A(n_323), .Y(n_998) );
BUFx2_ASAP7_75t_L g1065 ( .A(n_323), .Y(n_1065) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_323), .Y(n_1163) );
BUFx3_ASAP7_75t_L g1186 ( .A(n_323), .Y(n_1186) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g490 ( .A(n_324), .Y(n_490) );
INVx2_ASAP7_75t_L g337 ( .A(n_325), .Y(n_337) );
AND2x2_ASAP7_75t_L g343 ( .A(n_325), .B(n_330), .Y(n_343) );
BUFx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x6_ASAP7_75t_L g478 ( .A(n_328), .B(n_475), .Y(n_478) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_328), .B(n_475), .Y(n_1219) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_329), .Y(n_349) );
INVx2_ASAP7_75t_L g543 ( .A(n_329), .Y(n_543) );
BUFx6f_ASAP7_75t_L g708 ( .A(n_329), .Y(n_708) );
INVx1_ASAP7_75t_L g1578 ( .A(n_329), .Y(n_1578) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
INVx1_ASAP7_75t_L g489 ( .A(n_331), .Y(n_489) );
BUFx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g473 ( .A(n_334), .B(n_474), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_334), .A2(n_571), .B(n_572), .C(n_578), .Y(n_570) );
INVx2_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g723 ( .A(n_335), .Y(n_723) );
INVx1_ASAP7_75t_L g956 ( .A(n_335), .Y(n_956) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g480 ( .A(n_336), .B(n_363), .Y(n_480) );
INVx6_ASAP7_75t_L g568 ( .A(n_336), .Y(n_568) );
BUFx2_ASAP7_75t_L g1241 ( .A(n_336), .Y(n_1241) );
AND2x4_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
AND2x4_ASAP7_75t_L g724 ( .A(n_341), .B(n_725), .Y(n_724) );
BUFx6f_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g378 ( .A(n_342), .Y(n_378) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_342), .Y(n_642) );
INVx2_ASAP7_75t_L g989 ( .A(n_342), .Y(n_989) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_343), .Y(n_549) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g623 ( .A(n_349), .Y(n_623) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_349), .Y(n_644) );
BUFx6f_ASAP7_75t_L g945 ( .A(n_349), .Y(n_945) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_SL g898 ( .A1(n_351), .A2(n_899), .B1(n_901), .B2(n_905), .Y(n_898) );
INVx4_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx4f_ASAP7_75t_L g861 ( .A(n_352), .Y(n_861) );
AND2x4_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
AND2x4_ASAP7_75t_L g479 ( .A(n_353), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g1187 ( .A(n_353), .B(n_354), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_354), .Y(n_569) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_354), .Y(n_712) );
INVx2_ASAP7_75t_L g777 ( .A(n_354), .Y(n_777) );
INVx2_ASAP7_75t_SL g957 ( .A(n_354), .Y(n_957) );
INVx1_ASAP7_75t_L g990 ( .A(n_354), .Y(n_990) );
AND2x4_ASAP7_75t_L g363 ( .A(n_355), .B(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_368), .B1(n_369), .B2(n_375), .C(n_376), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_357), .A2(n_830), .B1(n_832), .B2(n_845), .Y(n_844) );
AOI221xp5_ASAP7_75t_L g1188 ( .A1(n_357), .A2(n_376), .B1(n_1189), .B2(n_1190), .C(n_1191), .Y(n_1188) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
OR2x2_ASAP7_75t_L g702 ( .A(n_359), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_360), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_574) );
AND2x4_ASAP7_75t_L g627 ( .A(n_360), .B(n_363), .Y(n_627) );
AND2x2_ASAP7_75t_L g965 ( .A(n_360), .B(n_363), .Y(n_965) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_360), .B(n_363), .Y(n_1062) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_SL g374 ( .A(n_362), .Y(n_374) );
INVx1_ASAP7_75t_L g379 ( .A(n_362), .Y(n_379) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .Y(n_362) );
BUFx2_ASAP7_75t_L g579 ( .A(n_363), .Y(n_579) );
AND2x4_ASAP7_75t_L g626 ( .A(n_363), .B(n_575), .Y(n_626) );
AND2x4_ASAP7_75t_L g701 ( .A(n_363), .B(n_575), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_363), .Y(n_703) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x6_ASAP7_75t_L g688 ( .A(n_366), .B(n_439), .Y(n_688) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g475 ( .A(n_367), .B(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g498 ( .A(n_367), .B(n_386), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_368), .A2(n_375), .B1(n_456), .B2(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g845 ( .A(n_370), .Y(n_845) );
INVx2_ASAP7_75t_L g1189 ( .A(n_370), .Y(n_1189) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_371), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g575 ( .A(n_372), .Y(n_575) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g896 ( .A(n_376), .B(n_897), .C(n_898), .Y(n_896) );
NOR3xp33_ASAP7_75t_L g1572 ( .A(n_376), .B(n_1573), .C(n_1598), .Y(n_1572) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
HB1xp67_ASAP7_75t_L g1555 ( .A(n_377), .Y(n_1555) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_379), .B(n_719), .Y(n_864) );
OAI31xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_397), .A3(n_461), .B(n_470), .Y(n_380) );
INVx3_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx3_ASAP7_75t_L g800 ( .A(n_383), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_383), .A2(n_466), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI221x1_ASAP7_75t_L g1193 ( .A1(n_383), .A2(n_466), .B1(n_1194), .B2(n_1195), .C(n_1196), .Y(n_1193) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_388), .Y(n_383) );
AND2x4_ASAP7_75t_L g393 ( .A(n_384), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g463 ( .A(n_386), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g466 ( .A(n_386), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g440 ( .A(n_387), .Y(n_440) );
INVx1_ASAP7_75t_L g510 ( .A(n_387), .Y(n_510) );
INVx1_ASAP7_75t_L g1202 ( .A(n_388), .Y(n_1202) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g513 ( .A(n_389), .Y(n_513) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_390), .Y(n_407) );
INVx3_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
AND2x4_ASAP7_75t_L g395 ( .A(n_391), .B(n_396), .Y(n_395) );
INVx8_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI221xp5_ASAP7_75t_SL g1204 ( .A1(n_393), .A2(n_1205), .B1(n_1206), .B2(n_1208), .C(n_1209), .Y(n_1204) );
BUFx6f_ASAP7_75t_L g758 ( .A(n_394), .Y(n_758) );
BUFx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_395), .Y(n_507) );
BUFx3_ASAP7_75t_L g522 ( .A(n_395), .Y(n_522) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_395), .Y(n_530) );
BUFx2_ASAP7_75t_L g593 ( .A(n_395), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_408), .B1(n_421), .B2(n_429), .C(n_442), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_405), .B2(n_406), .Y(n_398) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_SL g422 ( .A(n_401), .Y(n_422) );
BUFx3_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g605 ( .A(n_402), .Y(n_605) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g501 ( .A(n_403), .Y(n_501) );
BUFx2_ASAP7_75t_L g886 ( .A(n_403), .Y(n_886) );
INVx1_ASAP7_75t_L g460 ( .A(n_404), .Y(n_460) );
AND2x4_ASAP7_75t_L g467 ( .A(n_404), .B(n_468), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g931 ( .A1(n_406), .A2(n_932), .B1(n_933), .B2(n_935), .Y(n_931) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_SL g684 ( .A(n_407), .Y(n_684) );
INVx4_ASAP7_75t_L g761 ( .A(n_407), .Y(n_761) );
INVx2_ASAP7_75t_SL g806 ( .A(n_407), .Y(n_806) );
INVx2_ASAP7_75t_SL g1534 ( .A(n_407), .Y(n_1534) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_414), .B2(n_417), .C(n_418), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx3_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
BUFx2_ASAP7_75t_L g810 ( .A(n_410), .Y(n_810) );
INVx2_ASAP7_75t_L g817 ( .A(n_410), .Y(n_817) );
AND2x2_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_411), .B(n_412), .Y(n_431) );
INVx1_ASAP7_75t_L g590 ( .A(n_412), .Y(n_590) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g1023 ( .A(n_415), .Y(n_1023) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_SL g815 ( .A(n_420), .Y(n_815) );
OAI22xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_423), .B1(n_424), .B2(n_428), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_423), .A2(n_432), .B1(n_482), .B2(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g877 ( .A(n_426), .Y(n_877) );
INVx3_ASAP7_75t_L g1138 ( .A(n_426), .Y(n_1138) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g504 ( .A(n_427), .Y(n_504) );
INVx3_ASAP7_75t_L g534 ( .A(n_427), .Y(n_534) );
AOI222xp33_ASAP7_75t_L g472 ( .A1(n_428), .A2(n_435), .B1(n_452), .B2(n_473), .C1(n_477), .C2(n_479), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_432), .B1(n_433), .B2(n_435), .C(n_436), .Y(n_429) );
BUFx3_ASAP7_75t_L g926 ( .A(n_430), .Y(n_926) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_430), .A2(n_928), .B1(n_929), .B2(n_930), .Y(n_927) );
INVx2_ASAP7_75t_L g1101 ( .A(n_430), .Y(n_1101) );
BUFx3_ASAP7_75t_L g1606 ( .A(n_430), .Y(n_1606) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g822 ( .A(n_434), .Y(n_822) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_436), .A2(n_820), .B1(n_821), .B2(n_822), .C(n_823), .Y(n_819) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx2_ASAP7_75t_L g1615 ( .A(n_439), .Y(n_1615) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_452), .B(n_453), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NOR2xp67_ASAP7_75t_L g838 ( .A(n_444), .B(n_648), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_449), .Y(n_444) );
AND2x2_ASAP7_75t_L g831 ( .A(n_445), .B(n_586), .Y(n_831) );
AND2x2_ASAP7_75t_L g1618 ( .A(n_445), .B(n_586), .Y(n_1618) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_446), .A2(n_454), .B(n_455), .Y(n_453) );
OR2x6_ASAP7_75t_L g816 ( .A(n_446), .B(n_817), .Y(n_816) );
OR2x6_ASAP7_75t_L g834 ( .A(n_446), .B(n_460), .Y(n_834) );
INVx1_ASAP7_75t_L g882 ( .A(n_446), .Y(n_882) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g497 ( .A(n_449), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_SL g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g609 ( .A(n_450), .Y(n_609) );
INVx2_ASAP7_75t_L g1212 ( .A(n_450), .Y(n_1212) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_451), .Y(n_464) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_454), .A2(n_812), .B1(n_815), .B2(n_891), .C(n_892), .Y(n_890) );
INVx1_ASAP7_75t_L g1143 ( .A(n_454), .Y(n_1143) );
OAI21xp5_ASAP7_75t_SL g1197 ( .A1(n_454), .A2(n_1198), .B(n_1199), .Y(n_1197) );
NAND2x1_ASAP7_75t_SL g517 ( .A(n_456), .B(n_518), .Y(n_517) );
NAND2x1p5_ASAP7_75t_L g881 ( .A(n_456), .B(n_882), .Y(n_881) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_458), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g520 ( .A(n_459), .B(n_518), .Y(n_520) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
CKINVDCx6p67_ASAP7_75t_R g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g879 ( .A(n_464), .Y(n_879) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_464), .Y(n_1207) );
INVx3_ASAP7_75t_L g1609 ( .A(n_464), .Y(n_1609) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g799 ( .A(n_466), .Y(n_799) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_467), .Y(n_527) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_467), .Y(n_597) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_467), .Y(n_612) );
BUFx2_ASAP7_75t_L g1532 ( .A(n_467), .Y(n_1532) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g580 ( .A(n_470), .Y(n_580) );
BUFx8_ASAP7_75t_SL g893 ( .A(n_470), .Y(n_893) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g732 ( .A(n_471), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_473), .A2(n_482), .B1(n_823), .B2(n_827), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g909 ( .A1(n_473), .A2(n_482), .B1(n_910), .B2(n_911), .C(n_912), .Y(n_909) );
AND2x2_ASAP7_75t_L g482 ( .A(n_474), .B(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OR2x6_ASAP7_75t_L g486 ( .A(n_475), .B(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_475), .B(n_1215), .Y(n_1214) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_475), .B(n_1217), .Y(n_1216) );
INVx2_ASAP7_75t_L g541 ( .A(n_476), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_476), .B(n_543), .Y(n_542) );
OR2x2_ASAP7_75t_L g545 ( .A(n_476), .B(n_546), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g943 ( .A1(n_476), .A2(n_944), .B(n_946), .C(n_948), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_477), .A2(n_485), .B1(n_821), .B2(n_828), .Y(n_841) );
CKINVDCx6p67_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g692 ( .A(n_479), .Y(n_692) );
OR2x6_ASAP7_75t_L g837 ( .A(n_479), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g646 ( .A(n_480), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g966 ( .A(n_480), .B(n_967), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_483), .A2(n_930), .B1(n_932), .B2(n_947), .Y(n_946) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g630 ( .A(n_484), .Y(n_630) );
INVx2_ASAP7_75t_SL g1181 ( .A(n_484), .Y(n_1181) );
CKINVDCx6p67_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
OAI21xp33_ASAP7_75t_L g551 ( .A1(n_487), .A2(n_552), .B(n_553), .Y(n_551) );
OAI221xp5_ASAP7_75t_L g709 ( .A1(n_487), .A2(n_666), .B1(n_669), .B2(n_710), .C(n_712), .Y(n_709) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g564 ( .A(n_488), .Y(n_564) );
INVx1_ASAP7_75t_L g573 ( .A(n_488), .Y(n_573) );
BUFx2_ASAP7_75t_L g775 ( .A(n_488), .Y(n_775) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_488), .Y(n_903) );
INVx1_ASAP7_75t_L g1590 ( .A(n_488), .Y(n_1590) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
OR2x2_ASAP7_75t_L g546 ( .A(n_489), .B(n_490), .Y(n_546) );
XNOR2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_581), .Y(n_491) );
NAND3xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_523), .C(n_536), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_516), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x2_ASAP7_75t_L g526 ( .A(n_498), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g529 ( .A(n_498), .B(n_530), .Y(n_529) );
AND2x2_ASAP7_75t_L g533 ( .A(n_498), .B(n_534), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g603 ( .A1(n_498), .A2(n_515), .B1(n_604), .B2(n_611), .Y(n_603) );
AND2x4_ASAP7_75t_L g665 ( .A(n_498), .B(n_504), .Y(n_665) );
AND2x6_ASAP7_75t_L g667 ( .A(n_498), .B(n_522), .Y(n_667) );
AND2x4_ASAP7_75t_L g670 ( .A(n_498), .B(n_609), .Y(n_670) );
AND2x2_ASAP7_75t_L g672 ( .A(n_498), .B(n_527), .Y(n_672) );
AND2x2_ASAP7_75t_L g754 ( .A(n_498), .B(n_527), .Y(n_754) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_502), .B1(n_503), .B2(n_505), .C(n_506), .Y(n_499) );
INVx1_ASAP7_75t_L g826 ( .A(n_500), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g1611 ( .A1(n_500), .A2(n_806), .B1(n_1612), .B2(n_1613), .C(n_1614), .Y(n_1611) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g934 ( .A(n_501), .Y(n_934) );
INVx1_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g606 ( .A(n_504), .Y(n_606) );
INVx1_ASAP7_75t_L g888 ( .A(n_504), .Y(n_888) );
BUFx3_ASAP7_75t_L g1266 ( .A(n_504), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_505), .A2(n_557), .B1(n_558), .B2(n_560), .Y(n_556) );
OAI33xp33_ASAP7_75t_L g1021 ( .A1(n_508), .A2(n_1022), .A3(n_1026), .B1(n_1031), .B2(n_1035), .B3(n_1038), .Y(n_1021) );
OAI33xp33_ASAP7_75t_L g1084 ( .A1(n_508), .A2(n_1038), .A3(n_1085), .B1(n_1089), .B2(n_1095), .B3(n_1097), .Y(n_1084) );
OAI33xp33_ASAP7_75t_L g1122 ( .A1(n_508), .A2(n_1038), .A3(n_1123), .B1(n_1131), .B2(n_1135), .B3(n_1140), .Y(n_1122) );
OAI33xp33_ASAP7_75t_L g1256 ( .A1(n_508), .A2(n_688), .A3(n_1257), .B1(n_1260), .B2(n_1264), .B3(n_1267), .Y(n_1256) );
NAND3xp33_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .C(n_515), .Y(n_511) );
INVx1_ASAP7_75t_L g1262 ( .A(n_513), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1018 ( .A(n_517), .Y(n_1018) );
INVx2_ASAP7_75t_L g1082 ( .A(n_517), .Y(n_1082) );
NAND2x1p5_ASAP7_75t_L g521 ( .A(n_518), .B(n_522), .Y(n_521) );
AND2x4_ASAP7_75t_L g585 ( .A(n_518), .B(n_586), .Y(n_585) );
AND2x4_ASAP7_75t_L g588 ( .A(n_518), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g592 ( .A(n_518), .B(n_593), .Y(n_592) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx4f_ASAP7_75t_L g1019 ( .A(n_520), .Y(n_1019) );
BUFx4f_ASAP7_75t_L g1120 ( .A(n_520), .Y(n_1120) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_521), .Y(n_1020) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_521), .Y(n_1083) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_521), .Y(n_1121) );
NOR2xp33_ASAP7_75t_SL g523 ( .A(n_524), .B(n_531), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g939 ( .A(n_526), .Y(n_939) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g940 ( .A(n_529), .Y(n_940) );
INVx2_ASAP7_75t_SL g680 ( .A(n_530), .Y(n_680) );
BUFx6f_ASAP7_75t_L g764 ( .A(n_530), .Y(n_764) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g614 ( .A(n_534), .Y(n_614) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_534), .Y(n_922) );
INVx2_ASAP7_75t_L g1029 ( .A(n_534), .Y(n_1029) );
INVx2_ASAP7_75t_L g1034 ( .A(n_534), .Y(n_1034) );
INVx1_ASAP7_75t_L g1129 ( .A(n_534), .Y(n_1129) );
INVx2_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
AND2x4_ASAP7_75t_L g691 ( .A(n_535), .B(n_692), .Y(n_691) );
OAI31xp33_ASAP7_75t_SL g536 ( .A1(n_537), .A2(n_544), .A3(n_550), .B(n_580), .Y(n_536) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g985 ( .A1(n_539), .A2(n_986), .B1(n_991), .B2(n_992), .C(n_993), .Y(n_985) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_541), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_540), .A2(n_549), .B1(n_617), .B2(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g1217 ( .A(n_540), .Y(n_1217) );
BUFx4f_ASAP7_75t_L g1238 ( .A(n_540), .Y(n_1238) );
AND2x4_ASAP7_75t_L g548 ( .A(n_541), .B(n_549), .Y(n_548) );
AOI222xp33_ASAP7_75t_L g619 ( .A1(n_541), .A2(n_587), .B1(n_591), .B2(n_620), .C1(n_626), .C2(n_627), .Y(n_619) );
AND2x4_ASAP7_75t_L g697 ( .A(n_541), .B(n_698), .Y(n_697) );
INVx4_ASAP7_75t_L g730 ( .A(n_542), .Y(n_730) );
INVx1_ASAP7_75t_L g561 ( .A(n_543), .Y(n_561) );
INVx2_ASAP7_75t_L g1002 ( .A(n_543), .Y(n_1002) );
INVx6_ASAP7_75t_L g728 ( .A(n_545), .Y(n_728) );
INVx1_ASAP7_75t_L g559 ( .A(n_546), .Y(n_559) );
INVx1_ASAP7_75t_L g622 ( .A(n_546), .Y(n_622) );
INVx2_ASAP7_75t_L g711 ( .A(n_546), .Y(n_711) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_548), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g996 ( .A1(n_548), .A2(n_638), .B1(n_997), .B2(n_999), .C(n_1003), .Y(n_996) );
AOI221xp5_ASAP7_75t_L g1048 ( .A1(n_548), .A2(n_638), .B1(n_1049), .B2(n_1050), .C(n_1053), .Y(n_1048) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_548), .Y(n_1233) );
INVx2_ASAP7_75t_SL g632 ( .A(n_549), .Y(n_632) );
AND2x4_ASAP7_75t_L g638 ( .A(n_549), .B(n_579), .Y(n_638) );
BUFx6f_ASAP7_75t_L g719 ( .A(n_549), .Y(n_719) );
INVx1_ASAP7_75t_L g781 ( .A(n_549), .Y(n_781) );
BUFx3_ASAP7_75t_L g856 ( .A(n_549), .Y(n_856) );
BUFx4f_ASAP7_75t_L g947 ( .A(n_549), .Y(n_947) );
INVx1_ASAP7_75t_L g1237 ( .A(n_549), .Y(n_1237) );
OAI211xp5_ASAP7_75t_SL g550 ( .A1(n_551), .A2(n_556), .B(n_562), .C(n_570), .Y(n_550) );
INVx2_ASAP7_75t_L g1554 ( .A(n_554), .Y(n_1554) );
INVx2_ASAP7_75t_SL g1576 ( .A(n_554), .Y(n_1576) );
INVx1_ASAP7_75t_L g1593 ( .A(n_554), .Y(n_1593) );
INVx1_ASAP7_75t_L g721 ( .A(n_555), .Y(n_721) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_555), .Y(n_1153) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_558), .A2(n_750), .B1(n_752), .B2(n_774), .C(n_776), .Y(n_773) );
OAI221xp5_ASAP7_75t_L g905 ( .A1(n_558), .A2(n_902), .B1(n_906), .B2(n_907), .C(n_908), .Y(n_905) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OAI211xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B(n_565), .C(n_566), .Y(n_562) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_567), .Y(n_636) );
INVx1_ASAP7_75t_L g855 ( .A(n_567), .Y(n_855) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_L g641 ( .A(n_568), .Y(n_641) );
INVx1_ASAP7_75t_L g785 ( .A(n_568), .Y(n_785) );
INVx1_ASAP7_75t_L g987 ( .A(n_568), .Y(n_987) );
BUFx6f_ASAP7_75t_L g1055 ( .A(n_568), .Y(n_1055) );
INVx2_ASAP7_75t_SL g1549 ( .A(n_568), .Y(n_1549) );
NAND2xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g953 ( .A(n_573), .Y(n_953) );
BUFx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_649), .Y(n_581) );
INVx1_ASAP7_75t_L g651 ( .A(n_583), .Y(n_651) );
NAND3xp33_ASAP7_75t_SL g583 ( .A(n_584), .B(n_594), .C(n_603), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g584 ( .A1(n_585), .A2(n_587), .B1(n_588), .B2(n_591), .C(n_592), .Y(n_584) );
INVx1_ASAP7_75t_L g660 ( .A(n_585), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_585), .A2(n_742), .B1(n_744), .B2(n_745), .C(n_746), .Y(n_741) );
AOI221xp5_ASAP7_75t_L g968 ( .A1(n_585), .A2(n_588), .B1(n_592), .B2(n_969), .C(n_970), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g1516 ( .A1(n_585), .A2(n_588), .B1(n_592), .B2(n_1517), .C(n_1518), .Y(n_1516) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_588), .Y(n_657) );
INVx1_ASAP7_75t_L g743 ( .A(n_588), .Y(n_743) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_592), .A2(n_657), .B1(n_658), .B2(n_659), .C(n_661), .Y(n_656) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_592), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_593), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g1530 ( .A(n_593), .Y(n_1530) );
AOI22xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_596), .B1(n_601), .B2(n_602), .Y(n_594) );
AOI33xp33_ASAP7_75t_L g1526 ( .A1(n_595), .A2(n_687), .A3(n_1527), .B1(n_1531), .B2(n_1535), .B3(n_1536), .Y(n_1526) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_601), .A2(n_640), .B1(n_643), .B2(n_645), .Y(n_639) );
INVx2_ASAP7_75t_L g804 ( .A(n_605), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g1200 ( .A1(n_605), .A2(n_1201), .B1(n_1202), .B2(n_1203), .Y(n_1200) );
BUFx3_ASAP7_75t_L g678 ( .A(n_609), .Y(n_678) );
BUFx3_ASAP7_75t_L g682 ( .A(n_612), .Y(n_682) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g650 ( .A(n_618), .Y(n_650) );
AOI31xp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_628), .A3(n_639), .B(n_647), .Y(n_618) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g637 ( .A(n_623), .Y(n_637) );
INVx2_ASAP7_75t_L g994 ( .A(n_626), .Y(n_994) );
INVx2_ASAP7_75t_SL g995 ( .A(n_627), .Y(n_995) );
INVx2_ASAP7_75t_L g1231 ( .A(n_627), .Y(n_1231) );
AOI21xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_635), .B(n_638), .Y(n_628) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g852 ( .A(n_632), .Y(n_852) );
INVxp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g1239 ( .A(n_634), .Y(n_1239) );
INVx1_ASAP7_75t_L g948 ( .A(n_638), .Y(n_948) );
AOI221xp5_ASAP7_75t_L g1232 ( .A1(n_638), .A2(n_1233), .B1(n_1234), .B2(n_1235), .C(n_1240), .Y(n_1232) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_641), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_641), .A2(n_929), .B1(n_935), .B2(n_945), .Y(n_944) );
BUFx3_ASAP7_75t_L g1557 ( .A(n_641), .Y(n_1557) );
INVx1_ASAP7_75t_L g1067 ( .A(n_644), .Y(n_1067) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g1169 ( .A(n_647), .Y(n_1169) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_648), .A2(n_984), .B1(n_1007), .B2(n_1008), .Y(n_983) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .C(n_652), .Y(n_649) );
INVx2_ASAP7_75t_L g734 ( .A(n_653), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_655), .B(n_689), .Y(n_654) );
AND4x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_662), .C(n_668), .D(n_673), .Y(n_655) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_666), .B2(n_667), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_664), .A2(n_667), .B1(n_1068), .B2(n_1077), .Y(n_1076) );
BUFx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g749 ( .A(n_665), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_665), .A2(n_667), .B1(n_1012), .B2(n_1013), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1113 ( .A(n_665), .Y(n_1113) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_665), .A2(n_667), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
BUFx2_ASAP7_75t_L g1521 ( .A(n_665), .Y(n_1521) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_667), .A2(n_748), .B1(n_749), .B2(n_750), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_667), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_667), .A2(n_1520), .B1(n_1521), .B2(n_1522), .Y(n_1519) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_671), .B2(n_672), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_670), .A2(n_752), .B1(n_753), .B2(n_754), .Y(n_751) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_670), .A2(n_672), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_670), .A2(n_754), .B1(n_1066), .B2(n_1079), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g1115 ( .A1(n_670), .A2(n_672), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_670), .A2(n_672), .B1(n_1253), .B2(n_1254), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1523 ( .A1(n_670), .A2(n_672), .B1(n_1524), .B2(n_1525), .Y(n_1523) );
AOI33xp33_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_677), .A3(n_681), .B1(n_685), .B2(n_686), .B3(n_687), .Y(n_673) );
AOI33xp33_ASAP7_75t_L g755 ( .A1(n_674), .A2(n_687), .A3(n_756), .B1(n_759), .B2(n_762), .B3(n_763), .Y(n_755) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g824 ( .A1(n_684), .A2(n_825), .B1(n_827), .B2(n_828), .Y(n_824) );
INVx1_ASAP7_75t_L g936 ( .A(n_687), .Y(n_936) );
INVx6_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx5_ASAP7_75t_L g1039 ( .A(n_688), .Y(n_1039) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_693), .B(n_694), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_690), .A2(n_1046), .B1(n_1047), .B2(n_1073), .Y(n_1045) );
INVx1_ASAP7_75t_L g1108 ( .A(n_690), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g1539 ( .A1(n_690), .A2(n_1540), .B(n_1541), .Y(n_1539) );
INVx5_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g766 ( .A(n_691), .Y(n_766) );
INVx2_ASAP7_75t_SL g1008 ( .A(n_691), .Y(n_1008) );
INVx2_ASAP7_75t_L g1246 ( .A(n_691), .Y(n_1246) );
AOI31xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_713), .A3(n_726), .B(n_731), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B(n_699), .C(n_704), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g769 ( .A1(n_697), .A2(n_770), .B(n_771), .C(n_772), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_697), .B(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1156 ( .A(n_697), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1225 ( .A1(n_697), .A2(n_1226), .B1(n_1227), .B2(n_1228), .C(n_1230), .Y(n_1225) );
AOI21xp33_ASAP7_75t_SL g1542 ( .A1(n_697), .A2(n_1543), .B(n_1544), .Y(n_1542) );
BUFx3_ASAP7_75t_L g858 ( .A(n_698), .Y(n_858) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_SL g963 ( .A(n_701), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_701), .A2(n_1060), .B1(n_1061), .B2(n_1062), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_701), .A2(n_1158), .B1(n_1159), .B2(n_1160), .Y(n_1157) );
INVx1_ASAP7_75t_L g1159 ( .A(n_702), .Y(n_1159) );
INVx1_ASAP7_75t_SL g725 ( .A(n_703), .Y(n_725) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
BUFx3_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_708), .Y(n_849) );
INVx1_ASAP7_75t_L g860 ( .A(n_708), .Y(n_860) );
INVx1_ASAP7_75t_L g1595 ( .A(n_708), .Y(n_1595) );
OAI221xp5_ASAP7_75t_L g901 ( .A1(n_710), .A2(n_891), .B1(n_892), .B2(n_902), .C(n_904), .Y(n_901) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_711), .Y(n_1150) );
INVx1_ASAP7_75t_L g1215 ( .A(n_711), .Y(n_1215) );
INVx2_ASAP7_75t_L g1581 ( .A(n_711), .Y(n_1581) );
INVx2_ASAP7_75t_L g1586 ( .A(n_711), .Y(n_1586) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_715), .B1(n_716), .B2(n_722), .C(n_724), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g778 ( .A1(n_714), .A2(n_724), .B1(n_779), .B2(n_783), .C(n_786), .Y(n_778) );
INVx1_ASAP7_75t_L g1147 ( .A(n_714), .Y(n_1147) );
AOI221xp5_ASAP7_75t_L g1550 ( .A1(n_714), .A2(n_724), .B1(n_1551), .B2(n_1552), .C(n_1556), .Y(n_1550) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g1166 ( .A(n_719), .Y(n_1166) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g1154 ( .A(n_724), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_728), .A2(n_730), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g1004 ( .A1(n_728), .A2(n_730), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_728), .A2(n_730), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1242 ( .A1(n_728), .A2(n_730), .B1(n_1243), .B2(n_1244), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1558 ( .A1(n_728), .A2(n_730), .B1(n_1559), .B2(n_1560), .Y(n_1558) );
INVx1_ASAP7_75t_L g1046 ( .A(n_731), .Y(n_1046) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI31xp33_ASAP7_75t_L g942 ( .A1(n_732), .A2(n_943), .A3(n_949), .B(n_962), .Y(n_942) );
AOI21x1_ASAP7_75t_L g1192 ( .A1(n_732), .A2(n_1193), .B(n_1204), .Y(n_1192) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_866), .B1(n_973), .B2(n_974), .Y(n_735) );
INVx1_ASAP7_75t_L g973 ( .A(n_736), .Y(n_973) );
XNOR2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_794), .Y(n_736) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_765), .Y(n_739) );
AND4x1_ASAP7_75t_L g740 ( .A(n_741), .B(n_747), .C(n_751), .D(n_755), .Y(n_740) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
AOI21xp33_ASAP7_75t_SL g765 ( .A1(n_766), .A2(n_767), .B(n_768), .Y(n_765) );
AOI31xp33_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_778), .A3(n_787), .B(n_790), .Y(n_768) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx2_ASAP7_75t_SL g1583 ( .A(n_775), .Y(n_1583) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
BUFx2_ASAP7_75t_L g1167 ( .A(n_777), .Y(n_1167) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
HB1xp67_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI31xp33_ASAP7_75t_L g1541 ( .A1(n_790), .A2(n_1542), .A3(n_1550), .B(n_1558), .Y(n_1541) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
CKINVDCx8_ASAP7_75t_R g791 ( .A(n_792), .Y(n_791) );
OAI31xp33_ASAP7_75t_L g797 ( .A1(n_792), .A2(n_798), .A3(n_801), .B(n_818), .Y(n_797) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
NAND3xp33_ASAP7_75t_SL g796 ( .A(n_797), .B(n_835), .C(n_839), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g802 ( .A1(n_803), .A2(n_805), .B1(n_806), .B2(n_807), .Y(n_802) );
INVx2_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx2_ASAP7_75t_L g1090 ( .A(n_804), .Y(n_1090) );
INVx1_ASAP7_75t_L g1096 ( .A(n_804), .Y(n_1096) );
OAI221xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_811), .B1(n_812), .B2(n_814), .C(n_815), .Y(n_808) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g820 ( .A(n_810), .Y(n_820) );
INVx1_ASAP7_75t_L g1087 ( .A(n_810), .Y(n_1087) );
OAI22xp33_ASAP7_75t_L g923 ( .A1(n_812), .A2(n_924), .B1(n_925), .B2(n_926), .Y(n_923) );
INVx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OAI21xp5_ASAP7_75t_L g1196 ( .A1(n_816), .A2(n_1197), .B(n_1200), .Y(n_1196) );
INVx1_ASAP7_75t_L g1037 ( .A(n_817), .Y(n_1037) );
OAI22xp33_ASAP7_75t_L g1267 ( .A1(n_817), .A2(n_1023), .B1(n_1234), .B2(n_1243), .Y(n_1267) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_830), .A2(n_831), .B1(n_832), .B2(n_833), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1616 ( .A1(n_833), .A2(n_1617), .B1(n_1618), .B2(n_1619), .Y(n_1616) );
CKINVDCx11_ASAP7_75t_R g833 ( .A(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_837), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g894 ( .A(n_837), .B(n_895), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g1599 ( .A(n_837), .B(n_1600), .Y(n_1599) );
NOR2xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_843), .Y(n_839) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
NAND3xp33_ASAP7_75t_SL g843 ( .A(n_844), .B(n_846), .C(n_862), .Y(n_843) );
AOI33xp33_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_848), .A3(n_850), .B1(n_853), .B2(n_857), .B3(n_861), .Y(n_846) );
INVx2_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_864), .Y(n_863) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_867), .Y(n_974) );
XNOR2x1_ASAP7_75t_L g867 ( .A(n_868), .B(n_915), .Y(n_867) );
INVx1_ASAP7_75t_L g913 ( .A(n_869), .Y(n_913) );
NAND4xp25_ASAP7_75t_L g869 ( .A(n_870), .B(n_894), .C(n_896), .D(n_909), .Y(n_869) );
OAI21xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_883), .B(n_893), .Y(n_870) );
AOI21xp5_ASAP7_75t_L g875 ( .A1(n_876), .A2(n_878), .B(n_880), .Y(n_875) );
HB1xp67_ASAP7_75t_L g1528 ( .A(n_879), .Y(n_1528) );
INVx1_ASAP7_75t_L g1538 ( .A(n_879), .Y(n_1538) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_884) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_885), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_918) );
BUFx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
INVx2_ASAP7_75t_L g1125 ( .A(n_886), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1604 ( .A1(n_888), .A2(n_1124), .B1(n_1577), .B2(n_1579), .Y(n_1604) );
OAI31xp33_ASAP7_75t_L g1601 ( .A1(n_893), .A2(n_1602), .A3(n_1603), .B(n_1610), .Y(n_1601) );
INVx3_ASAP7_75t_L g1179 ( .A(n_899), .Y(n_1179) );
INVx2_ASAP7_75t_SL g902 ( .A(n_903), .Y(n_902) );
INVx1_ASAP7_75t_L g959 ( .A(n_903), .Y(n_959) );
INVx2_ASAP7_75t_L g1546 ( .A(n_903), .Y(n_1546) );
INVx1_ASAP7_75t_SL g972 ( .A(n_916), .Y(n_972) );
NAND4xp75_ASAP7_75t_L g916 ( .A(n_917), .B(n_937), .C(n_942), .D(n_968), .Y(n_916) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
OAI211xp5_ASAP7_75t_L g958 ( .A1(n_925), .A2(n_959), .B(n_960), .C(n_961), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g1022 ( .A1(n_926), .A2(n_1023), .B1(n_1024), .B2(n_1025), .Y(n_1022) );
BUFx3_ASAP7_75t_L g1133 ( .A(n_926), .Y(n_1133) );
INVx1_ASAP7_75t_L g1099 ( .A(n_928), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g1131 ( .A1(n_928), .A2(n_1132), .B1(n_1133), .B2(n_1134), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1140 ( .A1(n_928), .A2(n_1141), .B1(n_1142), .B2(n_1144), .Y(n_1140) );
BUFx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
BUFx2_ASAP7_75t_L g1027 ( .A(n_934), .Y(n_1027) );
NOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_941), .Y(n_937) );
INVx2_ASAP7_75t_SL g1151 ( .A(n_945), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_950), .B(n_958), .Y(n_949) );
OAI211xp5_ASAP7_75t_L g950 ( .A1(n_951), .A2(n_952), .B(n_954), .C(n_955), .Y(n_950) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx3_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
XNOR2xp5_ASAP7_75t_L g976 ( .A(n_977), .B(n_1172), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_978), .A2(n_979), .B1(n_1103), .B2(n_1104), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
AO22x1_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B1(n_1042), .B2(n_1043), .Y(n_979) );
INVx3_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g1040 ( .A(n_982), .Y(n_1040) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_983), .B(n_1009), .Y(n_982) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_996), .C(n_1004), .Y(n_984) );
INVx3_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_L g1184 ( .A(n_989), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g1031 ( .A1(n_992), .A2(n_1006), .B1(n_1027), .B2(n_1032), .Y(n_1031) );
INVx2_ASAP7_75t_SL g1000 ( .A(n_1001), .Y(n_1000) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1001), .Y(n_1229) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1035 ( .A1(n_1003), .A2(n_1005), .B1(n_1023), .B2(n_1036), .Y(n_1035) );
NOR3xp33_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1017), .C(n_1021), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1014), .Y(n_1010) );
OAI22xp33_ASAP7_75t_L g1085 ( .A1(n_1023), .A2(n_1086), .B1(n_1087), .B2(n_1088), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g1257 ( .A1(n_1023), .A2(n_1100), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_1027), .A2(n_1028), .B1(n_1029), .B2(n_1030), .Y(n_1026) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_1029), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1095 ( .A1(n_1029), .A2(n_1058), .B1(n_1072), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1036 ( .A(n_1037), .Y(n_1036) );
CKINVDCx8_ASAP7_75t_R g1038 ( .A(n_1039), .Y(n_1038) );
INVx2_ASAP7_75t_SL g1042 ( .A(n_1043), .Y(n_1042) );
XNOR2x1_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1102), .Y(n_1043) );
AND2x2_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1074), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_1046), .A2(n_1224), .B1(n_1245), .B2(n_1246), .Y(n_1223) );
NAND5xp2_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1056), .C(n_1059), .D(n_1063), .E(n_1071), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_1049), .A2(n_1057), .B1(n_1098), .B2(n_1100), .Y(n_1097) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1070 ( .A(n_1055), .Y(n_1070) );
OAI221xp5_ASAP7_75t_SL g1063 ( .A1(n_1064), .A2(n_1066), .B1(n_1067), .B2(n_1068), .C(n_1069), .Y(n_1063) );
INVx1_ASAP7_75t_L g1064 ( .A(n_1065), .Y(n_1064) );
NOR3xp33_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1080), .C(n_1084), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1078), .Y(n_1075) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1082), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1089 ( .A1(n_1090), .A2(n_1091), .B1(n_1092), .B2(n_1094), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g1260 ( .A1(n_1090), .A2(n_1261), .B1(n_1262), .B2(n_1263), .Y(n_1260) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_1096), .A2(n_1226), .B1(n_1244), .B2(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1098 ( .A(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1104 ( .A(n_1105), .Y(n_1104) );
INVx1_ASAP7_75t_L g1105 ( .A(n_1106), .Y(n_1105) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1107), .Y(n_1170) );
NOR3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1118), .C(n_1122), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1115), .Y(n_1110) );
OAI221xp5_ASAP7_75t_L g1161 ( .A1(n_1112), .A2(n_1117), .B1(n_1151), .B2(n_1162), .C(n_1164), .Y(n_1161) );
OAI22xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1126), .B1(n_1127), .B2(n_1130), .Y(n_1123) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_1124), .A2(n_1136), .B1(n_1137), .B2(n_1139), .Y(n_1135) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
INVx2_ASAP7_75t_SL g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_1130), .A2(n_1132), .B1(n_1149), .B2(n_1151), .C(n_1152), .Y(n_1148) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
OAI31xp33_ASAP7_75t_L g1145 ( .A1(n_1146), .A2(n_1155), .A3(n_1168), .B(n_1169), .Y(n_1145) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
HB1xp67_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
AO22x2_ASAP7_75t_L g1173 ( .A1(n_1174), .A2(n_1220), .B1(n_1221), .B2(n_1269), .Y(n_1173) );
INVxp67_ASAP7_75t_SL g1269 ( .A(n_1174), .Y(n_1269) );
INVxp67_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
NOR4xp75_ASAP7_75t_L g1176 ( .A(n_1177), .B(n_1192), .C(n_1213), .D(n_1218), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1188), .Y(n_1177) );
AOI33xp33_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1180), .A3(n_1182), .B1(n_1183), .B2(n_1185), .B3(n_1187), .Y(n_1178) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1187), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1210 ( .A(n_1211), .B(n_1212), .Y(n_1210) );
INVx2_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
XOR2x2_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1268), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1247), .Y(n_1222) );
NAND3xp33_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1232), .C(n_1242), .Y(n_1224) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
NOR3xp33_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1255), .C(n_1256), .Y(n_1247) );
NAND2xp5_ASAP7_75t_L g1248 ( .A(n_1249), .B(n_1252), .Y(n_1248) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1382 ( .A1(n_1268), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_1272), .A2(n_1510), .B1(n_1511), .B2(n_1562), .C(n_1565), .Y(n_1271) );
NOR2x1_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1450), .Y(n_1272) );
NAND4xp25_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1387), .C(n_1414), .D(n_1427), .Y(n_1273) );
A2O1A1Ixp33_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1300), .B(n_1330), .C(n_1376), .Y(n_1274) );
INVx1_ASAP7_75t_L g1420 ( .A(n_1275), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1426 ( .A(n_1275), .B(n_1364), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1275), .B(n_1334), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1504 ( .A(n_1275), .B(n_1438), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1296), .Y(n_1275) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1276), .Y(n_1356) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1276), .B(n_1297), .Y(n_1372) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1277), .B(n_1297), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1390 ( .A(n_1277), .B(n_1391), .Y(n_1390) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1290), .Y(n_1277) );
AND2x4_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1285), .Y(n_1279) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1326 ( .A(n_1281), .B(n_1286), .Y(n_1326) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1282), .B(n_1284), .Y(n_1281) );
HB1xp67_ASAP7_75t_L g1625 ( .A(n_1282), .Y(n_1625) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1284), .Y(n_1294) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1285), .B(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1286), .Y(n_1285) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1286), .B(n_1289), .Y(n_1329) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1292), .B(n_1293), .Y(n_1291) );
AND2x4_ASAP7_75t_L g1295 ( .A(n_1292), .B(n_1294), .Y(n_1295) );
AND2x4_ASAP7_75t_L g1307 ( .A(n_1292), .B(n_1293), .Y(n_1307) );
HB1xp67_ASAP7_75t_L g1626 ( .A(n_1293), .Y(n_1626) );
INVx1_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1295), .Y(n_1316) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1297), .Y(n_1333) );
INVxp67_ASAP7_75t_SL g1391 ( .A(n_1297), .Y(n_1391) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1297), .B(n_1334), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1299), .Y(n_1297) );
NOR2xp33_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1318), .Y(n_1300) );
OAI221xp5_ASAP7_75t_L g1500 ( .A1(n_1301), .A2(n_1501), .B1(n_1506), .B2(n_1507), .C(n_1508), .Y(n_1500) );
OR2x2_ASAP7_75t_L g1301 ( .A(n_1302), .B(n_1311), .Y(n_1301) );
INVx2_ASAP7_75t_L g1371 ( .A(n_1302), .Y(n_1371) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1302), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1303), .B(n_1308), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1303), .B(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1304), .Y(n_1344) );
AND2x2_ASAP7_75t_L g1362 ( .A(n_1304), .B(n_1308), .Y(n_1362) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1304), .B(n_1311), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1304), .B(n_1340), .Y(n_1403) );
BUFx6f_ASAP7_75t_L g1415 ( .A(n_1304), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1306), .Y(n_1304) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1307), .Y(n_1314) );
BUFx3_ASAP7_75t_L g1380 ( .A(n_1307), .Y(n_1380) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1308), .Y(n_1340) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1308), .Y(n_1354) );
INVx1_ASAP7_75t_L g1360 ( .A(n_1308), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1308), .B(n_1343), .Y(n_1406) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1308), .B(n_1320), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1310), .Y(n_1308) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1311), .B(n_1339), .Y(n_1338) );
CKINVDCx6p67_ASAP7_75t_R g1343 ( .A(n_1311), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1311), .B(n_1349), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1357 ( .A(n_1311), .B(n_1344), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1311), .B(n_1344), .Y(n_1407) );
NAND2xp5_ASAP7_75t_L g1462 ( .A(n_1311), .B(n_1353), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1506 ( .A(n_1311), .B(n_1378), .Y(n_1506) );
OR2x6_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1312), .B(n_1313), .Y(n_1368) );
OAI22xp5_ASAP7_75t_SL g1313 ( .A1(n_1314), .A2(n_1315), .B1(n_1316), .B2(n_1317), .Y(n_1313) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1316), .Y(n_1322) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1316), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1318), .B(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_1319), .B(n_1363), .Y(n_1395) );
NOR2xp33_ASAP7_75t_L g1502 ( .A(n_1319), .B(n_1503), .Y(n_1502) );
BUFx3_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_1320), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1359 ( .A(n_1320), .B(n_1360), .Y(n_1359) );
NOR2xp33_ASAP7_75t_L g1375 ( .A(n_1320), .B(n_1340), .Y(n_1375) );
BUFx2_ASAP7_75t_L g1423 ( .A(n_1320), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1320), .B(n_1334), .Y(n_1438) );
INVx2_ASAP7_75t_SL g1320 ( .A(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1321), .B(n_1340), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1321), .B(n_1364), .Y(n_1392) );
OAI22xp33_ASAP7_75t_L g1323 ( .A1(n_1324), .A2(n_1325), .B1(n_1327), .B2(n_1328), .Y(n_1323) );
BUFx3_ASAP7_75t_L g1383 ( .A(n_1325), .Y(n_1383) );
BUFx6f_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1328 ( .A(n_1329), .Y(n_1328) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1329), .Y(n_1386) );
OAI211xp5_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1337), .B(n_1341), .C(n_1370), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1334), .Y(n_1332) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1333), .B(n_1359), .Y(n_1358) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1333), .Y(n_1478) );
OR2x2_ASAP7_75t_L g1490 ( .A(n_1333), .B(n_1334), .Y(n_1490) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1334), .B(n_1346), .Y(n_1345) );
CKINVDCx5p33_ASAP7_75t_R g1364 ( .A(n_1334), .Y(n_1364) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_1334), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1429 ( .A(n_1334), .B(n_1355), .Y(n_1429) );
NOR2xp33_ASAP7_75t_L g1445 ( .A(n_1334), .B(n_1356), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1468 ( .A(n_1334), .B(n_1390), .Y(n_1468) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1334), .B(n_1356), .Y(n_1475) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1334), .B(n_1478), .Y(n_1477) );
AND2x4_ASAP7_75t_SL g1334 ( .A(n_1335), .B(n_1336), .Y(n_1334) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
AOI221xp5_ASAP7_75t_L g1463 ( .A1(n_1338), .A2(n_1390), .B1(n_1464), .B2(n_1465), .C(n_1466), .Y(n_1463) );
NAND3xp33_ASAP7_75t_L g1410 ( .A(n_1339), .B(n_1411), .C(n_1412), .Y(n_1410) );
AOI221xp5_ASAP7_75t_L g1491 ( .A1(n_1339), .A2(n_1354), .B1(n_1454), .B2(n_1492), .C(n_1495), .Y(n_1491) );
AOI211xp5_ASAP7_75t_L g1341 ( .A1(n_1342), .A2(n_1345), .B(n_1347), .C(n_1365), .Y(n_1341) );
AOI331xp33_ASAP7_75t_L g1414 ( .A1(n_1342), .A2(n_1376), .A3(n_1389), .B1(n_1415), .B2(n_1416), .B3(n_1421), .C1(n_1424), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1342 ( .A(n_1343), .B(n_1344), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1343), .B(n_1403), .Y(n_1402) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1343), .B(n_1377), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1397 ( .A(n_1344), .B(n_1377), .Y(n_1397) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1344), .Y(n_1440) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1345), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1509 ( .A(n_1345), .B(n_1422), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1363 ( .A(n_1346), .B(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1346), .Y(n_1369) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1346), .B(n_1375), .Y(n_1374) );
OAI321xp33_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1351), .A3(n_1355), .B1(n_1357), .B2(n_1358), .C(n_1361), .Y(n_1347) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1348), .Y(n_1411) );
INVxp67_ASAP7_75t_L g1349 ( .A(n_1350), .Y(n_1349) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1350), .B(n_1429), .Y(n_1428) );
NOR2xp33_ASAP7_75t_L g1457 ( .A(n_1350), .B(n_1458), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g1461 ( .A(n_1350), .Y(n_1461) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1350), .B(n_1372), .Y(n_1494) );
O2A1O1Ixp33_ASAP7_75t_SL g1404 ( .A1(n_1351), .A2(n_1376), .B(n_1405), .C(n_1407), .Y(n_1404) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1351), .B(n_1454), .Y(n_1453) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1352), .Y(n_1433) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1353), .B(n_1389), .Y(n_1388) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1353), .B(n_1437), .Y(n_1436) );
INVx3_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
NAND2xp5_ASAP7_75t_L g1431 ( .A(n_1354), .B(n_1393), .Y(n_1431) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
AOI222xp33_ASAP7_75t_L g1501 ( .A1(n_1356), .A2(n_1362), .B1(n_1415), .B2(n_1502), .C1(n_1504), .C2(n_1505), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1455 ( .A(n_1360), .B(n_1456), .Y(n_1455) );
OAI221xp5_ASAP7_75t_SL g1486 ( .A1(n_1360), .A2(n_1487), .B1(n_1489), .B2(n_1490), .C(n_1491), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1361 ( .A(n_1362), .B(n_1363), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_1362), .B(n_1423), .Y(n_1497) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1362), .Y(n_1503) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1364), .B(n_1390), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1435 ( .A(n_1364), .B(n_1372), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1364), .B(n_1457), .Y(n_1456) );
OR2x2_ASAP7_75t_L g1493 ( .A(n_1364), .B(n_1494), .Y(n_1493) );
NOR2xp33_ASAP7_75t_L g1495 ( .A(n_1364), .B(n_1496), .Y(n_1495) );
NOR3xp33_ASAP7_75t_L g1365 ( .A(n_1366), .B(n_1368), .C(n_1369), .Y(n_1365) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
A2O1A1Ixp33_ASAP7_75t_L g1370 ( .A1(n_1368), .A2(n_1371), .B(n_1372), .C(n_1373), .Y(n_1370) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1368), .B(n_1425), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1369), .B(n_1420), .Y(n_1419) );
OR2x2_ASAP7_75t_L g1469 ( .A(n_1369), .B(n_1470), .Y(n_1469) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1372), .B(n_1392), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1488 ( .A(n_1372), .B(n_1438), .Y(n_1488) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1375), .B(n_1426), .Y(n_1425) );
INVx3_ASAP7_75t_L g1484 ( .A(n_1376), .Y(n_1484) );
A2O1A1Ixp33_ASAP7_75t_L g1508 ( .A1(n_1376), .A2(n_1433), .B(n_1439), .C(n_1509), .Y(n_1508) );
INVx2_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1379), .B(n_1440), .Y(n_1439) );
CKINVDCx5p33_ASAP7_75t_R g1510 ( .A(n_1380), .Y(n_1510) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
AOI221xp5_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1393), .B1(n_1394), .B2(n_1396), .C(n_1398), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1392), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1390), .B(n_1438), .Y(n_1437) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1390), .Y(n_1458) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1392), .Y(n_1470) );
AOI21xp5_ASAP7_75t_L g1472 ( .A1(n_1393), .A2(n_1473), .B(n_1479), .Y(n_1472) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_L g1398 ( .A1(n_1399), .A2(n_1401), .B1(n_1404), .B2(n_1408), .C(n_1410), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1464 ( .A(n_1399), .B(n_1442), .Y(n_1464) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1403), .Y(n_1471) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1403), .B(n_1423), .Y(n_1489) );
CKINVDCx5p33_ASAP7_75t_R g1405 ( .A(n_1406), .Y(n_1405) );
AOI211xp5_ASAP7_75t_L g1451 ( .A1(n_1407), .A2(n_1452), .B(n_1455), .C(n_1459), .Y(n_1451) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1481 ( .A(n_1413), .B(n_1482), .Y(n_1481) );
NAND2xp5_ASAP7_75t_L g1480 ( .A(n_1415), .B(n_1481), .Y(n_1480) );
NOR2xp33_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1418), .Y(n_1416) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1419), .Y(n_1418) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1505 ( .A(n_1422), .B(n_1477), .Y(n_1505) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1423), .B(n_1440), .Y(n_1465) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1423), .B(n_1477), .Y(n_1476) );
AOI221xp5_ASAP7_75t_L g1427 ( .A1(n_1428), .A2(n_1430), .B1(n_1432), .B2(n_1439), .C(n_1441), .Y(n_1427) );
INVx1_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
OAI21xp33_ASAP7_75t_L g1432 ( .A1(n_1433), .A2(n_1434), .B(n_1436), .Y(n_1432) );
OAI21xp33_ASAP7_75t_L g1473 ( .A1(n_1433), .A2(n_1474), .B(n_1476), .Y(n_1473) );
AOI21xp33_ASAP7_75t_SL g1459 ( .A1(n_1434), .A2(n_1460), .B(n_1462), .Y(n_1459) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
AOI21xp5_ASAP7_75t_L g1441 ( .A1(n_1442), .A2(n_1443), .B(n_1446), .Y(n_1441) );
INVx1_ASAP7_75t_L g1443 ( .A(n_1444), .Y(n_1443) );
HB1xp67_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1448), .Y(n_1447) );
A2O1A1Ixp33_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1463), .B(n_1483), .C(n_1485), .Y(n_1450) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1454), .B(n_1461), .Y(n_1460) );
A2O1A1Ixp33_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1469), .B(n_1471), .C(n_1472), .Y(n_1466) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
NOR2xp33_ASAP7_75t_L g1487 ( .A(n_1468), .B(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
AOI21xp33_ASAP7_75t_SL g1485 ( .A1(n_1486), .A2(n_1498), .B(n_1500), .Y(n_1485) );
INVx2_ASAP7_75t_L g1492 ( .A(n_1493), .Y(n_1492) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1499), .Y(n_1498) );
INVxp67_ASAP7_75t_L g1507 ( .A(n_1505), .Y(n_1507) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1513), .Y(n_1561) );
BUFx2_ASAP7_75t_L g1513 ( .A(n_1514), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1539), .Y(n_1514) );
AND4x1_ASAP7_75t_L g1515 ( .A(n_1516), .B(n_1519), .C(n_1523), .D(n_1526), .Y(n_1515) );
OAI211xp5_ASAP7_75t_L g1545 ( .A1(n_1522), .A2(n_1546), .B(n_1547), .C(n_1548), .Y(n_1545) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1537 ( .A(n_1538), .Y(n_1537) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1562 ( .A(n_1563), .Y(n_1562) );
A2O1A1Ixp33_ASAP7_75t_L g1623 ( .A1(n_1564), .A2(n_1624), .B(n_1626), .C(n_1627), .Y(n_1623) );
BUFx2_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
HB1xp67_ASAP7_75t_L g1569 ( .A(n_1570), .Y(n_1569) );
AND4x1_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1599), .C(n_1601), .D(n_1620), .Y(n_1571) );
OAI33xp33_ASAP7_75t_L g1573 ( .A1(n_1574), .A2(n_1575), .A3(n_1580), .B1(n_1585), .B2(n_1592), .B3(n_1597), .Y(n_1573) );
OAI22xp33_ASAP7_75t_L g1575 ( .A1(n_1576), .A2(n_1577), .B1(n_1578), .B2(n_1579), .Y(n_1575) );
OAI22xp33_ASAP7_75t_L g1580 ( .A1(n_1581), .A2(n_1582), .B1(n_1583), .B2(n_1584), .Y(n_1580) );
OAI21xp33_ASAP7_75t_SL g1605 ( .A1(n_1584), .A2(n_1606), .B(n_1607), .Y(n_1605) );
OAI22xp5_ASAP7_75t_L g1585 ( .A1(n_1586), .A2(n_1587), .B1(n_1588), .B2(n_1591), .Y(n_1585) );
INVx2_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
OAI22xp5_ASAP7_75t_L g1592 ( .A1(n_1593), .A2(n_1594), .B1(n_1595), .B2(n_1596), .Y(n_1592) );
INVx2_ASAP7_75t_SL g1608 ( .A(n_1609), .Y(n_1608) );
NOR2xp33_ASAP7_75t_L g1620 ( .A(n_1621), .B(n_1622), .Y(n_1620) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
endmodule