module fake_jpeg_557_n_426 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_426);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_426;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx8_ASAP7_75t_L g184 ( 
.A(n_53),
.Y(n_184)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_55),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_6),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_58),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_5),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_5),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_60),
.B(n_74),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_24),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_67),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_21),
.B(n_8),
.C(n_12),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_91),
.Y(n_114)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_70),
.Y(n_177)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_72),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_25),
.B(n_9),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_75),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_76),
.Y(n_151)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_20),
.B(n_16),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_79),
.B(n_81),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_80),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_29),
.B(n_9),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_19),
.Y(n_82)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_82),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_83),
.Y(n_166)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_84),
.Y(n_155)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_19),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_85),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_37),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_86),
.B(n_90),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_87),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_88),
.Y(n_167)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_12),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_26),
.B(n_0),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_93),
.Y(n_171)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_29),
.B(n_0),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_0),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_107),
.Y(n_117)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_18),
.B(n_1),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_101),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

BUFx2_ASAP7_75t_SL g162 ( 
.A(n_100),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_27),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_103),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_43),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_41),
.B(n_1),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_42),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_113),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_112),
.B(n_1),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_42),
.B(n_47),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_L g115 ( 
.A1(n_63),
.A2(n_50),
.B1(n_34),
.B2(n_48),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_126),
.B1(n_172),
.B2(n_190),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_99),
.A2(n_47),
.B1(n_49),
.B2(n_44),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_91),
.B(n_44),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_129),
.B(n_132),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_111),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_56),
.A2(n_49),
.B1(n_50),
.B2(n_34),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_138),
.A2(n_142),
.B1(n_146),
.B2(n_152),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_53),
.A2(n_33),
.B1(n_37),
.B2(n_48),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_33),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_144),
.B(n_149),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_53),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_73),
.Y(n_149)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_45),
.CON(n_150),
.SN(n_150)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_150),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_100),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_78),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_153),
.A2(n_168),
.B1(n_176),
.B2(n_133),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_76),
.B(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_170),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_108),
.A2(n_36),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_159),
.A2(n_145),
.B1(n_187),
.B2(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_68),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_160),
.B(n_185),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_163),
.B(n_133),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_72),
.A2(n_2),
.B1(n_36),
.B2(n_102),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_107),
.B(n_87),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_104),
.A2(n_105),
.B1(n_59),
.B2(n_101),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_103),
.A2(n_85),
.B1(n_92),
.B2(n_88),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_87),
.B(n_93),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_179),
.B(n_180),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_84),
.B(n_77),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_82),
.B(n_64),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_181),
.B(n_188),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_66),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g186 ( 
.A1(n_70),
.A2(n_79),
.B(n_90),
.Y(n_186)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_186),
.B(n_146),
.CI(n_142),
.CON(n_225),
.SN(n_225)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_113),
.B(n_79),
.Y(n_188)
);

OAI22xp33_ASAP7_75t_L g190 ( 
.A1(n_63),
.A2(n_72),
.B1(n_68),
.B2(n_78),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g266 ( 
.A(n_191),
.Y(n_266)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_192),
.Y(n_255)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_193),
.A2(n_246),
.B1(n_216),
.B2(n_212),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_195),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_119),
.A2(n_172),
.B1(n_114),
.B2(n_135),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_196),
.A2(n_198),
.B(n_204),
.Y(n_290)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_198),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_127),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_199),
.B(n_210),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_120),
.B1(n_115),
.B2(n_116),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_200),
.A2(n_207),
.B1(n_217),
.B2(n_224),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_138),
.B1(n_152),
.B2(n_159),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_202),
.A2(n_194),
.B1(n_247),
.B2(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_203),
.Y(n_264)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_204),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_140),
.Y(n_206)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_143),
.A2(n_157),
.B1(n_183),
.B2(n_154),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_208),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_209),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_164),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_211),
.Y(n_260)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_166),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_215),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_119),
.A2(n_145),
.B1(n_124),
.B2(n_121),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_230),
.B1(n_237),
.B2(n_241),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_148),
.B1(n_154),
.B2(n_122),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_178),
.Y(n_218)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_218),
.Y(n_270)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_221),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_175),
.A2(n_182),
.B1(n_130),
.B2(n_141),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_225),
.B(n_229),
.Y(n_284)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_174),
.Y(n_227)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_227),
.Y(n_287)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_228),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_117),
.B(n_165),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_124),
.A2(n_137),
.B1(n_187),
.B2(n_118),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_165),
.Y(n_231)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_156),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_233),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_166),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_234),
.Y(n_296)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_161),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_235),
.Y(n_261)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_236),
.Y(n_275)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_173),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_238),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_148),
.A2(n_147),
.B1(n_131),
.B2(n_169),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_239),
.A2(n_248),
.B1(n_200),
.B2(n_217),
.Y(n_273)
);

INVx6_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_242),
.Y(n_265)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_249),
.Y(n_289)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_167),
.Y(n_245)
);

AO22x1_ASAP7_75t_SL g246 ( 
.A1(n_133),
.A2(n_119),
.B1(n_126),
.B2(n_99),
.Y(n_246)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_177),
.A2(n_119),
.B1(n_126),
.B2(n_114),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_247),
.B(n_253),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_177),
.A2(n_126),
.B1(n_114),
.B2(n_190),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_167),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_250),
.B(n_252),
.Y(n_299)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_182),
.B(n_175),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_254),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_283),
.B1(n_254),
.B2(n_268),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_246),
.C(n_233),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_271),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_222),
.C(n_223),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g326 ( 
.A1(n_273),
.A2(n_255),
.B1(n_291),
.B2(n_285),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_226),
.B(n_193),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_286),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_201),
.B(n_202),
.C(n_237),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_283),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_201),
.B(n_208),
.C(n_215),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_214),
.B(n_206),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_201),
.A2(n_207),
.B1(n_230),
.B2(n_205),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_288),
.A2(n_272),
.B1(n_265),
.B2(n_294),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_290),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_191),
.A2(n_211),
.B(n_252),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_293),
.A2(n_240),
.B(n_257),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_195),
.B(n_245),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_255),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_300),
.A2(n_320),
.B(n_308),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_284),
.A3(n_263),
.B1(n_282),
.B2(n_262),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_305),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_274),
.A2(n_254),
.B1(n_289),
.B2(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_311),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_254),
.A2(n_288),
.B1(n_290),
.B2(n_286),
.Y(n_304)
);

AO21x2_ASAP7_75t_L g351 ( 
.A1(n_307),
.A2(n_320),
.B(n_327),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_266),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_271),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_265),
.A2(n_296),
.B1(n_299),
.B2(n_293),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_275),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_313),
.B(n_323),
.Y(n_356)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_299),
.Y(n_314)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_266),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_258),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_287),
.A2(n_264),
.B1(n_277),
.B2(n_260),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_317),
.A2(n_326),
.B1(n_320),
.B2(n_315),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_264),
.B(n_292),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_261),
.A2(n_256),
.B1(n_295),
.B2(n_277),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_319),
.A2(n_314),
.B1(n_330),
.B2(n_311),
.Y(n_337)
);

AOI22x1_ASAP7_75t_L g320 ( 
.A1(n_267),
.A2(n_281),
.B1(n_259),
.B2(n_258),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_292),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_332),
.Y(n_349)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_270),
.Y(n_322)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_322),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_269),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_276),
.A2(n_281),
.B(n_278),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_324),
.A2(n_318),
.B(n_317),
.Y(n_354)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_267),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_327),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_291),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_328),
.B(n_329),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_199),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_299),
.Y(n_330)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_330),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_274),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_274),
.B(n_286),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_309),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_310),
.C(n_305),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_334),
.B(n_348),
.C(n_322),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_313),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_337),
.B(n_354),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_323),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_340),
.B(n_350),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_312),
.A2(n_307),
.B1(n_306),
.B2(n_303),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_341),
.A2(n_351),
.B1(n_349),
.B2(n_336),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_302),
.B1(n_306),
.B2(n_331),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_342),
.A2(n_300),
.B1(n_320),
.B2(n_316),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_325),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_345),
.B(n_352),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_346),
.A2(n_355),
.B1(n_316),
.B2(n_319),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_310),
.B(n_301),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_329),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_356),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_366),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_359),
.B(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_335),
.B(n_328),
.Y(n_361)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_361),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_348),
.B(n_321),
.C(n_324),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_334),
.C(n_340),
.Y(n_380)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_365),
.Y(n_377)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_371),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_368),
.B(n_370),
.Y(n_379)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_373),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_338),
.Y(n_373)
);

AND2x6_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_340),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_378),
.A2(n_336),
.B1(n_351),
.B2(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_380),
.B(n_384),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_361),
.Y(n_381)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_359),
.B(n_362),
.C(n_341),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_382),
.B(n_342),
.C(n_358),
.Y(n_387)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_357),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_383),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_392),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_380),
.B(n_364),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_358),
.B(n_371),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_391),
.A2(n_393),
.B(n_394),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_382),
.B(n_369),
.C(n_373),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_367),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_384),
.B(n_352),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_368),
.B(n_365),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_376),
.Y(n_399)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_386),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_401),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_376),
.Y(n_401)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_403),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_397),
.B(n_363),
.C(n_346),
.Y(n_404)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_404),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_389),
.B(n_344),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_406),
.B(n_389),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_404),
.A2(n_396),
.B(n_391),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_408),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_410),
.B(n_411),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_401),
.B(n_390),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_412),
.B(n_400),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_415),
.C(n_388),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_412),
.B(n_402),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_416),
.A2(n_409),
.B(n_408),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_417),
.A2(n_418),
.B1(n_419),
.B2(n_405),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_413),
.A2(n_387),
.B(n_407),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_420),
.B(n_421),
.C(n_385),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_417),
.A2(n_385),
.B1(n_399),
.B2(n_379),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_421),
.C(n_395),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_363),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_424),
.B(n_350),
.C(n_377),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_425),
.B(n_356),
.Y(n_426)
);


endmodule