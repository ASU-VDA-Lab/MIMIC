module fake_jpeg_9924_n_45 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_45);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_45;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_0),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.Y(n_37)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_0),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_12),
.B1(n_17),
.B2(n_16),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_2),
.Y(n_29)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_2),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_18),
.B(n_3),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_22),
.B1(n_4),
.B2(n_3),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_30),
.A2(n_4),
.B1(n_20),
.B2(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_36),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_40),
.B(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_41),
.B(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_42),
.B(n_38),
.Y(n_43)
);

INVxp33_ASAP7_75t_SL g44 ( 
.A(n_43),
.Y(n_44)
);

AOI21x1_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_39),
.B(n_32),
.Y(n_45)
);


endmodule