module real_jpeg_6270_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_28),
.B2(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_1),
.A2(n_28),
.B1(n_135),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_1),
.A2(n_28),
.B1(n_255),
.B2(n_258),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_1),
.A2(n_28),
.B1(n_177),
.B2(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_2),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_2),
.A2(n_54),
.B1(n_64),
.B2(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_2),
.A2(n_64),
.B1(n_86),
.B2(n_270),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_3),
.Y(n_85)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_3),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_4),
.A2(n_57),
.B1(n_262),
.B2(n_264),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_4),
.A2(n_57),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_5),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_5),
.Y(n_164)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_7),
.A2(n_125),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_7),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_7),
.A2(n_128),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_7),
.A2(n_65),
.B1(n_128),
.B2(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_7),
.A2(n_128),
.B1(n_293),
.B2(n_295),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_8),
.Y(n_162)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_8),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_9),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_9),
.A2(n_65),
.B1(n_158),
.B2(n_212),
.Y(n_211)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_10),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_12),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_12),
.Y(n_105)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_12),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_12),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_12),
.Y(n_203)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_13),
.Y(n_73)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_13),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_14),
.A2(n_95),
.B1(n_173),
.B2(n_176),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_15),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_15),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_15),
.B(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_15),
.B(n_230),
.C(n_234),
.Y(n_229)
);

OAI22xp33_ASAP7_75t_L g239 ( 
.A1(n_15),
.A2(n_240),
.B1(n_241),
.B2(n_244),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_15),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_15),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_15),
.A2(n_145),
.B1(n_292),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_217),
.B1(n_218),
.B2(n_362),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_18),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_215),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_189),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_20),
.B(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_131),
.C(n_168),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_21),
.B(n_360),
.Y(n_359)
);

BUFx24_ASAP7_75t_SL g364 ( 
.A(n_21),
.Y(n_364)
);

FAx1_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_60),
.CI(n_98),
.CON(n_21),
.SN(n_21)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_22),
.B(n_60),
.C(n_98),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_34),
.B2(n_52),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_23),
.A2(n_32),
.B1(n_34),
.B2(n_183),
.Y(n_182)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_24),
.Y(n_334)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_26),
.Y(n_322)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_27),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_27),
.Y(n_134)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_27),
.Y(n_188)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_33),
.A2(n_53),
.B(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_33),
.A2(n_184),
.B1(n_252),
.B2(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_46),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_34),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_34),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_36),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_37),
.Y(n_244)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_37),
.Y(n_257)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_37),
.Y(n_258)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_37),
.Y(n_329)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_40),
.Y(n_325)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx5_ASAP7_75t_L g247 ( 
.A(n_41),
.Y(n_247)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_42),
.Y(n_213)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_42),
.Y(n_228)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_42),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_42),
.Y(n_339)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_48),
.Y(n_196)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_51),
.Y(n_319)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_66),
.B(n_88),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_61),
.B(n_90),
.Y(n_353)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_66),
.A2(n_90),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_66),
.A2(n_351),
.B(n_352),
.Y(n_350)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_67),
.A2(n_89),
.B1(n_239),
.B2(n_245),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_67),
.A2(n_89),
.B1(n_245),
.B2(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_67),
.A2(n_89),
.B1(n_254),
.B2(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_79),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_71),
.B1(n_74),
.B2(n_77),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_76),
.Y(n_233)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_85),
.Y(n_266)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_85),
.Y(n_308)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_90),
.B(n_240),
.Y(n_290)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_91),
.Y(n_210)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_97),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_106),
.B1(n_123),
.B2(n_130),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_100),
.A2(n_108),
.B1(n_110),
.B2(n_112),
.Y(n_107)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp33_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_106),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_124),
.A2(n_181),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_130),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_131),
.B(n_168),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_144),
.Y(n_191)
);

OAI32xp33_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_135),
.A3(n_137),
.B1(n_139),
.B2(n_143),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_154),
.B1(n_161),
.B2(n_163),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_163),
.B(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_145),
.A2(n_261),
.B(n_267),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_145),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_145),
.A2(n_279),
.B1(n_292),
.B2(n_296),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_145),
.A2(n_207),
.B(n_269),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_146),
.Y(n_280)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_148),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_150),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_155),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_151),
.B(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_SL g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_153),
.Y(n_304)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_179),
.C(n_182),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_169),
.A2(n_170),
.B1(n_179),
.B2(n_180),
.Y(n_346)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_175),
.Y(n_272)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_182),
.B(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI32xp33_ASAP7_75t_L g316 ( 
.A1(n_187),
.A2(n_317),
.A3(n_319),
.B1(n_320),
.B2(n_323),
.Y(n_316)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_204),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_214),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_209),
.Y(n_205)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_357),
.B(n_361),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_341),
.B(n_356),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_312),
.B(n_340),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_275),
.B(n_311),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_248),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_223),
.B(n_248),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_238),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_224),
.B(n_238),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_240),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_240),
.B(n_321),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_SL g333 ( 
.A1(n_240),
.A2(n_320),
.B(n_334),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_260),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_259),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_259),
.C(n_260),
.Y(n_313)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_253),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx8_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_288),
.B(n_310),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_287),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_287),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_298),
.B(n_309),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_290),
.B(n_291),
.Y(n_309)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_313),
.B(n_314),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_331),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_332),
.C(n_335),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_330),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_316),
.B(n_330),
.Y(n_349)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_326),
.Y(n_323)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_328),
.Y(n_337)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_342),
.B(n_343),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_345),
.B1(n_347),
.B2(n_348),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_350),
.C(n_354),
.Y(n_358)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_349),
.A2(n_350),
.B1(n_354),
.B2(n_355),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_359),
.Y(n_361)
);


endmodule