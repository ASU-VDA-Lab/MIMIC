module real_jpeg_21219_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_110;
wire n_61;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_97;
wire n_75;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_0),
.A2(n_72),
.B1(n_78),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_0),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_150),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_1),
.Y(n_148)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_14),
.B(n_34),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_148),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_1),
.A2(n_59),
.B1(n_203),
.B2(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_1),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_1),
.B(n_46),
.Y(n_230)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_1),
.A2(n_46),
.B(n_230),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_2),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_3),
.A2(n_72),
.B1(n_78),
.B2(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_3),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_128),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_128),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_3),
.A2(n_27),
.B1(n_30),
.B2(n_128),
.Y(n_221)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_4),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_4),
.A2(n_87),
.B(n_157),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_4),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_5),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_7),
.A2(n_29),
.B1(n_72),
.B2(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_7),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_8),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_38),
.B1(n_72),
.B2(n_78),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_8),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_9),
.A2(n_46),
.B1(n_47),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_53),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_53),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_11),
.A2(n_72),
.B1(n_78),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_11),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_96),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_96),
.Y(n_237)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_71),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_30),
.B(n_32),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_131),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_130),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_105),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_20),
.B(n_105),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_104),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_55),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_54),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_24),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_25),
.A2(n_40),
.B(n_237),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_26),
.Y(n_141)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_27),
.A2(n_35),
.B(n_148),
.C(n_195),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_27),
.B(n_44),
.Y(n_231)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_30),
.A2(n_45),
.A3(n_47),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_31),
.B(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_32),
.A2(n_40),
.B1(n_64),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_32),
.A2(n_36),
.B(n_92),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_32),
.A2(n_40),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_32),
.B(n_148),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_32),
.A2(n_40),
.B1(n_199),
.B2(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_32),
.A2(n_40),
.B1(n_221),
.B2(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_33),
.B(n_209),
.Y(n_208)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_64),
.B(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_40),
.A2(n_65),
.B(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_42)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_43),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_43),
.A2(n_49),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_43),
.A2(n_49),
.B1(n_144),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_43),
.A2(n_49),
.B1(n_175),
.B2(n_234),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_46),
.B(n_71),
.Y(n_154)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_47),
.A2(n_74),
.B1(n_147),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_50),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_49),
.B(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_49),
.B(n_123),
.Y(n_166)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_66),
.B2(n_67),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_63),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_68),
.B1(n_81),
.B2(n_82),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_58),
.A2(n_63),
.B1(n_82),
.B2(n_110),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B(n_61),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_59),
.A2(n_118),
.B(n_119),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_59),
.A2(n_118),
.B1(n_156),
.B2(n_158),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_59),
.A2(n_189),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_59),
.A2(n_89),
.B(n_191),
.Y(n_222)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_88),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_60),
.B(n_148),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_62),
.A2(n_120),
.B(n_187),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_76),
.B(n_79),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_95),
.B(n_97),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_69),
.A2(n_95),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_69),
.A2(n_127),
.B1(n_129),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_75),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_72),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g147 ( 
.A(n_72),
.B(n_148),
.CON(n_147),
.SN(n_147)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_83),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.C(n_98),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_91),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_85),
.B(n_91),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_89),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_101),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_101),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.C(n_111),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_106),
.A2(n_107),
.B1(n_109),
.B2(n_280),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_109),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_111),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_121),
.C(n_125),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_112),
.A2(n_113),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_117),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_121),
.A2(n_125),
.B1(n_126),
.B2(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_121),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_148),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_276),
.B(n_281),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_179),
.B(n_261),
.C(n_275),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_168),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_134),
.B(n_168),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_151),
.B2(n_167),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_137),
.B(n_138),
.C(n_167),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_146),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_139),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_170),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_149),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_152),
.B(n_160),
.C(n_164),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_155),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_164),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_171),
.C(n_173),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_169),
.B(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_171),
.A2(n_172),
.B1(n_173),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_174),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_176),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_260),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_254),
.B(n_259),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_242),
.B(n_253),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_224),
.B(n_241),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_212),
.B(n_223),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_200),
.B(n_211),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_186),
.B(n_192),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_206),
.B(n_210),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_205),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_213),
.B(n_214),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_220),
.C(n_222),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_232),
.B1(n_239),
.B2(n_240),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_232),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_235),
.B1(n_236),
.B2(n_238),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_251),
.C(n_252),
.Y(n_255)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_256),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_273),
.B2(n_274),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_269),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule