module fake_jpeg_13751_n_524 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_524);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_524;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g115 ( 
.A(n_61),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_62),
.Y(n_111)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_66),
.Y(n_104)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_69),
.B(n_76),
.Y(n_113)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_75),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_0),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_84),
.Y(n_148)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_32),
.B(n_2),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_96),
.B(n_99),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_97),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_100),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_30),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_21),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_40),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_31),
.B1(n_36),
.B2(n_40),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_109),
.A2(n_121),
.B1(n_130),
.B2(n_138),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_120),
.B(n_81),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_95),
.A2(n_31),
.B1(n_40),
.B2(n_28),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_79),
.B(n_39),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_37),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_54),
.A2(n_31),
.B1(n_40),
.B2(n_28),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_19),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_134),
.B(n_145),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_58),
.A2(n_30),
.B1(n_25),
.B2(n_49),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_19),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_59),
.A2(n_45),
.B1(n_50),
.B2(n_18),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_146),
.A2(n_147),
.B1(n_153),
.B2(n_34),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_61),
.A2(n_70),
.B1(n_99),
.B2(n_68),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_101),
.A2(n_45),
.B1(n_50),
.B2(n_18),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_81),
.B(n_47),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_154),
.B(n_53),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_109),
.A2(n_98),
.B1(n_62),
.B2(n_71),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_159),
.A2(n_166),
.B1(n_185),
.B2(n_158),
.Y(n_234)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_160),
.Y(n_240)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_122),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_162),
.Y(n_217)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_167),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_164),
.B(n_199),
.Y(n_253)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_141),
.A2(n_86),
.B1(n_65),
.B2(n_92),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_113),
.B(n_47),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_169),
.B(n_170),
.Y(n_216)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_173),
.Y(n_225)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_172),
.Y(n_222)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_174),
.Y(n_236)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_135),
.Y(n_176)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_177),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_91),
.B1(n_89),
.B2(n_66),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_178),
.A2(n_206),
.B1(n_147),
.B2(n_49),
.Y(n_214)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_105),
.B(n_35),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_180),
.B(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_126),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_94),
.B1(n_73),
.B2(n_52),
.Y(n_185)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_107),
.Y(n_186)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_187),
.A2(n_190),
.B1(n_209),
.B2(n_136),
.Y(n_230)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_123),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

OA22x2_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_85),
.B1(n_72),
.B2(n_82),
.Y(n_190)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_191),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_129),
.Y(n_192)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_106),
.B(n_34),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_193),
.B(n_195),
.Y(n_252)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_196),
.B(n_198),
.Y(n_259)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_110),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_118),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_116),
.B(n_35),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_201),
.B(n_204),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_202),
.A2(n_207),
.B1(n_212),
.B2(n_213),
.Y(n_251)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_137),
.B(n_44),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_144),
.A2(n_51),
.B1(n_22),
.B2(n_41),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_104),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_144),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_208),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g209 ( 
.A1(n_149),
.A2(n_87),
.B1(n_42),
.B2(n_41),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_132),
.B(n_80),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_210),
.Y(n_255)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_158),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_214),
.A2(n_20),
.B1(n_4),
.B2(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_162),
.B(n_39),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_244),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_230),
.A2(n_245),
.B1(n_20),
.B2(n_4),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_115),
.B(n_136),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_231),
.A2(n_237),
.B(n_207),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_194),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_118),
.B(n_125),
.Y(n_237)
);

AOI32xp33_ASAP7_75t_L g238 ( 
.A1(n_197),
.A2(n_53),
.A3(n_143),
.B1(n_102),
.B2(n_37),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_238),
.B(n_258),
.C(n_26),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_165),
.B(n_155),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_159),
.A2(n_108),
.B1(n_149),
.B2(n_155),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_209),
.B(n_108),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_246),
.B(n_260),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_178),
.A2(n_139),
.B1(n_111),
.B2(n_150),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_256),
.B1(n_261),
.B2(n_160),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_182),
.A2(n_206),
.B1(n_139),
.B2(n_111),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_209),
.A3(n_190),
.B1(n_189),
.B2(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_188),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_190),
.A2(n_41),
.B1(n_25),
.B2(n_49),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_215),
.B(n_44),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_262),
.B(n_264),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_263),
.A2(n_278),
.B1(n_298),
.B2(n_235),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_215),
.B(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_265),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_260),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_266),
.B(n_285),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_225),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_267),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_200),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_268),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_213),
.B(n_22),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_270),
.A2(n_279),
.B(n_223),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_272),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_256),
.A2(n_214),
.B1(n_249),
.B2(n_230),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_273),
.A2(n_281),
.B1(n_286),
.B2(n_293),
.Y(n_330)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_228),
.B(n_211),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_275),
.B(n_294),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_234),
.A2(n_161),
.B1(n_202),
.B2(n_192),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_276),
.A2(n_287),
.B1(n_288),
.B2(n_295),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_277),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_258),
.A2(n_177),
.B(n_175),
.Y(n_279)
);

XOR2x1_ASAP7_75t_L g323 ( 
.A(n_280),
.B(n_302),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_217),
.A2(n_131),
.B1(n_97),
.B2(n_176),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_221),
.Y(n_282)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_241),
.Y(n_284)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_284),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_26),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_217),
.A2(n_42),
.B1(n_26),
.B2(n_25),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_228),
.A2(n_42),
.B1(n_22),
.B2(n_20),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_255),
.B(n_20),
.C(n_4),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_297),
.C(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_221),
.Y(n_290)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_290),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_216),
.B(n_2),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_292),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_225),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_239),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_238),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_222),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_296),
.B(n_299),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_233),
.B(n_219),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_304),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g298 ( 
.A1(n_255),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_222),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_233),
.B(n_17),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_301),
.Y(n_324)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_236),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_252),
.B(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_241),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_303),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_259),
.B(n_5),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_231),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_305),
.Y(n_321)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_232),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_307),
.B(n_341),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_310),
.Y(n_368)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_283),
.A2(n_253),
.B(n_254),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_313),
.A2(n_281),
.B(n_287),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_283),
.A2(n_250),
.B1(n_232),
.B2(n_226),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_317),
.B1(n_318),
.B2(n_320),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_273),
.A2(n_251),
.B1(n_250),
.B2(n_239),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_315),
.A2(n_332),
.B1(n_333),
.B2(n_336),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_232),
.B1(n_240),
.B2(n_218),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_240),
.B1(n_218),
.B2(n_243),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_288),
.A2(n_276),
.B1(n_265),
.B2(n_266),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_248),
.C(n_243),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_269),
.C(n_289),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_279),
.A2(n_263),
.B1(n_280),
.B2(n_305),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_271),
.A2(n_224),
.B1(n_240),
.B2(n_257),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_271),
.A2(n_224),
.B1(n_248),
.B2(n_229),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_270),
.A2(n_229),
.B1(n_235),
.B2(n_241),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_338),
.A2(n_330),
.B1(n_333),
.B2(n_336),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_339),
.A2(n_343),
.B1(n_285),
.B2(n_292),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_275),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_295),
.A2(n_272),
.B1(n_294),
.B2(n_267),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_286),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_341),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_369),
.C(n_370),
.Y(n_412)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_316),
.Y(n_350)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_350),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_315),
.A2(n_306),
.B1(n_303),
.B2(n_284),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_351),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_316),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_356),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_322),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_353),
.B(n_362),
.Y(n_387)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_354),
.Y(n_392)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_317),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_365),
.B1(n_371),
.B2(n_376),
.Y(n_403)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_311),
.B(n_264),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_359),
.B(n_360),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_300),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_361),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_337),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_311),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_363),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_364),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_320),
.A2(n_262),
.B1(n_299),
.B2(n_296),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_312),
.B(n_301),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_366),
.B(n_381),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_367),
.A2(n_380),
.B1(n_326),
.B2(n_344),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_323),
.B(n_282),
.C(n_277),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_290),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_308),
.A2(n_274),
.B1(n_220),
.B2(n_236),
.Y(n_371)
);

XOR2x2_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_227),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_375),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_319),
.B(n_220),
.Y(n_373)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_338),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_379),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_SL g375 ( 
.A(n_323),
.B(n_7),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_308),
.A2(n_319),
.B1(n_310),
.B2(n_343),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_324),
.B(n_242),
.Y(n_377)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

NAND2x1p5_ASAP7_75t_L g378 ( 
.A(n_321),
.B(n_242),
.Y(n_378)
);

OA22x2_ASAP7_75t_L g406 ( 
.A1(n_378),
.A2(n_325),
.B1(n_340),
.B2(n_328),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_314),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_332),
.A2(n_227),
.B1(n_8),
.B2(n_9),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_345),
.A2(n_7),
.B(n_8),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_366),
.B(n_329),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_368),
.A2(n_318),
.B(n_313),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_406),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_307),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_389),
.B(n_394),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_373),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g432 ( 
.A1(n_391),
.A2(n_396),
.B1(n_399),
.B2(n_400),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_313),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_313),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_395),
.B(n_405),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_359),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_377),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_376),
.A2(n_330),
.B1(n_331),
.B2(n_321),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_404),
.A2(n_408),
.B1(n_355),
.B2(n_352),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_358),
.B(n_326),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_406),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_325),
.B1(n_324),
.B2(n_328),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_354),
.Y(n_409)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_402),
.Y(n_413)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_413),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_347),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_414),
.B(n_421),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_312),
.B1(n_367),
.B2(n_355),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_416),
.A2(n_418),
.B1(n_419),
.B2(n_429),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_388),
.A2(n_379),
.B1(n_348),
.B2(n_350),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_368),
.C(n_378),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_420),
.B(n_433),
.C(n_401),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_375),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_392),
.Y(n_422)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_424),
.B(n_426),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_365),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_408),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_387),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_387),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_427),
.B(n_428),
.Y(n_449)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_390),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_388),
.A2(n_356),
.B1(n_371),
.B2(n_363),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_406),
.Y(n_430)
);

A2O1A1Ixp33_ASAP7_75t_SL g456 ( 
.A1(n_430),
.A2(n_356),
.B(n_364),
.C(n_397),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_394),
.C(n_386),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_435),
.Y(n_459)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_393),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_407),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_437),
.A2(n_353),
.B1(n_362),
.B2(n_349),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_386),
.Y(n_439)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_439),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_436),
.B(n_404),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_440),
.B(n_452),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_444),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_411),
.C(n_378),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_447),
.B(n_450),
.Y(n_460)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_438),
.B(n_406),
.C(n_403),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_438),
.B(n_415),
.C(n_433),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_453),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_436),
.B(n_403),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_393),
.C(n_400),
.Y(n_453)
);

FAx1_ASAP7_75t_SL g454 ( 
.A(n_432),
.B(n_360),
.CI(n_342),
.CON(n_454),
.SN(n_454)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_418),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_419),
.B(n_380),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_429),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_456),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_446),
.A2(n_413),
.B(n_424),
.Y(n_461)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_461),
.Y(n_485)
);

OAI221xp5_ASAP7_75t_L g462 ( 
.A1(n_459),
.A2(n_342),
.B1(n_435),
.B2(n_430),
.C(n_431),
.Y(n_462)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_462),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_464),
.A2(n_441),
.B1(n_454),
.B2(n_452),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_327),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_431),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_469),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_442),
.B(n_423),
.C(n_421),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_453),
.B(n_397),
.C(n_410),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_471),
.B(n_475),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_384),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_473),
.B(n_381),
.Y(n_488)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_457),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_461),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_477),
.B(n_482),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_466),
.A2(n_458),
.B1(n_455),
.B2(n_450),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_478),
.A2(n_479),
.B1(n_470),
.B2(n_471),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_474),
.A2(n_417),
.B1(n_447),
.B2(n_353),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_335),
.B1(n_346),
.B2(n_12),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_443),
.C(n_456),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_456),
.C(n_410),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_484),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_486),
.B(n_489),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_465),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_469),
.B(n_340),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_456),
.C(n_346),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_465),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_491),
.B(n_7),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g493 ( 
.A(n_480),
.B(n_467),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_493),
.B(n_500),
.Y(n_504)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_495),
.Y(n_506)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_496),
.Y(n_511)
);

AOI21xp33_ASAP7_75t_L g498 ( 
.A1(n_483),
.A2(n_468),
.B(n_473),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_498),
.B(n_499),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_485),
.A2(n_335),
.B1(n_10),
.B2(n_12),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_501),
.B(n_502),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g502 ( 
.A(n_487),
.B(n_16),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_503),
.B(n_491),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_482),
.C(n_484),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_497),
.C(n_500),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_509),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_492),
.B(n_490),
.Y(n_510)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_510),
.A2(n_499),
.B(n_503),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_508),
.Y(n_517)
);

AOI21x1_ASAP7_75t_SL g518 ( 
.A1(n_513),
.A2(n_515),
.B(n_507),
.Y(n_518)
);

AOI21x1_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_501),
.B(n_12),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_514),
.B(n_511),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_516),
.B(n_517),
.C(n_518),
.Y(n_519)
);

NAND3xp33_ASAP7_75t_L g520 ( 
.A(n_517),
.B(n_506),
.C(n_504),
.Y(n_520)
);

A2O1A1O1Ixp25_ASAP7_75t_L g521 ( 
.A1(n_520),
.A2(n_509),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_519),
.B1(n_13),
.B2(n_14),
.Y(n_522)
);

AO21x2_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_16),
.B(n_10),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_15),
.B(n_16),
.Y(n_524)
);


endmodule