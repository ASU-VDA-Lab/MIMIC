module fake_netlist_1_8455_n_814 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_814);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_814;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_808;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_802;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_223;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_33), .Y(n_103) );
INVx2_ASAP7_75t_SL g104 ( .A(n_22), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_58), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_25), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_19), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_81), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_17), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_43), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_68), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_41), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_36), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_88), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_8), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_14), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_39), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_8), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_69), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_53), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_51), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_36), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_95), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_17), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_31), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_57), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_100), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_101), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_60), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_34), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_74), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_92), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_31), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_18), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_25), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_22), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_70), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_2), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_10), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_35), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_63), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_44), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_65), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_111), .B(n_0), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_107), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_111), .B(n_0), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_130), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_104), .B(n_1), .Y(n_151) );
INVxp67_ASAP7_75t_L g152 ( .A(n_104), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_104), .B(n_1), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_130), .B(n_2), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_109), .B(n_3), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_130), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_107), .B(n_3), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_128), .B(n_4), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_128), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
AND2x4_ASAP7_75t_L g161 ( .A(n_113), .B(n_4), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_133), .B(n_5), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_133), .B(n_5), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_146), .Y(n_164) );
BUFx12f_ASAP7_75t_L g165 ( .A(n_105), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_113), .B(n_6), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_123), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_138), .B(n_6), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_123), .Y(n_169) );
AO22x2_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_146), .B1(n_125), .B2(n_126), .Y(n_170) );
INVx11_ASAP7_75t_L g171 ( .A(n_165), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_169), .Y(n_172) );
AO22x2_ASAP7_75t_L g173 ( .A1(n_151), .A2(n_134), .B1(n_132), .B2(n_126), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_169), .Y(n_174) );
OA22x2_ASAP7_75t_L g175 ( .A1(n_148), .A2(n_138), .B1(n_139), .B2(n_143), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
NOR2x1p5_ASAP7_75t_L g177 ( .A(n_147), .B(n_139), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_151), .A2(n_112), .B1(n_122), .B2(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_169), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_148), .B(n_141), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_147), .B(n_103), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_169), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_169), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_148), .B(n_141), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_159), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_159), .B(n_142), .Y(n_186) );
AND2x2_ASAP7_75t_L g187 ( .A(n_159), .B(n_142), .Y(n_187) );
INVxp67_ASAP7_75t_SL g188 ( .A(n_147), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_169), .Y(n_189) );
AO22x2_ASAP7_75t_L g190 ( .A1(n_151), .A2(n_125), .B1(n_132), .B2(n_134), .Y(n_190) );
AO22x2_ASAP7_75t_L g191 ( .A1(n_151), .A2(n_143), .B1(n_116), .B2(n_115), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_169), .Y(n_192) );
OAI22xp33_ASAP7_75t_L g193 ( .A1(n_149), .A2(n_120), .B1(n_106), .B2(n_119), .Y(n_193) );
XNOR2xp5_ASAP7_75t_L g194 ( .A(n_149), .B(n_145), .Y(n_194) );
OAI22xp33_ASAP7_75t_L g195 ( .A1(n_149), .A2(n_110), .B1(n_114), .B2(n_137), .Y(n_195) );
OAI22xp33_ASAP7_75t_SL g196 ( .A1(n_157), .A2(n_124), .B1(n_136), .B2(n_117), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_152), .B(n_108), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_151), .A2(n_154), .B1(n_166), .B2(n_161), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_153), .B(n_118), .Y(n_199) );
NOR2xp33_ASAP7_75t_R g200 ( .A(n_165), .B(n_121), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_169), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_151), .A2(n_127), .B1(n_116), .B2(n_115), .Y(n_202) );
BUFx2_ASAP7_75t_L g203 ( .A(n_165), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_169), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_152), .B(n_129), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_169), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_153), .B(n_135), .Y(n_207) );
AO22x2_ASAP7_75t_L g208 ( .A1(n_151), .A2(n_7), .B1(n_9), .B2(n_10), .Y(n_208) );
AO22x2_ASAP7_75t_L g209 ( .A1(n_166), .A2(n_7), .B1(n_9), .B2(n_11), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_152), .B(n_140), .Y(n_210) );
OA22x2_ASAP7_75t_L g211 ( .A1(n_154), .A2(n_144), .B1(n_12), .B2(n_13), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_154), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_154), .Y(n_214) );
AND2x2_ASAP7_75t_L g215 ( .A(n_153), .B(n_14), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_154), .B(n_15), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_214), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_188), .B(n_153), .Y(n_218) );
NOR2xp67_ASAP7_75t_L g219 ( .A(n_198), .B(n_164), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_194), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_214), .Y(n_221) );
OR2x6_ASAP7_75t_L g222 ( .A(n_208), .B(n_166), .Y(n_222) );
AND2x2_ASAP7_75t_L g223 ( .A(n_185), .B(n_154), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_216), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_214), .Y(n_225) );
CKINVDCx20_ASAP7_75t_R g226 ( .A(n_194), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_181), .B(n_165), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_214), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_181), .B(n_166), .Y(n_229) );
INVx1_ASAP7_75t_SL g230 ( .A(n_199), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_198), .A2(n_164), .B(n_166), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_212), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_212), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_199), .B(n_154), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_207), .B(n_166), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_180), .B(n_160), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_216), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_215), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_216), .Y(n_239) );
INVxp33_ASAP7_75t_L g240 ( .A(n_184), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_184), .B(n_161), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVxp67_ASAP7_75t_SL g243 ( .A(n_215), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_176), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_203), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_170), .Y(n_246) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_203), .B(n_161), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_170), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_170), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g250 ( .A(n_193), .B(n_161), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g251 ( .A(n_178), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_177), .B(n_154), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_177), .B(n_161), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g254 ( .A(n_195), .B(n_161), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_186), .B(n_161), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_186), .B(n_157), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_170), .Y(n_257) );
NOR2xp33_ASAP7_75t_SL g258 ( .A(n_213), .B(n_157), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_170), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_190), .Y(n_260) );
CKINVDCx20_ASAP7_75t_R g261 ( .A(n_178), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_190), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_190), .Y(n_263) );
BUFx6f_ASAP7_75t_SL g264 ( .A(n_209), .Y(n_264) );
XOR2xp5_ASAP7_75t_L g265 ( .A(n_202), .B(n_158), .Y(n_265) );
XOR2x2_ASAP7_75t_L g266 ( .A(n_196), .B(n_158), .Y(n_266) );
AND2x2_ASAP7_75t_L g267 ( .A(n_187), .B(n_158), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_173), .B(n_162), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_190), .Y(n_269) );
INVxp33_ASAP7_75t_L g270 ( .A(n_197), .Y(n_270) );
XNOR2xp5_ASAP7_75t_L g271 ( .A(n_202), .B(n_162), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_172), .A2(n_164), .B(n_160), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_205), .B(n_164), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_210), .B(n_155), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_217), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_224), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_217), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_256), .B(n_190), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_224), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
AND2x4_ASAP7_75t_L g281 ( .A(n_219), .B(n_167), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_224), .B(n_211), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_256), .B(n_173), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_231), .A2(n_175), .B(n_211), .Y(n_284) );
NOR2xp33_ASAP7_75t_R g285 ( .A(n_264), .B(n_171), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_267), .B(n_173), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_267), .B(n_173), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_221), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_224), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_270), .B(n_171), .Y(n_290) );
AND2x4_ASAP7_75t_L g291 ( .A(n_219), .B(n_167), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_221), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_268), .B(n_191), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_268), .B(n_191), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_238), .B(n_191), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_247), .B(n_191), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_245), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
INVx2_ASAP7_75t_SL g299 ( .A(n_237), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_225), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_247), .B(n_191), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_229), .A2(n_175), .B(n_211), .Y(n_302) );
INVx2_ASAP7_75t_SL g303 ( .A(n_237), .Y(n_303) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_245), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_247), .B(n_208), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_243), .B(n_175), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_234), .B(n_208), .Y(n_307) );
INVxp67_ASAP7_75t_L g308 ( .A(n_245), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_228), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_234), .B(n_222), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_245), .Y(n_311) );
INVx1_ASAP7_75t_SL g312 ( .A(n_245), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_218), .B(n_160), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_228), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_232), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_232), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_222), .B(n_208), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_222), .B(n_208), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_246), .Y(n_319) );
OAI21xp5_ASAP7_75t_L g320 ( .A1(n_235), .A2(n_172), .B(n_206), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_271), .B(n_160), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_233), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_222), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_233), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_222), .B(n_209), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_315), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_278), .B(n_240), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_278), .B(n_283), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_304), .Y(n_330) );
BUFx2_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_315), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_321), .B(n_265), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_278), .B(n_283), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_323), .B(n_246), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_321), .B(n_230), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_283), .B(n_271), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_283), .B(n_252), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_316), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_292), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_286), .B(n_252), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_323), .B(n_248), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_316), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_286), .B(n_255), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_323), .B(n_248), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_286), .B(n_265), .Y(n_349) );
AND2x4_ASAP7_75t_L g350 ( .A(n_323), .B(n_249), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_304), .Y(n_352) );
BUFx6f_ASAP7_75t_L g353 ( .A(n_304), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_292), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_285), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_316), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_327), .B(n_286), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_341), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_327), .B(n_287), .Y(n_361) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
BUFx4_ASAP7_75t_SL g363 ( .A(n_331), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_341), .Y(n_364) );
INVxp67_ASAP7_75t_SL g365 ( .A(n_341), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_343), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_330), .Y(n_367) );
INVx3_ASAP7_75t_L g368 ( .A(n_343), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_330), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_343), .Y(n_370) );
CKINVDCx20_ASAP7_75t_R g371 ( .A(n_331), .Y(n_371) );
INVx5_ASAP7_75t_L g372 ( .A(n_330), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_333), .B(n_251), .Y(n_373) );
NAND2x1p5_ASAP7_75t_L g374 ( .A(n_343), .B(n_317), .Y(n_374) );
INVx4_ASAP7_75t_L g375 ( .A(n_330), .Y(n_375) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_354), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_354), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_354), .B(n_287), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_354), .Y(n_380) );
INVx1_ASAP7_75t_SL g381 ( .A(n_352), .Y(n_381) );
BUFx4_ASAP7_75t_SL g382 ( .A(n_331), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_330), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_352), .Y(n_384) );
INVx5_ASAP7_75t_L g385 ( .A(n_330), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_355), .Y(n_386) );
OAI21xp5_ASAP7_75t_SL g387 ( .A1(n_374), .A2(n_301), .B(n_296), .Y(n_387) );
CKINVDCx16_ASAP7_75t_R g388 ( .A(n_371), .Y(n_388) );
BUFx8_ASAP7_75t_SL g389 ( .A(n_371), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_359), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_379), .B(n_327), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_364), .Y(n_392) );
INVx1_ASAP7_75t_SL g393 ( .A(n_372), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_365), .Y(n_394) );
AOI22xp5_ASAP7_75t_L g395 ( .A1(n_373), .A2(n_264), .B1(n_305), .B2(n_301), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_359), .B(n_357), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_373), .A2(n_305), .B1(n_296), .B2(n_301), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g398 ( .A1(n_386), .A2(n_264), .B1(n_301), .B2(n_296), .Y(n_398) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_359), .B(n_295), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_364), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_379), .B(n_332), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_372), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_386), .A2(n_296), .B1(n_305), .B2(n_318), .Y(n_403) );
AOI22xp33_ASAP7_75t_SL g404 ( .A1(n_374), .A2(n_305), .B1(n_318), .B2(n_317), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_364), .Y(n_406) );
BUFx3_ASAP7_75t_L g407 ( .A(n_372), .Y(n_407) );
BUFx12f_ASAP7_75t_L g408 ( .A(n_374), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_365), .A2(n_295), .B1(n_294), .B2(n_293), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_363), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_379), .A2(n_333), .B1(n_349), .B2(n_338), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g418 ( .A1(n_376), .A2(n_295), .B1(n_294), .B2(n_293), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_370), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_370), .Y(n_420) );
AOI22x1_ASAP7_75t_SL g421 ( .A1(n_363), .A2(n_261), .B1(n_220), .B2(n_226), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_379), .A2(n_337), .B1(n_258), .B2(n_287), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_370), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_376), .A2(n_293), .B1(n_294), .B2(n_318), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_374), .A2(n_333), .B1(n_349), .B2(n_338), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_358), .B(n_332), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_374), .A2(n_293), .B1(n_294), .B2(n_318), .Y(n_428) );
BUFx12f_ASAP7_75t_L g429 ( .A(n_375), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_358), .B(n_332), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_398), .A2(n_317), .B1(n_325), .B2(n_209), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_426), .A2(n_325), .B1(n_317), .B2(n_307), .Y(n_432) );
CKINVDCx5p33_ASAP7_75t_R g433 ( .A(n_389), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_325), .B1(n_209), .B2(n_355), .Y(n_434) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_395), .A2(n_394), .B1(n_408), .B2(n_403), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_429), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
BUFx2_ASAP7_75t_SL g438 ( .A(n_407), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_378), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_395), .A2(n_325), .B1(n_209), .B2(n_355), .Y(n_440) );
INVx5_ASAP7_75t_SL g441 ( .A(n_410), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_415), .B(n_378), .Y(n_442) );
NOR2x1_ASAP7_75t_R g443 ( .A(n_414), .B(n_382), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_394), .A2(n_380), .B1(n_337), .B2(n_339), .Y(n_444) );
INVx4_ASAP7_75t_L g445 ( .A(n_429), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_390), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_429), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_409), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_409), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_426), .A2(n_307), .B1(n_326), .B2(n_344), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_415), .B(n_380), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_422), .A2(n_227), .B1(n_250), .B2(n_266), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_392), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_394), .A2(n_408), .B1(n_403), .B2(n_404), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_407), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_411), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_407), .Y(n_457) );
INVx3_ASAP7_75t_L g458 ( .A(n_407), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_392), .Y(n_460) );
OAI22xp5_ASAP7_75t_L g461 ( .A1(n_404), .A2(n_380), .B1(n_346), .B2(n_339), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_411), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_422), .A2(n_307), .B1(n_326), .B2(n_340), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_413), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_428), .A2(n_307), .B1(n_344), .B2(n_340), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_388), .A2(n_357), .B1(n_346), .B2(n_342), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_413), .Y(n_467) );
AOI22xp33_ASAP7_75t_SL g468 ( .A1(n_388), .A2(n_385), .B1(n_372), .B2(n_368), .Y(n_468) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_428), .A2(n_340), .B1(n_344), .B2(n_329), .Y(n_469) );
INVx6_ASAP7_75t_L g470 ( .A(n_402), .Y(n_470) );
OAI22xp33_ASAP7_75t_L g471 ( .A1(n_414), .A2(n_342), .B1(n_346), .B2(n_361), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_392), .Y(n_472) );
BUFx2_ASAP7_75t_L g473 ( .A(n_402), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_387), .A2(n_342), .B1(n_361), .B2(n_319), .Y(n_474) );
OAI21xp5_ASAP7_75t_SL g475 ( .A1(n_387), .A2(n_287), .B(n_382), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_424), .A2(n_329), .B1(n_334), .B2(n_282), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_424), .A2(n_334), .B1(n_282), .B2(n_347), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_421), .B(n_155), .C(n_302), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_397), .A2(n_347), .B1(n_328), .B2(n_310), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_396), .B(n_328), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_391), .B(n_328), .Y(n_481) );
INVx4_ASAP7_75t_L g482 ( .A(n_410), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g483 ( .A1(n_397), .A2(n_347), .B1(n_310), .B2(n_266), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_412), .A2(n_310), .B1(n_368), .B2(n_284), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_400), .Y(n_485) );
AOI22xp33_ASAP7_75t_SL g486 ( .A1(n_421), .A2(n_385), .B1(n_372), .B2(n_368), .Y(n_486) );
INVx4_ASAP7_75t_L g487 ( .A(n_410), .Y(n_487) );
OAI22xp5_ASAP7_75t_L g488 ( .A1(n_393), .A2(n_319), .B1(n_368), .B2(n_310), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_416), .Y(n_489) );
OAI222xp33_ASAP7_75t_L g490 ( .A1(n_412), .A2(n_418), .B1(n_401), .B2(n_391), .C1(n_423), .C2(n_420), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_418), .A2(n_310), .B1(n_368), .B2(n_284), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_416), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_416), .A2(n_385), .B1(n_372), .B2(n_375), .Y(n_493) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_417), .A2(n_385), .B1(n_372), .B2(n_375), .Y(n_494) );
OAI222xp33_ASAP7_75t_L g495 ( .A1(n_401), .A2(n_384), .B1(n_381), .B2(n_375), .C1(n_385), .C2(n_372), .Y(n_495) );
OAI21xp33_ASAP7_75t_L g496 ( .A1(n_417), .A2(n_163), .B(n_162), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_400), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_417), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_478), .A2(n_168), .B1(n_163), .B2(n_284), .C(n_302), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_435), .A2(n_399), .B1(n_336), .B2(n_345), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g501 ( .A1(n_440), .A2(n_430), .B1(n_427), .B2(n_399), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_454), .A2(n_350), .B1(n_336), .B2(n_348), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_475), .A2(n_430), .B1(n_425), .B2(n_423), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_482), .B(n_419), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_482), .B(n_419), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_434), .A2(n_350), .B1(n_348), .B2(n_345), .Y(n_506) );
OAI22xp33_ASAP7_75t_SL g507 ( .A1(n_445), .A2(n_425), .B1(n_423), .B2(n_420), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_439), .B(n_420), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_483), .A2(n_348), .B1(n_336), .B2(n_345), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_437), .B(n_425), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_452), .A2(n_302), .B1(n_254), .B2(n_348), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_482), .B(n_400), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_483), .A2(n_336), .B1(n_348), .B2(n_345), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_466), .A2(n_163), .B1(n_168), .B2(n_274), .C(n_167), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_431), .A2(n_336), .B1(n_345), .B2(n_348), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g516 ( .A1(n_486), .A2(n_406), .B1(n_405), .B2(n_381), .Y(n_516) );
OA21x2_ASAP7_75t_L g517 ( .A1(n_495), .A2(n_383), .B(n_405), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_474), .A2(n_336), .B1(n_345), .B2(n_350), .Y(n_518) );
AOI222xp33_ASAP7_75t_L g519 ( .A1(n_490), .A2(n_168), .B1(n_306), .B2(n_281), .C1(n_291), .C2(n_167), .Y(n_519) );
OAI221xp5_ASAP7_75t_SL g520 ( .A1(n_450), .A2(n_306), .B1(n_167), .B2(n_150), .C(n_384), .Y(n_520) );
OAI222xp33_ASAP7_75t_L g521 ( .A1(n_445), .A2(n_375), .B1(n_405), .B2(n_406), .C1(n_372), .C2(n_385), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_450), .A2(n_350), .B1(n_281), .B2(n_291), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_487), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_468), .A2(n_406), .B1(n_385), .B2(n_375), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_471), .A2(n_385), .B1(n_306), .B2(n_377), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_463), .A2(n_350), .B1(n_291), .B2(n_281), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_463), .A2(n_350), .B1(n_291), .B2(n_281), .Y(n_527) );
OAI222xp33_ASAP7_75t_L g528 ( .A1(n_445), .A2(n_385), .B1(n_383), .B2(n_377), .C1(n_369), .C2(n_156), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_447), .B(n_150), .C(n_156), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_484), .A2(n_259), .B1(n_257), .B2(n_249), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_484), .A2(n_291), .B1(n_281), .B2(n_150), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_461), .A2(n_369), .B1(n_377), .B2(n_257), .Y(n_532) );
OAI222xp33_ASAP7_75t_L g533 ( .A1(n_436), .A2(n_383), .B1(n_377), .B2(n_369), .C1(n_156), .C2(n_269), .Y(n_533) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_447), .A2(n_369), .B1(n_367), .B2(n_362), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_436), .B(n_150), .C(n_156), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_487), .Y(n_536) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_438), .A2(n_367), .B1(n_362), .B2(n_383), .Y(n_537) );
OA21x2_ASAP7_75t_L g538 ( .A1(n_442), .A2(n_308), .B(n_356), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_441), .A2(n_263), .B1(n_259), .B2(n_260), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_487), .B(n_362), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_446), .B(n_156), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_448), .B(n_449), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_453), .Y(n_543) );
OAI211xp5_ASAP7_75t_SL g544 ( .A1(n_476), .A2(n_479), .B(n_469), .C(n_477), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_469), .A2(n_291), .B1(n_281), .B2(n_322), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_491), .A2(n_291), .B1(n_281), .B2(n_150), .Y(n_546) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_441), .A2(n_269), .B1(n_263), .B2(n_260), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_470), .A2(n_367), .B1(n_362), .B2(n_330), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_473), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_491), .A2(n_262), .B1(n_156), .B2(n_322), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_432), .A2(n_322), .B1(n_324), .B2(n_367), .Y(n_551) );
NAND3xp33_ASAP7_75t_L g552 ( .A(n_493), .B(n_304), .C(n_311), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_498), .B(n_362), .Y(n_553) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_470), .A2(n_367), .B1(n_362), .B2(n_353), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_455), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_465), .A2(n_253), .B1(n_297), .B2(n_312), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_476), .A2(n_367), .B1(n_362), .B2(n_304), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_465), .A2(n_367), .B1(n_304), .B2(n_311), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_456), .B(n_160), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_462), .B(n_160), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_451), .A2(n_311), .B1(n_280), .B2(n_289), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_480), .A2(n_311), .B1(n_280), .B2(n_289), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_494), .A2(n_297), .B1(n_312), .B2(n_290), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g564 ( .A1(n_444), .A2(n_312), .B1(n_353), .B2(n_335), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_496), .A2(n_433), .B1(n_481), .B2(n_457), .C(n_458), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_470), .A2(n_311), .B1(n_289), .B2(n_280), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_453), .B(n_15), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_464), .B(n_16), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_488), .A2(n_311), .B1(n_298), .B2(n_292), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_455), .A2(n_311), .B1(n_300), .B2(n_298), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_459), .B(n_353), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_467), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_489), .B(n_16), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g574 ( .A(n_459), .B(n_353), .C(n_351), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_492), .B(n_18), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_459), .A2(n_298), .B1(n_300), .B2(n_277), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_460), .B(n_19), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_459), .A2(n_298), .B1(n_300), .B2(n_277), .Y(n_578) );
OAI22x1_ASAP7_75t_L g579 ( .A1(n_460), .A2(n_20), .B1(n_21), .B2(n_23), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_472), .A2(n_298), .B1(n_300), .B2(n_277), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_497), .A2(n_300), .B1(n_288), .B2(n_309), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_497), .A2(n_275), .B1(n_309), .B2(n_288), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_485), .A2(n_275), .B1(n_309), .B2(n_288), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_485), .A2(n_275), .B1(n_314), .B2(n_335), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_443), .A2(n_241), .B1(n_273), .B2(n_255), .C(n_236), .Y(n_585) );
NAND3xp33_ASAP7_75t_L g586 ( .A(n_529), .B(n_353), .C(n_351), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_523), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_544), .A2(n_314), .B1(n_351), .B2(n_335), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_508), .B(n_504), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_521), .B(n_335), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_529), .B(n_351), .C(n_335), .Y(n_591) );
OA21x2_ASAP7_75t_L g592 ( .A1(n_552), .A2(n_320), .B(n_242), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_572), .B(n_21), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_572), .B(n_23), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_549), .B(n_24), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_542), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_501), .B(n_24), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_512), .B(n_26), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_512), .B(n_26), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_501), .B(n_27), .Y(n_600) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_499), .B(n_239), .C(n_320), .Y(n_601) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_503), .A2(n_223), .B(n_313), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_504), .B(n_27), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_505), .B(n_28), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_543), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_505), .B(n_28), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g607 ( .A1(n_502), .A2(n_320), .B1(n_313), .B2(n_314), .C(n_223), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_553), .B(n_29), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_579), .A2(n_313), .B1(n_192), .B2(n_206), .C(n_174), .Y(n_609) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_565), .A2(n_299), .B1(n_303), .B2(n_32), .C(n_33), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_535), .B(n_351), .C(n_276), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g612 ( .A(n_535), .B(n_276), .C(n_279), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_540), .B(n_30), .Y(n_613) );
NAND3xp33_ASAP7_75t_L g614 ( .A(n_519), .B(n_568), .C(n_552), .Y(n_614) );
NOR3xp33_ASAP7_75t_SL g615 ( .A(n_520), .B(n_30), .C(n_32), .Y(n_615) );
INVxp67_ASAP7_75t_SL g616 ( .A(n_507), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_567), .B(n_37), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_507), .A2(n_200), .B(n_176), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_516), .B(n_276), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_540), .B(n_37), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_579), .A2(n_174), .B1(n_189), .B2(n_192), .C(n_201), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_567), .B(n_38), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_536), .B(n_39), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_510), .B(n_40), .Y(n_624) );
NAND3xp33_ASAP7_75t_L g625 ( .A(n_519), .B(n_276), .C(n_279), .Y(n_625) );
OA21x2_ASAP7_75t_L g626 ( .A1(n_574), .A2(n_189), .B(n_176), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_500), .B(n_40), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_541), .B(n_42), .Y(n_628) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_509), .A2(n_303), .B1(n_299), .B2(n_204), .C(n_201), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_538), .B(n_45), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_573), .B(n_46), .Y(n_631) );
OAI221xp5_ASAP7_75t_SL g632 ( .A1(n_513), .A2(n_303), .B1(n_299), .B2(n_204), .C(n_201), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_575), .B(n_47), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_538), .B(n_555), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_577), .B(n_279), .C(n_276), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_555), .B(n_49), .Y(n_636) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_563), .B(n_279), .C(n_276), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_506), .B(n_50), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_511), .B(n_52), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_559), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_511), .B(n_54), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_518), .B(n_55), .Y(n_642) );
AOI221x1_ASAP7_75t_SL g643 ( .A1(n_530), .A2(n_204), .B1(n_183), .B2(n_182), .C(n_179), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_517), .B(n_56), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g645 ( .A(n_537), .B(n_279), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_515), .A2(n_279), .B1(n_276), .B2(n_303), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_532), .B(n_59), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_556), .A2(n_279), .B1(n_276), .B2(n_299), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_517), .B(n_557), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_525), .B(n_61), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_524), .A2(n_272), .B(n_276), .C(n_279), .Y(n_651) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_534), .A2(n_279), .B(n_276), .C(n_183), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_530), .B(n_62), .Y(n_653) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_574), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_560), .B(n_64), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_556), .B(n_66), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_545), .A2(n_279), .B1(n_183), .B2(n_182), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_581), .B(n_67), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_517), .B(n_548), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g660 ( .A1(n_528), .A2(n_71), .B(n_72), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_585), .B(n_182), .C(n_179), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_554), .B(n_73), .Y(n_662) );
NOR2xp33_ASAP7_75t_SL g663 ( .A(n_533), .B(n_75), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_514), .B(n_179), .C(n_78), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_551), .B(n_77), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_545), .A2(n_79), .B1(n_80), .B2(n_82), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_522), .A2(n_244), .B1(n_84), .B2(n_85), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_531), .A2(n_83), .B1(n_86), .B2(n_87), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_582), .B(n_90), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_583), .B(n_91), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_517), .B(n_93), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_580), .B(n_94), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_550), .B(n_569), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_561), .B(n_96), .Y(n_674) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_558), .B(n_97), .C(n_98), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_564), .B(n_99), .Y(n_676) );
INVx2_ASAP7_75t_L g677 ( .A(n_571), .Y(n_677) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_598), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_596), .B(n_584), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_587), .B(n_570), .C(n_562), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_614), .A2(n_673), .B1(n_625), .B2(n_640), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_598), .B(n_547), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_605), .B(n_578), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_610), .A2(n_526), .B1(n_527), .B2(n_546), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_620), .B(n_566), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_620), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_608), .B(n_576), .Y(n_687) );
NOR3xp33_ASAP7_75t_L g688 ( .A(n_595), .B(n_539), .C(n_102), .Y(n_688) );
NAND4xp25_ASAP7_75t_L g689 ( .A(n_588), .B(n_244), .C(n_602), .D(n_597), .Y(n_689) );
BUFx3_ASAP7_75t_L g690 ( .A(n_634), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_590), .A2(n_645), .B(n_619), .Y(n_691) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_660), .A2(n_618), .B(n_588), .C(n_600), .Y(n_692) );
NAND4xp75_ASAP7_75t_L g693 ( .A(n_599), .B(n_604), .C(n_603), .D(n_608), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_645), .B(n_659), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_624), .B(n_594), .C(n_593), .Y(n_695) );
AND2x4_ASAP7_75t_SL g696 ( .A(n_603), .B(n_604), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g697 ( .A(n_651), .B(n_659), .C(n_619), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_637), .B(n_649), .C(n_606), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_623), .B(n_643), .Y(n_699) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_627), .B(n_617), .C(n_622), .Y(n_700) );
NAND4xp75_ASAP7_75t_L g701 ( .A(n_649), .B(n_623), .C(n_671), .D(n_644), .Y(n_701) );
NAND4xp75_ASAP7_75t_L g702 ( .A(n_644), .B(n_671), .C(n_639), .D(n_641), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_661), .B(n_664), .C(n_633), .Y(n_703) );
OR2x2_ASAP7_75t_L g704 ( .A(n_677), .B(n_635), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_609), .B(n_621), .C(n_612), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_615), .A2(n_632), .B1(n_611), .B2(n_648), .Y(n_706) );
OAI221xp5_ASAP7_75t_L g707 ( .A1(n_663), .A2(n_667), .B1(n_607), .B2(n_631), .C(n_656), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_630), .B(n_592), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g709 ( .A(n_646), .Y(n_709) );
NAND4xp75_ASAP7_75t_L g710 ( .A(n_592), .B(n_650), .C(n_642), .D(n_638), .Y(n_710) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_592), .B(n_653), .C(n_647), .D(n_636), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_601), .A2(n_655), .B1(n_628), .B2(n_665), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_586), .B(n_591), .Y(n_713) );
AOI22x1_ASAP7_75t_L g714 ( .A1(n_652), .A2(n_667), .B1(n_675), .B2(n_666), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_626), .B(n_676), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g716 ( .A(n_662), .B(n_657), .C(n_670), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_669), .A2(n_629), .B1(n_658), .B2(n_672), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_674), .B(n_668), .Y(n_718) );
AND4x1_ASAP7_75t_L g719 ( .A(n_590), .B(n_663), .C(n_615), .D(n_625), .Y(n_719) );
AND2x4_ASAP7_75t_L g720 ( .A(n_634), .B(n_587), .Y(n_720) );
NAND4xp75_ASAP7_75t_L g721 ( .A(n_598), .B(n_599), .C(n_620), .D(n_613), .Y(n_721) );
NAND4xp75_ASAP7_75t_L g722 ( .A(n_598), .B(n_599), .C(n_620), .D(n_613), .Y(n_722) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_616), .B(n_587), .C(n_654), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_616), .A2(n_435), .B1(n_590), .B2(n_454), .Y(n_724) );
NOR3xp33_ASAP7_75t_L g725 ( .A(n_610), .B(n_595), .C(n_597), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_610), .B(n_595), .C(n_597), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_590), .B(n_507), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_616), .A2(n_596), .B1(n_614), .B2(n_595), .C(n_600), .Y(n_728) );
OR2x2_ASAP7_75t_L g729 ( .A(n_589), .B(n_587), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_616), .B(n_587), .C(n_654), .Y(n_730) );
NAND3xp33_ASAP7_75t_L g731 ( .A(n_616), .B(n_587), .C(n_654), .Y(n_731) );
NOR4xp25_ASAP7_75t_SL g732 ( .A(n_727), .B(n_728), .C(n_678), .D(n_682), .Y(n_732) );
XOR2x2_ASAP7_75t_L g733 ( .A(n_693), .B(n_721), .Y(n_733) );
INVx2_ASAP7_75t_SL g734 ( .A(n_690), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_724), .A2(n_725), .B1(n_726), .B2(n_722), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_690), .B(n_720), .Y(n_736) );
NAND4xp75_ASAP7_75t_SL g737 ( .A(n_718), .B(n_715), .C(n_724), .D(n_719), .Y(n_737) );
NAND4xp75_ASAP7_75t_L g738 ( .A(n_727), .B(n_691), .C(n_699), .D(n_694), .Y(n_738) );
NOR4xp25_ASAP7_75t_L g739 ( .A(n_723), .B(n_731), .C(n_730), .D(n_681), .Y(n_739) );
XOR2xp5_ASAP7_75t_L g740 ( .A(n_709), .B(n_701), .Y(n_740) );
XNOR2x2_ASAP7_75t_L g741 ( .A(n_697), .B(n_694), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_729), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_720), .Y(n_743) );
NAND4xp75_ASAP7_75t_L g744 ( .A(n_679), .B(n_687), .C(n_685), .D(n_708), .Y(n_744) );
XNOR2x1_ASAP7_75t_L g745 ( .A(n_702), .B(n_686), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_696), .Y(n_746) );
AND2x2_ASAP7_75t_L g747 ( .A(n_704), .B(n_698), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_683), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_713), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_705), .Y(n_750) );
HB1xp67_ASAP7_75t_L g751 ( .A(n_680), .Y(n_751) );
NOR3xp33_ASAP7_75t_L g752 ( .A(n_692), .B(n_707), .C(n_716), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_695), .B(n_700), .Y(n_753) );
NAND4xp75_ASAP7_75t_SL g754 ( .A(n_711), .B(n_710), .C(n_714), .D(n_689), .Y(n_754) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_706), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_700), .Y(n_756) );
INVx2_ASAP7_75t_SL g757 ( .A(n_688), .Y(n_757) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_703), .A2(n_716), .B1(n_712), .B2(n_717), .Y(n_758) );
INVx1_ASAP7_75t_SL g759 ( .A(n_746), .Y(n_759) );
INVxp67_ASAP7_75t_L g760 ( .A(n_755), .Y(n_760) );
XOR2x2_ASAP7_75t_L g761 ( .A(n_733), .B(n_737), .Y(n_761) );
INVxp67_ASAP7_75t_SL g762 ( .A(n_741), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_745), .A2(n_712), .B1(n_717), .B2(n_684), .Y(n_763) );
AND2x2_ASAP7_75t_L g764 ( .A(n_749), .B(n_703), .Y(n_764) );
INVxp67_ASAP7_75t_SL g765 ( .A(n_741), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_733), .Y(n_766) );
INVxp33_ASAP7_75t_L g767 ( .A(n_740), .Y(n_767) );
INVxp33_ASAP7_75t_SL g768 ( .A(n_735), .Y(n_768) );
XNOR2xp5_ASAP7_75t_L g769 ( .A(n_740), .B(n_684), .Y(n_769) );
OA22x2_ASAP7_75t_L g770 ( .A1(n_758), .A2(n_750), .B1(n_751), .B2(n_756), .Y(n_770) );
XNOR2x1_ASAP7_75t_L g771 ( .A(n_738), .B(n_754), .Y(n_771) );
BUFx2_ASAP7_75t_L g772 ( .A(n_734), .Y(n_772) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_752), .A2(n_757), .B1(n_753), .B2(n_756), .Y(n_773) );
XNOR2xp5_ASAP7_75t_L g774 ( .A(n_745), .B(n_744), .Y(n_774) );
INVxp67_ASAP7_75t_L g775 ( .A(n_738), .Y(n_775) );
XNOR2xp5_ASAP7_75t_L g776 ( .A(n_757), .B(n_739), .Y(n_776) );
OA22x2_ASAP7_75t_L g777 ( .A1(n_774), .A2(n_747), .B1(n_734), .B2(n_732), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_759), .Y(n_778) );
AO22x1_ASAP7_75t_L g779 ( .A1(n_762), .A2(n_747), .B1(n_743), .B2(n_736), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_761), .B(n_748), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_772), .Y(n_781) );
XNOR2xp5_ASAP7_75t_L g782 ( .A(n_761), .B(n_742), .Y(n_782) );
INVx2_ASAP7_75t_SL g783 ( .A(n_772), .Y(n_783) );
BUFx3_ASAP7_75t_L g784 ( .A(n_771), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_778), .B(n_760), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_783), .Y(n_786) );
INVx1_ASAP7_75t_L g787 ( .A(n_783), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_780), .B(n_765), .Y(n_788) );
INVx5_ASAP7_75t_L g789 ( .A(n_781), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_781), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_785), .Y(n_791) );
INVx2_ASAP7_75t_L g792 ( .A(n_790), .Y(n_792) );
AO22x2_ASAP7_75t_L g793 ( .A1(n_788), .A2(n_784), .B1(n_771), .B2(n_763), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_785), .Y(n_794) );
NOR4xp25_ASAP7_75t_L g795 ( .A(n_788), .B(n_775), .C(n_770), .D(n_784), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_792), .Y(n_796) );
OAI221xp5_ASAP7_75t_L g797 ( .A1(n_795), .A2(n_776), .B1(n_777), .B2(n_770), .C(n_780), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_792), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_796), .Y(n_799) );
INVx1_ASAP7_75t_L g800 ( .A(n_798), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_799), .Y(n_801) );
HB1xp67_ASAP7_75t_L g802 ( .A(n_800), .Y(n_802) );
AO22x2_ASAP7_75t_L g803 ( .A1(n_801), .A2(n_794), .B1(n_791), .B2(n_787), .Y(n_803) );
AOI22x1_ASAP7_75t_L g804 ( .A1(n_802), .A2(n_793), .B1(n_776), .B2(n_782), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_803), .Y(n_805) );
BUFx2_ASAP7_75t_L g806 ( .A(n_804), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g807 ( .A1(n_806), .A2(n_793), .B1(n_797), .B2(n_766), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_807), .Y(n_808) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_808), .A2(n_793), .B1(n_805), .B2(n_768), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_809), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_810), .A2(n_786), .B1(n_782), .B2(n_767), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_811), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g813 ( .A1(n_812), .A2(n_779), .B1(n_789), .B2(n_773), .C(n_769), .Y(n_813) );
AOI211xp5_ASAP7_75t_L g814 ( .A1(n_813), .A2(n_769), .B(n_773), .C(n_764), .Y(n_814) );
endmodule