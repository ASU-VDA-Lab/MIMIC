module fake_ibex_447_n_367 (n_85, n_84, n_64, n_3, n_73, n_65, n_95, n_55, n_63, n_29, n_2, n_76, n_8, n_67, n_9, n_38, n_37, n_47, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_48, n_57, n_59, n_28, n_39, n_5, n_62, n_71, n_93, n_13, n_61, n_14, n_0, n_94, n_12, n_42, n_77, n_88, n_44, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_22, n_4, n_33, n_30, n_6, n_72, n_26, n_34, n_15, n_24, n_52, n_1, n_25, n_36, n_41, n_45, n_18, n_89, n_83, n_32, n_53, n_50, n_11, n_92, n_68, n_79, n_81, n_35, n_31, n_56, n_23, n_91, n_54, n_19, n_367);

input n_85;
input n_84;
input n_64;
input n_3;
input n_73;
input n_65;
input n_95;
input n_55;
input n_63;
input n_29;
input n_2;
input n_76;
input n_8;
input n_67;
input n_9;
input n_38;
input n_37;
input n_47;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_48;
input n_57;
input n_59;
input n_28;
input n_39;
input n_5;
input n_62;
input n_71;
input n_93;
input n_13;
input n_61;
input n_14;
input n_0;
input n_94;
input n_12;
input n_42;
input n_77;
input n_88;
input n_44;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_22;
input n_4;
input n_33;
input n_30;
input n_6;
input n_72;
input n_26;
input n_34;
input n_15;
input n_24;
input n_52;
input n_1;
input n_25;
input n_36;
input n_41;
input n_45;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_50;
input n_11;
input n_92;
input n_68;
input n_79;
input n_81;
input n_35;
input n_31;
input n_56;
input n_23;
input n_91;
input n_54;
input n_19;

output n_367;

wire n_151;
wire n_171;
wire n_103;
wire n_204;
wire n_274;
wire n_130;
wire n_177;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_293;
wire n_341;
wire n_124;
wire n_256;
wire n_193;
wire n_108;
wire n_350;
wire n_165;
wire n_255;
wire n_175;
wire n_125;
wire n_304;
wire n_191;
wire n_153;
wire n_194;
wire n_249;
wire n_334;
wire n_312;
wire n_239;
wire n_134;
wire n_357;
wire n_142;
wire n_226;
wire n_336;
wire n_258;
wire n_176;
wire n_216;
wire n_166;
wire n_163;
wire n_114;
wire n_236;
wire n_189;
wire n_280;
wire n_317;
wire n_340;
wire n_105;
wire n_187;
wire n_154;
wire n_182;
wire n_196;
wire n_327;
wire n_326;
wire n_170;
wire n_144;
wire n_270;
wire n_346;
wire n_113;
wire n_117;
wire n_265;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_210;
wire n_348;
wire n_220;
wire n_287;
wire n_243;
wire n_228;
wire n_147;
wire n_251;
wire n_244;
wire n_343;
wire n_310;
wire n_323;
wire n_143;
wire n_106;
wire n_224;
wire n_183;
wire n_333;
wire n_110;
wire n_306;
wire n_169;
wire n_242;
wire n_278;
wire n_316;
wire n_109;
wire n_127;
wire n_121;
wire n_325;
wire n_301;
wire n_296;
wire n_120;
wire n_168;
wire n_155;
wire n_315;
wire n_122;
wire n_116;
wire n_289;
wire n_150;
wire n_286;
wire n_321;
wire n_133;
wire n_215;
wire n_279;
wire n_235;
wire n_136;
wire n_261;
wire n_221;
wire n_355;
wire n_102;
wire n_99;
wire n_269;
wire n_156;
wire n_126;
wire n_356;
wire n_104;
wire n_141;
wire n_222;
wire n_186;
wire n_349;
wire n_295;
wire n_331;
wire n_230;
wire n_96;
wire n_185;
wire n_352;
wire n_290;
wire n_174;
wire n_157;
wire n_219;
wire n_246;
wire n_146;
wire n_207;
wire n_167;
wire n_128;
wire n_253;
wire n_208;
wire n_234;
wire n_152;
wire n_300;
wire n_145;
wire n_358;
wire n_205;
wire n_139;
wire n_275;
wire n_98;
wire n_129;
wire n_267;
wire n_245;
wire n_229;
wire n_209;
wire n_347;
wire n_335;
wire n_263;
wire n_353;
wire n_359;
wire n_299;
wire n_262;
wire n_137;
wire n_338;
wire n_173;
wire n_363;
wire n_180;
wire n_201;
wire n_351;
wire n_257;
wire n_305;
wire n_307;
wire n_192;
wire n_140;
wire n_365;
wire n_100;
wire n_179;
wire n_354;
wire n_206;
wire n_329;
wire n_188;
wire n_200;
wire n_199;
wire n_308;
wire n_135;
wire n_283;
wire n_366;
wire n_111;
wire n_322;
wire n_227;
wire n_115;
wire n_248;
wire n_101;
wire n_190;
wire n_138;
wire n_238;
wire n_214;
wire n_332;
wire n_211;
wire n_218;
wire n_314;
wire n_132;
wire n_277;
wire n_337;
wire n_225;
wire n_360;
wire n_272;
wire n_223;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_291;
wire n_318;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_148;
wire n_342;
wire n_233;
wire n_118;
wire n_164;
wire n_198;
wire n_264;
wire n_217;
wire n_324;
wire n_178;
wire n_303;
wire n_362;
wire n_162;
wire n_240;
wire n_282;
wire n_266;
wire n_294;
wire n_112;
wire n_284;
wire n_172;
wire n_250;
wire n_313;
wire n_345;
wire n_119;
wire n_361;
wire n_319;
wire n_195;
wire n_212;
wire n_311;
wire n_97;
wire n_197;
wire n_181;
wire n_131;
wire n_123;
wire n_260;
wire n_302;
wire n_344;
wire n_297;
wire n_252;
wire n_107;
wire n_149;
wire n_254;
wire n_213;
wire n_271;
wire n_241;
wire n_292;
wire n_364;
wire n_159;
wire n_231;
wire n_202;
wire n_298;
wire n_160;
wire n_184;
wire n_232;
wire n_281;

INVxp67_ASAP7_75t_L g96 ( 
.A(n_75),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_24),
.Y(n_98)
);

INVxp67_ASAP7_75t_SL g99 ( 
.A(n_54),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVxp33_ASAP7_75t_SL g105 ( 
.A(n_44),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_95),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_87),
.Y(n_115)
);

INVxp33_ASAP7_75t_SL g116 ( 
.A(n_42),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_67),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVxp33_ASAP7_75t_SL g120 ( 
.A(n_83),
.Y(n_120)
);

INVxp33_ASAP7_75t_SL g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_31),
.Y(n_122)
);

CKINVDCx5p33_ASAP7_75t_R g123 ( 
.A(n_52),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_4),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_59),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_37),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_13),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_0),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_19),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_49),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_32),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_88),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_86),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_26),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_22),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_64),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_27),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_36),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_4),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_16),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_63),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_82),
.Y(n_152)
);

INVxp33_ASAP7_75t_SL g153 ( 
.A(n_25),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_12),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVxp33_ASAP7_75t_SL g158 ( 
.A(n_1),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_62),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_89),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_20),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_71),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_51),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_50),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_29),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_40),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_47),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_18),
.Y(n_171)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_7),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_74),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_14),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_45),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_23),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_46),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_2),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_57),
.Y(n_181)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_17),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_43),
.Y(n_183)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_132),
.B(n_0),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_170),
.Y(n_188)
);

AND3x2_ASAP7_75t_L g189 ( 
.A(n_146),
.B(n_180),
.C(n_181),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_1),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_155),
.B(n_168),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g192 ( 
.A(n_124),
.B(n_3),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_117),
.B(n_3),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g194 ( 
.A1(n_150),
.A2(n_5),
.B1(n_10),
.B2(n_21),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_157),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_103),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_101),
.B(n_28),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_102),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_158),
.B(n_30),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_98),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_122),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_110),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_111),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_112),
.Y(n_209)
);

AND3x2_ASAP7_75t_L g210 ( 
.A(n_99),
.B(n_56),
.C(n_85),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_119),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_125),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_126),
.B(n_183),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_L g217 ( 
.A(n_106),
.B(n_176),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_127),
.B(n_178),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_137),
.B(n_162),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_139),
.B(n_142),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_99),
.B(n_181),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_140),
.B(n_152),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_143),
.B(n_179),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_113),
.A2(n_153),
.B1(n_105),
.B2(n_116),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_145),
.B(n_169),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_147),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_120),
.A2(n_121),
.B1(n_177),
.B2(n_175),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_167),
.B(n_96),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_128),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_123),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_143),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_96),
.B(n_174),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_179),
.Y(n_239)
);

BUFx6f_ASAP7_75t_SL g240 ( 
.A(n_141),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_136),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_174),
.Y(n_243)
);

AND2x6_ASAP7_75t_SL g244 ( 
.A(n_192),
.B(n_161),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_203),
.B(n_136),
.Y(n_246)
);

OR2x6_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_149),
.Y(n_247)
);

BUFx4f_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NOR2x1p5_ASAP7_75t_L g249 ( 
.A(n_186),
.B(n_182),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_192),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_149),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_156),
.B1(n_151),
.B2(n_172),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_241),
.B(n_131),
.Y(n_254)
);

NOR3xp33_ASAP7_75t_SL g255 ( 
.A(n_187),
.B(n_135),
.C(n_138),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_188),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_185),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_196),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_197),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_184),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_184),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_236),
.B(n_160),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_225),
.B(n_173),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_198),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

AND2x4_ASAP7_75t_L g270 ( 
.A(n_239),
.B(n_164),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g271 ( 
.A(n_241),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_165),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_210),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_193),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_235),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_214),
.B(n_211),
.Y(n_277)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_200),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_215),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_205),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_231),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_233),
.B(n_227),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_209),
.B(n_218),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_204),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_189),
.Y(n_286)
);

AND3x1_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_206),
.C(n_222),
.Y(n_287)
);

BUFx4f_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_216),
.B(n_228),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_240),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_222),
.B(n_224),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_221),
.A2(n_189),
.B1(n_217),
.B2(n_202),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_240),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_243),
.B(n_224),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_269),
.Y(n_296)
);

OAI21x1_ASAP7_75t_SL g297 ( 
.A1(n_286),
.A2(n_206),
.B(n_199),
.Y(n_297)
);

OA21x2_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_199),
.B(n_191),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_292),
.B(n_226),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_249),
.B(n_219),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_262),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_274),
.B(n_220),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_257),
.A2(n_252),
.B(n_273),
.Y(n_303)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_229),
.Y(n_304)
);

AO31x2_ASAP7_75t_L g305 ( 
.A1(n_282),
.A2(n_230),
.A3(n_232),
.B(n_194),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g306 ( 
.A1(n_284),
.A2(n_194),
.B(n_210),
.C(n_290),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_254),
.A2(n_277),
.B(n_256),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_281),
.A2(n_285),
.B(n_246),
.C(n_268),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

OAI21x1_ASAP7_75t_L g310 ( 
.A1(n_245),
.A2(n_260),
.B(n_264),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_279),
.Y(n_311)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_272),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_274),
.B(n_293),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_287),
.A2(n_283),
.B1(n_247),
.B2(n_270),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_247),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_288),
.B(n_271),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_275),
.Y(n_318)
);

AOI21x1_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_255),
.B(n_291),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_301),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_306),
.A2(n_258),
.B(n_261),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_263),
.B(n_253),
.Y(n_322)
);

AOI21x1_ASAP7_75t_SL g323 ( 
.A1(n_311),
.A2(n_294),
.B(n_248),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_315),
.A2(n_295),
.B1(n_296),
.B2(n_314),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_276),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_280),
.Y(n_326)
);

OR2x6_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_244),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_288),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_308),
.A2(n_248),
.B1(n_278),
.B2(n_265),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_265),
.B1(n_278),
.B2(n_304),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_312),
.A2(n_265),
.B1(n_278),
.B2(n_304),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_307),
.Y(n_332)
);

BUFx8_ASAP7_75t_L g333 ( 
.A(n_300),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

AOI211xp5_ASAP7_75t_L g335 ( 
.A1(n_300),
.A2(n_317),
.B(n_302),
.C(n_309),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_305),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_320),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_305),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_333),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_332),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_322),
.Y(n_342)
);

NOR4xp25_ASAP7_75t_SL g343 ( 
.A(n_327),
.B(n_305),
.C(n_298),
.D(n_303),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_298),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_327),
.B(n_321),
.Y(n_346)
);

BUFx8_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_337),
.Y(n_348)
);

OR2x6_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_327),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_345),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_339),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_345),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_351),
.B(n_344),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_338),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g356 ( 
.A(n_349),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_353),
.Y(n_357)
);

NOR2x1p5_ASAP7_75t_L g358 ( 
.A(n_354),
.B(n_346),
.Y(n_358)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_349),
.B(n_326),
.Y(n_359)
);

A2O1A1Ixp33_ASAP7_75t_L g360 ( 
.A1(n_358),
.A2(n_356),
.B(n_338),
.C(n_355),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_359),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_361),
.B(n_360),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_336),
.A3(n_352),
.B1(n_347),
.B2(n_342),
.C1(n_319),
.C2(n_343),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_363),
.A2(n_342),
.B1(n_341),
.B2(n_322),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_364),
.A2(n_333),
.B1(n_330),
.B2(n_331),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_365),
.A2(n_341),
.B1(n_329),
.B2(n_335),
.Y(n_366)
);

AOI221xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_323),
.B1(n_335),
.B2(n_341),
.C(n_365),
.Y(n_367)
);


endmodule