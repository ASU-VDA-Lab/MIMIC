module fake_jpeg_21871_n_74 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_74);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_64;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_73;
wire n_20;
wire n_59;
wire n_71;
wire n_48;
wire n_35;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_72;
wire n_49;
wire n_44;
wire n_28;
wire n_24;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_25;
wire n_67;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;
wire n_70;
wire n_66;

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_19),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_10),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_30),
.B(n_2),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_29),
.B(n_4),
.CON(n_42),
.SN(n_42)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_45),
.C(n_46),
.Y(n_57)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_6),
.B(n_9),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_23),
.B(n_17),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_54),
.A2(n_42),
.B(n_33),
.C(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_50),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_39),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_43),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_63),
.B(n_60),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_50),
.B(n_25),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_57),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_57),
.C(n_55),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_68),
.A2(n_22),
.B1(n_24),
.B2(n_38),
.Y(n_70)
);

OAI31xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_70),
.A3(n_53),
.B(n_32),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_18),
.C(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_52),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_49),
.Y(n_74)
);


endmodule