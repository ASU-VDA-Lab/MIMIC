module fake_jpeg_19982_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx5_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_8),
.B(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_16),
.B(n_19),
.C(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_22),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_29),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_35),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_42),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_24),
.B1(n_25),
.B2(n_16),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_17),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_49),
.B(n_60),
.Y(n_75)
);

OAI22x1_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_50),
.A2(n_37),
.B1(n_39),
.B2(n_43),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_25),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_56),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_30),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_55),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_30),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_21),
.C(n_31),
.Y(n_56)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_40),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_32),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_57),
.A2(n_39),
.B1(n_43),
.B2(n_37),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_65),
.A2(n_59),
.B(n_47),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_47),
.C(n_50),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_56),
.C(n_48),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_53),
.A2(n_41),
.B1(n_15),
.B2(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_15),
.B1(n_12),
.B2(n_3),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_80),
.B(n_76),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_54),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_88),
.C(n_84),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_56),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_89),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_12),
.B(n_2),
.C(n_3),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_92),
.B(n_101),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_86),
.C(n_81),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_70),
.C(n_62),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_102),
.C(n_93),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_68),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_97),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_90),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_83),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_69),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_105),
.C(n_108),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_64),
.C(n_87),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_79),
.B1(n_75),
.B2(n_72),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_91),
.B1(n_101),
.B2(n_96),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_111),
.B(n_99),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_79),
.B1(n_99),
.B2(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_98),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_107),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_102),
.C(n_77),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_105),
.C(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_124),
.B(n_9),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_112),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g129 ( 
.A1(n_125),
.A2(n_128),
.A3(n_120),
.B1(n_119),
.B2(n_9),
.C1(n_51),
.C2(n_0),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_100),
.B(n_11),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_51),
.A3(n_2),
.B1(n_4),
.B2(n_5),
.C(n_6),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_131),
.B(n_5),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_0),
.B(n_2),
.C(n_4),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_125),
.C(n_51),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);


endmodule