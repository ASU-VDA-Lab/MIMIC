module fake_jpeg_31758_n_62 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_62);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_62;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

INVx11_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_22),
.Y(n_28)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_25),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_10),
.B1(n_14),
.B2(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_12),
.B(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_14),
.B1(n_17),
.B2(n_11),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_15),
.C(n_8),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_26),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_24),
.A2(n_13),
.B(n_10),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_1),
.B(n_2),
.Y(n_37)
);

NAND3xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_17),
.C(n_12),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_3),
.B(n_4),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_41),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_27),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_23),
.B1(n_26),
.B2(n_20),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_26),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_45),
.A2(n_41),
.B1(n_30),
.B2(n_23),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_39),
.C(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_50),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_51),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_37),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_11),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_52),
.B(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_50),
.B1(n_49),
.B2(n_45),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_57),
.A2(n_55),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_4),
.C(n_5),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_57),
.B(n_59),
.C(n_11),
.D(n_20),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_31),
.Y(n_62)
);


endmodule