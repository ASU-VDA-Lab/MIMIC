module fake_jpeg_32003_n_518 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_518);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_518;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_16),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_16),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_5),
.Y(n_48)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_50),
.Y(n_110)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_17),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_52),
.B(n_87),
.Y(n_127)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_64),
.Y(n_125)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_66),
.Y(n_161)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_70),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_43),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_73),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_74),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_18),
.B(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_19),
.Y(n_107)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_76),
.Y(n_157)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_81),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_84),
.Y(n_139)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_17),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_91),
.B(n_92),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_45),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_93),
.Y(n_149)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_95),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_96),
.Y(n_122)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

BUFx10_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_100),
.A2(n_21),
.B1(n_22),
.B2(n_49),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_103),
.A2(n_130),
.B1(n_156),
.B2(n_4),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_107),
.B(n_114),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_52),
.B(n_38),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_142),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_57),
.B(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_126),
.B(n_128),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_24),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_36),
.B1(n_49),
.B2(n_34),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_129),
.B(n_138),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_62),
.A2(n_21),
.B1(n_22),
.B2(n_49),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_94),
.B(n_44),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_98),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_76),
.B(n_44),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_93),
.C(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_70),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_53),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_58),
.A2(n_44),
.B1(n_48),
.B2(n_42),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_177)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_72),
.A2(n_22),
.B1(n_40),
.B2(n_31),
.Y(n_156)
);

NAND2x1_ASAP7_75t_SL g158 ( 
.A(n_89),
.B(n_22),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_158),
.A2(n_162),
.B(n_2),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_79),
.A2(n_15),
.B(n_14),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_133),
.Y(n_165)
);

BUFx2_ASAP7_75t_SL g263 ( 
.A(n_165),
.Y(n_263)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_166),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_158),
.A2(n_84),
.B1(n_31),
.B2(n_48),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_97),
.B1(n_69),
.B2(n_90),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_169),
.A2(n_177),
.B1(n_201),
.B2(n_216),
.Y(n_244)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_136),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_171),
.B(n_178),
.Y(n_246)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_173),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_127),
.B(n_25),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_184),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_176),
.Y(n_227)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_180),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_181),
.B(n_185),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_123),
.B(n_83),
.C(n_81),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_219),
.C(n_160),
.Y(n_254)
);

CKINVDCx12_ASAP7_75t_R g183 ( 
.A(n_122),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_30),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_186),
.Y(n_238)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_113),
.Y(n_187)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_187),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_31),
.B1(n_80),
.B2(n_55),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g252 ( 
.A1(n_188),
.A2(n_215),
.B(n_117),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_103),
.B1(n_130),
.B2(n_155),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_190),
.A2(n_148),
.B1(n_115),
.B2(n_145),
.Y(n_253)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_119),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_192),
.B(n_214),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_111),
.B(n_42),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_193),
.B(n_195),
.Y(n_245)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_127),
.B(n_39),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_196),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_159),
.A2(n_39),
.B1(n_30),
.B2(n_28),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_197),
.A2(n_199),
.B1(n_139),
.B2(n_116),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_207),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_119),
.A2(n_28),
.B1(n_27),
.B2(n_25),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_153),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

BUFx16f_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_138),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_205),
.A2(n_5),
.B(n_6),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_206),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_122),
.B(n_133),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_102),
.Y(n_208)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_141),
.Y(n_209)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_143),
.B(n_0),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_211),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_124),
.B(n_0),
.Y(n_211)
);

BUFx12_ASAP7_75t_L g212 ( 
.A(n_141),
.Y(n_212)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_124),
.B(n_1),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_153),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_101),
.Y(n_217)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_218),
.A2(n_108),
.B1(n_154),
.B2(n_149),
.Y(n_228)
);

AND2x2_ASAP7_75t_SL g219 ( 
.A(n_157),
.B(n_4),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_121),
.Y(n_220)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_104),
.Y(n_222)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_222),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_228),
.A2(n_230),
.B1(n_243),
.B2(n_253),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_177),
.B1(n_190),
.B2(n_108),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_242),
.A2(n_264),
.B(n_269),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_149),
.B1(n_148),
.B2(n_115),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_254),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g257 ( 
.A(n_188),
.B(n_109),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_188),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_202),
.A2(n_160),
.B1(n_145),
.B2(n_140),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_179),
.B1(n_166),
.B2(n_192),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_117),
.B(n_6),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_188),
.A2(n_140),
.B1(n_151),
.B2(n_139),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_266),
.A2(n_187),
.B1(n_168),
.B2(n_163),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_267),
.Y(n_272)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

INVx13_ASAP7_75t_L g274 ( 
.A(n_225),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_274),
.Y(n_332)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_225),
.Y(n_276)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_277),
.A2(n_312),
.B1(n_313),
.B2(n_315),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_L g278 ( 
.A1(n_227),
.A2(n_213),
.B(n_219),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_278),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_223),
.B(n_231),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_279),
.B(n_286),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_292),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_244),
.A2(n_219),
.B1(n_178),
.B2(n_172),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_281),
.A2(n_283),
.B1(n_291),
.B2(n_305),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_229),
.A2(n_165),
.B1(n_196),
.B2(n_189),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_282),
.A2(n_308),
.B1(n_226),
.B2(n_259),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_257),
.A2(n_180),
.B1(n_170),
.B2(n_194),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_254),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g336 ( 
.A(n_285),
.B(n_116),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_245),
.B(n_203),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_287),
.Y(n_333)
);

OR2x2_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_205),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_288),
.A2(n_301),
.B(n_302),
.Y(n_319)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_263),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_289),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_264),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_294),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_229),
.A2(n_182),
.B1(n_189),
.B2(n_220),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_252),
.B(n_246),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_191),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_293),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_261),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_265),
.Y(n_296)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

INVx13_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_236),
.B(n_204),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_298),
.Y(n_347)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_300),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_251),
.Y(n_300)
);

AND2x6_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_204),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_249),
.A2(n_221),
.B(n_209),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_255),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_303),
.B(n_306),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_249),
.B(n_216),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_304),
.A2(n_228),
.B(n_242),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_253),
.A2(n_206),
.B1(n_151),
.B2(n_171),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_173),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_307),
.B(n_309),
.Y(n_337)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_311),
.Y(n_351)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_267),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_232),
.B(n_212),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_238),
.B(n_248),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_317),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_285),
.B(n_256),
.C(n_259),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_322),
.B(n_324),
.C(n_336),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_226),
.C(n_235),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_288),
.A2(n_281),
.B1(n_306),
.B2(n_280),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_326),
.B(n_339),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_280),
.A2(n_251),
.B1(n_234),
.B2(n_250),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_335),
.A2(n_273),
.B1(n_272),
.B2(n_312),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_275),
.B(n_270),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_338),
.B(n_349),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_304),
.A2(n_250),
.B1(n_224),
.B2(n_233),
.Y(n_339)
);

AND2x2_ASAP7_75t_SL g341 ( 
.A(n_314),
.B(n_258),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_341),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_292),
.A2(n_271),
.B(n_233),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_345),
.B(n_353),
.Y(n_380)
);

OA22x2_ASAP7_75t_L g344 ( 
.A1(n_283),
.A2(n_305),
.B1(n_301),
.B2(n_277),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_295),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_292),
.A2(n_209),
.B(n_241),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_271),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_304),
.B(n_212),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_SL g359 ( 
.A(n_350),
.B(n_354),
.C(n_274),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_241),
.C(n_112),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_352),
.B(n_273),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_104),
.B(n_8),
.Y(n_353)
);

AOI32xp33_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_355),
.Y(n_388)
);

NOR2x1_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_308),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_363),
.Y(n_389)
);

INVx13_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_357),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_379),
.B(n_342),
.Y(n_393)
);

INVx13_ASAP7_75t_L g360 ( 
.A(n_332),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_361),
.Y(n_391)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_362),
.A2(n_344),
.B(n_346),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_321),
.A2(n_284),
.B1(n_296),
.B2(n_300),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_330),
.B(n_284),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_365),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_330),
.B(n_287),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_318),
.B(n_303),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_381),
.Y(n_403)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_332),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_372),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_294),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_378),
.Y(n_400)
);

OAI22x1_ASAP7_75t_L g370 ( 
.A1(n_341),
.A2(n_353),
.B1(n_342),
.B2(n_319),
.Y(n_370)
);

A2O1A1Ixp33_ASAP7_75t_SL g409 ( 
.A1(n_370),
.A2(n_341),
.B(n_344),
.C(n_350),
.Y(n_409)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_351),
.Y(n_371)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_371),
.Y(n_399)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_351),
.Y(n_374)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_347),
.B(n_307),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_375),
.B(n_320),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_337),
.B(n_311),
.Y(n_376)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_376),
.Y(n_411)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_333),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_377),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_328),
.Y(n_378)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_289),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_328),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_382),
.B(n_383),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_334),
.B(n_276),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_337),
.B(n_310),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_386),
.B(n_323),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_393),
.B(n_410),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_373),
.A2(n_345),
.B(n_318),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_416),
.B(n_380),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_405),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_368),
.B(n_349),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_402),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_338),
.Y(n_402)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_362),
.A2(n_317),
.B1(n_352),
.B2(n_344),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_375),
.B(n_297),
.Y(n_406)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_406),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_336),
.C(n_322),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_407),
.B(n_358),
.C(n_385),
.Y(n_425)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_370),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_L g410 ( 
.A(n_370),
.B(n_329),
.C(n_320),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_387),
.B(n_324),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_414),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_413),
.B(n_415),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_371),
.B(n_343),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_363),
.B(n_335),
.Y(n_416)
);

XNOR2x1_ASAP7_75t_L g449 ( 
.A(n_417),
.B(n_389),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_400),
.A2(n_384),
.B1(n_358),
.B2(n_359),
.Y(n_418)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_404),
.B(n_369),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_421),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_395),
.B(n_364),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_430),
.C(n_441),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_400),
.A2(n_366),
.B1(n_365),
.B2(n_385),
.Y(n_426)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_426),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_374),
.B1(n_382),
.B2(n_378),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_428),
.A2(n_429),
.B1(n_433),
.B2(n_438),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_403),
.A2(n_355),
.B1(n_377),
.B2(n_361),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_407),
.C(n_398),
.Y(n_430)
);

CKINVDCx16_ASAP7_75t_R g431 ( 
.A(n_388),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_431),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_392),
.B(n_357),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_432),
.A2(n_391),
.B(n_388),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_380),
.B1(n_316),
.B2(n_376),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_402),
.B(n_386),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_436),
.B(n_409),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_414),
.B(n_346),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_440),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_379),
.B1(n_331),
.B2(n_333),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_439),
.A2(n_391),
.B1(n_401),
.B2(n_397),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_411),
.B(n_356),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_408),
.C(n_399),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_437),
.A2(n_405),
.B1(n_416),
.B2(n_399),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_442),
.A2(n_454),
.B1(n_327),
.B2(n_325),
.Y(n_472)
);

NOR2xp67_ASAP7_75t_SL g447 ( 
.A(n_417),
.B(n_379),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_447),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_430),
.B(n_419),
.C(n_425),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_456),
.C(n_457),
.Y(n_466)
);

A2O1A1Ixp33_ASAP7_75t_SL g474 ( 
.A1(n_449),
.A2(n_367),
.B(n_360),
.C(n_327),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_450),
.B(n_451),
.Y(n_476)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_417),
.B(n_409),
.C(n_411),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_417),
.A2(n_416),
.B1(n_408),
.B2(n_356),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g455 ( 
.A(n_417),
.B(n_389),
.CI(n_409),
.CON(n_455),
.SN(n_455)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_455),
.B(n_381),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_419),
.B(n_396),
.C(n_390),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_397),
.Y(n_457)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_458),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_461),
.A2(n_422),
.B1(n_452),
.B2(n_459),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_462),
.B(n_472),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_L g463 ( 
.A1(n_446),
.A2(n_440),
.B1(n_434),
.B2(n_441),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_474),
.Y(n_481)
);

A2O1A1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_460),
.A2(n_427),
.B(n_434),
.C(n_438),
.Y(n_464)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_464),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_455),
.B(n_435),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g483 ( 
.A(n_465),
.Y(n_483)
);

AO221x1_ASAP7_75t_L g467 ( 
.A1(n_453),
.A2(n_331),
.B1(n_423),
.B2(n_357),
.C(n_367),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_467),
.A2(n_454),
.B(n_442),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_424),
.C(n_436),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_468),
.B(n_450),
.C(n_457),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_444),
.B(n_325),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_470),
.B(n_475),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_471),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_309),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_451),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_477),
.B(n_455),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_SL g478 ( 
.A(n_469),
.B(n_456),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_485),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_473),
.A2(n_460),
.B(n_448),
.Y(n_480)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_482),
.B(n_488),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_466),
.B(n_443),
.C(n_449),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_490),
.C(n_468),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_466),
.B(n_443),
.C(n_299),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_484),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_476),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_484),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_479),
.A2(n_465),
.B1(n_473),
.B2(n_463),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_494),
.B(n_497),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_483),
.B(n_464),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_490),
.B(n_474),
.C(n_312),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_498),
.B(n_499),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_486),
.B(n_474),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_360),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_7),
.C(n_9),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_487),
.B1(n_481),
.B2(n_482),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_504),
.A2(n_481),
.B1(n_474),
.B2(n_493),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_498),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_508),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_505),
.A2(n_496),
.B1(n_492),
.B2(n_491),
.Y(n_508)
);

OAI31xp67_ASAP7_75t_L g512 ( 
.A1(n_509),
.A2(n_510),
.A3(n_503),
.B(n_501),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_512),
.A2(n_510),
.B1(n_507),
.B2(n_502),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_513),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_511),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_506),
.C(n_9),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_7),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_11),
.B(n_12),
.Y(n_518)
);


endmodule