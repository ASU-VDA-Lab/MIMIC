module fake_aes_6947_n_556 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_556);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_556;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_69;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_70;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_68;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g68 ( .A(n_28), .Y(n_68) );
INVx2_ASAP7_75t_L g69 ( .A(n_65), .Y(n_69) );
INVx1_ASAP7_75t_L g70 ( .A(n_67), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_16), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_57), .Y(n_72) );
INVx1_ASAP7_75t_L g73 ( .A(n_60), .Y(n_73) );
INVxp67_ASAP7_75t_SL g74 ( .A(n_50), .Y(n_74) );
INVxp67_ASAP7_75t_L g75 ( .A(n_43), .Y(n_75) );
CKINVDCx20_ASAP7_75t_R g76 ( .A(n_56), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_0), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_62), .Y(n_78) );
INVx2_ASAP7_75t_L g79 ( .A(n_29), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_66), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_33), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_15), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_20), .Y(n_84) );
INVxp33_ASAP7_75t_L g85 ( .A(n_45), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_17), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_12), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_14), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_63), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_16), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_49), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_44), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_4), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_48), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_22), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g97 ( .A(n_11), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_6), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_5), .Y(n_99) );
INVxp67_ASAP7_75t_SL g100 ( .A(n_21), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_52), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_35), .Y(n_104) );
INVxp67_ASAP7_75t_SL g105 ( .A(n_37), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_10), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_34), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_30), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_53), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_24), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
CKINVDCx14_ASAP7_75t_R g112 ( .A(n_31), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
INVx2_ASAP7_75t_SL g114 ( .A(n_12), .Y(n_114) );
INVxp33_ASAP7_75t_L g115 ( .A(n_25), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_10), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_114), .B(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_70), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_98), .B(n_1), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_90), .B(n_1), .Y(n_121) );
BUFx6f_ASAP7_75t_L g122 ( .A(n_91), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_76), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_69), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_70), .Y(n_125) );
BUFx10_ASAP7_75t_L g126 ( .A(n_78), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_97), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_72), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_84), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_72), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_94), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_111), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_114), .B(n_2), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_85), .B(n_3), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_73), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_113), .B(n_3), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_112), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_79), .B(n_4), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_73), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_80), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g141 ( .A(n_91), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_80), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_108), .B(n_5), .Y(n_144) );
NOR2xp33_ASAP7_75t_R g145 ( .A(n_89), .B(n_36), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_108), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_81), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_81), .B(n_6), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_71), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_93), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_115), .B(n_90), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_68), .Y(n_152) );
AND2x6_ASAP7_75t_L g153 ( .A(n_93), .B(n_38), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_71), .B(n_7), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_77), .B(n_8), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_95), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_77), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_95), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_92), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_154), .A2(n_116), .B1(n_99), .B2(n_82), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_146), .Y(n_164) );
INVx3_ASAP7_75t_L g165 ( .A(n_154), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_146), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_154), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_153), .Y(n_169) );
AND2x4_ASAP7_75t_L g170 ( .A(n_151), .B(n_116), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_146), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_126), .B(n_75), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_146), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_119), .A2(n_110), .B(n_96), .C(n_101), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_154), .Y(n_176) );
CKINVDCx8_ASAP7_75t_R g177 ( .A(n_123), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_121), .B(n_110), .Y(n_178) );
AND2x2_ASAP7_75t_L g179 ( .A(n_151), .B(n_87), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
NAND2x1p5_ASAP7_75t_L g181 ( .A(n_121), .B(n_103), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_122), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_121), .B(n_82), .Y(n_183) );
NAND2x1p5_ASAP7_75t_L g184 ( .A(n_121), .B(n_101), .Y(n_184) );
AO22x2_ASAP7_75t_L g185 ( .A1(n_119), .A2(n_104), .B1(n_102), .B2(n_103), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_122), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_156), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_122), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_159), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_122), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_159), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_117), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_127), .Y(n_194) );
BUFx4f_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_157), .B(n_83), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_125), .B(n_83), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_122), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_126), .B(n_109), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_125), .B(n_86), .Y(n_201) );
CKINVDCx16_ASAP7_75t_R g202 ( .A(n_137), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_117), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_122), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_128), .B(n_86), .Y(n_205) );
NOR2x1p5_ASAP7_75t_L g206 ( .A(n_129), .B(n_87), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_126), .B(n_102), .Y(n_207) );
BUFx3_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_128), .B(n_88), .Y(n_209) );
AND2x4_ASAP7_75t_L g210 ( .A(n_130), .B(n_88), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_126), .B(n_104), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_117), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_124), .Y(n_213) );
CKINVDCx8_ASAP7_75t_R g214 ( .A(n_132), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_124), .Y(n_215) );
INVx3_ASAP7_75t_L g216 ( .A(n_142), .Y(n_216) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_155), .B(n_106), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_124), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_147), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
NOR2x1p5_ASAP7_75t_L g222 ( .A(n_152), .B(n_106), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_147), .Y(n_223) );
CKINVDCx16_ASAP7_75t_R g224 ( .A(n_194), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_218), .B(n_134), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_174), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_217), .B(n_134), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_221), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_217), .A2(n_153), .B1(n_147), .B2(n_155), .Y(n_229) );
INVx4_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_174), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_207), .B(n_139), .Y(n_232) );
NOR3xp33_ASAP7_75t_SL g233 ( .A(n_202), .B(n_160), .C(n_120), .Y(n_233) );
INVx5_ASAP7_75t_L g234 ( .A(n_221), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
INVx3_ASAP7_75t_SL g236 ( .A(n_196), .Y(n_236) );
INVx3_ASAP7_75t_L g237 ( .A(n_216), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_178), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_168), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_178), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_211), .B(n_139), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_169), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_178), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_181), .Y(n_244) );
NAND2x1_ASAP7_75t_L g245 ( .A(n_165), .B(n_150), .Y(n_245) );
AND2x4_ASAP7_75t_L g246 ( .A(n_196), .B(n_141), .Y(n_246) );
BUFx2_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_180), .Y(n_248) );
INVx5_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_172), .B(n_135), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_185), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_187), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_205), .B(n_143), .Y(n_253) );
BUFx10_ASAP7_75t_L g254 ( .A(n_222), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_183), .B(n_133), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_218), .B(n_150), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_217), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_181), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_200), .B(n_135), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_181), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_197), .Y(n_261) );
BUFx2_ASAP7_75t_L g262 ( .A(n_185), .Y(n_262) );
NOR2xp33_ASAP7_75t_R g263 ( .A(n_214), .B(n_149), .Y(n_263) );
BUFx3_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_184), .Y(n_265) );
BUFx2_ASAP7_75t_L g266 ( .A(n_185), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_222), .A2(n_118), .B1(n_143), .B2(n_140), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_184), .Y(n_268) );
NOR3xp33_ASAP7_75t_SL g269 ( .A(n_202), .B(n_136), .C(n_148), .Y(n_269) );
AO22x1_ASAP7_75t_L g270 ( .A1(n_183), .A2(n_74), .B1(n_100), .B2(n_105), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g271 ( .A1(n_184), .A2(n_140), .B1(n_130), .B2(n_144), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_170), .B(n_138), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_187), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_216), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_189), .Y(n_275) );
AND2x4_ASAP7_75t_L g276 ( .A(n_183), .B(n_158), .Y(n_276) );
A2O1A1Ixp33_ASAP7_75t_L g277 ( .A1(n_165), .A2(n_158), .B(n_142), .C(n_99), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_214), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_170), .B(n_142), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_179), .B(n_107), .Y(n_280) );
NOR2xp33_ASAP7_75t_R g281 ( .A(n_177), .B(n_40), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_179), .B(n_145), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_195), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_256), .A2(n_195), .B(n_165), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_258), .B(n_206), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_236), .B(n_167), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_276), .Y(n_287) );
BUFx12f_ASAP7_75t_L g288 ( .A(n_239), .Y(n_288) );
AO22x1_ASAP7_75t_L g289 ( .A1(n_239), .A2(n_177), .B1(n_205), .B2(n_167), .Y(n_289) );
O2A1O1Ixp5_ASAP7_75t_SL g290 ( .A1(n_271), .A2(n_166), .B(n_171), .C(n_219), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_236), .B(n_167), .Y(n_291) );
INVx2_ASAP7_75t_SL g292 ( .A(n_258), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_251), .A2(n_266), .B1(n_262), .B2(n_260), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_246), .B(n_206), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_260), .B(n_205), .Y(n_295) );
BUFx6f_ASAP7_75t_L g296 ( .A(n_228), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_226), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_230), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_238), .B(n_198), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_247), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_226), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_277), .A2(n_176), .B(n_189), .C(n_191), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_SL g304 ( .A1(n_229), .A2(n_176), .B(n_199), .C(n_188), .Y(n_304) );
BUFx4f_ASAP7_75t_SL g305 ( .A(n_246), .Y(n_305) );
NOR3xp33_ASAP7_75t_L g306 ( .A(n_224), .B(n_175), .C(n_176), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
BUFx12f_ASAP7_75t_L g308 ( .A(n_254), .Y(n_308) );
NOR2x1_ASAP7_75t_SL g309 ( .A(n_240), .B(n_192), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_251), .A2(n_185), .B1(n_198), .B2(n_201), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_246), .B(n_198), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_230), .Y(n_312) );
INVx4_ASAP7_75t_L g313 ( .A(n_262), .Y(n_313) );
BUFx8_ASAP7_75t_SL g314 ( .A(n_257), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_253), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_230), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_231), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_266), .A2(n_201), .B1(n_198), .B2(n_209), .Y(n_318) );
OAI21xp33_ASAP7_75t_L g319 ( .A1(n_272), .A2(n_162), .B(n_209), .Y(n_319) );
BUFx4_ASAP7_75t_SL g320 ( .A(n_243), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_256), .A2(n_195), .B(n_220), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_255), .B(n_210), .Y(n_322) );
BUFx3_ASAP7_75t_L g323 ( .A(n_244), .Y(n_323) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_265), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_268), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_225), .A2(n_220), .B(n_223), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
O2A1O1Ixp33_ASAP7_75t_SL g328 ( .A1(n_277), .A2(n_171), .B(n_166), .C(n_191), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_234), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_228), .Y(n_330) );
BUFx6f_ASAP7_75t_L g331 ( .A(n_228), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_228), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_235), .Y(n_333) );
INVx3_ASAP7_75t_L g334 ( .A(n_237), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_305), .A2(n_257), .B1(n_227), .B2(n_255), .Y(n_335) );
OAI22xp5_ASAP7_75t_L g336 ( .A1(n_310), .A2(n_255), .B1(n_241), .B2(n_232), .Y(n_336) );
INVx2_ASAP7_75t_SL g337 ( .A(n_323), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_311), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_318), .A2(n_280), .B1(n_273), .B2(n_252), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_323), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_322), .A2(n_280), .B1(n_273), .B2(n_252), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_329), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_300), .B(n_283), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_294), .B(n_278), .Y(n_344) );
INVx6_ASAP7_75t_L g345 ( .A(n_308), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_329), .Y(n_346) );
BUFx8_ASAP7_75t_L g347 ( .A(n_288), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_315), .B(n_235), .Y(n_348) );
CKINVDCx5p33_ASAP7_75t_R g349 ( .A(n_320), .Y(n_349) );
CKINVDCx5p33_ASAP7_75t_R g350 ( .A(n_288), .Y(n_350) );
O2A1O1Ixp33_ASAP7_75t_SL g351 ( .A1(n_304), .A2(n_192), .B(n_225), .C(n_203), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_300), .B(n_280), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_300), .B(n_282), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_324), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_285), .B(n_267), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_295), .B(n_270), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_306), .A2(n_282), .B1(n_263), .B2(n_279), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_325), .B(n_295), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_307), .Y(n_360) );
AND2x4_ASAP7_75t_L g361 ( .A(n_309), .B(n_283), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_290), .A2(n_326), .B(n_321), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_298), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_289), .B(n_248), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_295), .B(n_250), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_287), .Y(n_366) );
AOI221xp5_ASAP7_75t_L g367 ( .A1(n_319), .A2(n_269), .B1(n_233), .B2(n_259), .C(n_210), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_338), .B(n_285), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_336), .A2(n_313), .B1(n_293), .B2(n_333), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_341), .A2(n_313), .B1(n_327), .B2(n_292), .Y(n_370) );
AOI22xp33_ASAP7_75t_SL g371 ( .A1(n_347), .A2(n_313), .B1(n_281), .B2(n_285), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_348), .B(n_298), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_348), .Y(n_373) );
INVx3_ASAP7_75t_L g374 ( .A(n_342), .Y(n_374) );
OAI22xp5_ASAP7_75t_SL g375 ( .A1(n_357), .A2(n_308), .B1(n_314), .B2(n_292), .Y(n_375) );
AOI221xp5_ASAP7_75t_L g376 ( .A1(n_356), .A2(n_297), .B1(n_303), .B2(n_209), .C(n_210), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g377 ( .A1(n_339), .A2(n_210), .B1(n_209), .B2(n_201), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_363), .B(n_302), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_363), .Y(n_379) );
OAI211xp5_ASAP7_75t_SL g380 ( .A1(n_358), .A2(n_303), .B(n_212), .C(n_215), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_362), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_366), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_357), .A2(n_286), .B1(n_291), .B2(n_201), .Y(n_383) );
NAND2xp33_ASAP7_75t_SL g384 ( .A(n_337), .B(n_302), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_337), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g386 ( .A1(n_364), .A2(n_317), .B1(n_248), .B2(n_275), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_357), .B(n_317), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_357), .A2(n_286), .B1(n_291), .B2(n_334), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_354), .A2(n_328), .B1(n_203), .B2(n_193), .C(n_212), .Y(n_389) );
AOI21x1_ASAP7_75t_L g390 ( .A1(n_362), .A2(n_186), .B(n_182), .Y(n_390) );
AO21x2_ASAP7_75t_L g391 ( .A1(n_351), .A2(n_304), .B(n_328), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_353), .B(n_275), .Y(n_392) );
AND2x6_ASAP7_75t_SL g393 ( .A(n_347), .B(n_314), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g394 ( .A1(n_367), .A2(n_245), .B(n_193), .C(n_215), .Y(n_394) );
OAI211xp5_ASAP7_75t_SL g395 ( .A1(n_344), .A2(n_219), .B(n_213), .C(n_254), .Y(n_395) );
AOI222xp33_ASAP7_75t_L g396 ( .A1(n_375), .A2(n_347), .B1(n_335), .B2(n_352), .C1(n_360), .C2(n_355), .Y(n_396) );
AOI21x1_ASAP7_75t_L g397 ( .A1(n_390), .A2(n_364), .B(n_190), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_372), .B(n_340), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_375), .B(n_350), .Y(n_399) );
OAI211xp5_ASAP7_75t_SL g400 ( .A1(n_368), .A2(n_359), .B(n_365), .C(n_340), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
OR2x6_ASAP7_75t_L g402 ( .A(n_386), .B(n_340), .Y(n_402) );
BUFx3_ASAP7_75t_L g403 ( .A(n_372), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_390), .A2(n_351), .B(n_284), .Y(n_404) );
INVx4_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_377), .A2(n_383), .B1(n_386), .B2(n_371), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_378), .B(n_342), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_376), .A2(n_343), .B1(n_342), .B2(n_346), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_382), .B(n_350), .Y(n_409) );
INVxp67_ASAP7_75t_SL g410 ( .A(n_379), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_373), .B(n_346), .Y(n_411) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_388), .A2(n_345), .B1(n_349), .B2(n_346), .C(n_334), .Y(n_412) );
AND2x4_ASAP7_75t_L g413 ( .A(n_387), .B(n_361), .Y(n_413) );
OAI21xp33_ASAP7_75t_L g414 ( .A1(n_377), .A2(n_361), .B(n_349), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_387), .B(n_361), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_373), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_380), .A2(n_343), .B1(n_345), .B2(n_312), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_382), .Y(n_418) );
BUFx3_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_395), .A2(n_343), .B1(n_213), .B2(n_237), .C(n_274), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_381), .Y(n_421) );
CKINVDCx8_ASAP7_75t_R g422 ( .A(n_393), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_374), .B(n_9), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_381), .Y(n_424) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_369), .A2(n_274), .B1(n_299), .B2(n_312), .C(n_316), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_381), .Y(n_426) );
CKINVDCx20_ASAP7_75t_R g427 ( .A(n_393), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_414), .B(n_384), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_401), .B(n_391), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_421), .Y(n_430) );
AND2x4_ASAP7_75t_L g431 ( .A(n_424), .B(n_374), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_418), .B(n_374), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_410), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_424), .Y(n_434) );
OAI31xp33_ASAP7_75t_L g435 ( .A1(n_406), .A2(n_370), .A3(n_394), .B(n_385), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_426), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_401), .B(n_391), .Y(n_437) );
OAI33xp33_ASAP7_75t_L g438 ( .A1(n_400), .A2(n_392), .A3(n_11), .B1(n_13), .B2(n_14), .B3(n_15), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_416), .B(n_389), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_405), .Y(n_440) );
NAND4xp25_ASAP7_75t_SL g441 ( .A(n_396), .B(n_9), .C(n_13), .D(n_17), .Y(n_441) );
BUFx3_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
INVx1_ASAP7_75t_SL g443 ( .A(n_419), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_403), .B(n_18), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_397), .Y(n_445) );
AND2x4_ASAP7_75t_L g446 ( .A(n_402), .B(n_330), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_398), .B(n_19), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_398), .B(n_19), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_402), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_397), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_414), .A2(n_316), .B1(n_312), .B2(n_299), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_419), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
AOI31xp33_ASAP7_75t_L g456 ( .A1(n_399), .A2(n_254), .A3(n_223), .B(n_27), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_402), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_409), .B(n_329), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_402), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_407), .B(n_186), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_408), .B(n_199), .C(n_182), .D(n_188), .Y(n_461) );
AOI211xp5_ASAP7_75t_L g462 ( .A1(n_412), .A2(n_204), .B(n_161), .C(n_173), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_411), .B(n_204), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_413), .B(n_23), .Y(n_464) );
INVx3_ASAP7_75t_SL g465 ( .A(n_413), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_442), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_441), .B(n_422), .Y(n_467) );
OAI211xp5_ASAP7_75t_L g468 ( .A1(n_435), .A2(n_422), .B(n_427), .C(n_417), .Y(n_468) );
NOR2xp33_ASAP7_75t_SL g469 ( .A(n_444), .B(n_405), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_457), .B(n_405), .Y(n_470) );
OAI21xp33_ASAP7_75t_L g471 ( .A1(n_441), .A2(n_423), .B(n_411), .Y(n_471) );
OAI211xp5_ASAP7_75t_SL g472 ( .A1(n_435), .A2(n_420), .B(n_425), .C(n_161), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_465), .B(n_415), .Y(n_473) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_456), .B(n_413), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_444), .B(n_330), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_444), .B(n_26), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_447), .B(n_173), .Y(n_477) );
BUFx2_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g479 ( .A(n_442), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_447), .B(n_32), .Y(n_480) );
NOR3xp33_ASAP7_75t_L g481 ( .A(n_456), .B(n_164), .C(n_163), .Y(n_481) );
NAND2x1_ASAP7_75t_L g482 ( .A(n_440), .B(n_332), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_430), .Y(n_483) );
NOR2xp33_ASAP7_75t_R g484 ( .A(n_440), .B(n_330), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_440), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_448), .B(n_39), .Y(n_486) );
INVx5_ASAP7_75t_L g487 ( .A(n_440), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_448), .B(n_41), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_451), .A2(n_330), .B1(n_331), .B2(n_332), .Y(n_489) );
NOR2xp33_ASAP7_75t_R g490 ( .A(n_464), .B(n_47), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_438), .A2(n_332), .B1(n_331), .B2(n_296), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_458), .B(n_51), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_479), .B(n_433), .Y(n_493) );
AOI32xp33_ASAP7_75t_L g494 ( .A1(n_467), .A2(n_464), .A3(n_449), .B1(n_462), .B2(n_443), .Y(n_494) );
AND2x4_ASAP7_75t_SL g495 ( .A(n_473), .B(n_446), .Y(n_495) );
AOI32xp33_ASAP7_75t_L g496 ( .A1(n_467), .A2(n_453), .A3(n_443), .B1(n_428), .B2(n_446), .Y(n_496) );
INVxp33_ASAP7_75t_L g497 ( .A(n_490), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_L g498 ( .A1(n_481), .A2(n_439), .B(n_463), .C(n_432), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_474), .A2(n_446), .B(n_433), .C(n_459), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_483), .B(n_429), .Y(n_500) );
XNOR2x2_ASAP7_75t_L g501 ( .A(n_474), .B(n_432), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_484), .Y(n_502) );
OAI321xp33_ASAP7_75t_L g503 ( .A1(n_468), .A2(n_459), .A3(n_461), .B1(n_460), .B2(n_437), .C(n_439), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g504 ( .A1(n_481), .A2(n_460), .B1(n_437), .B2(n_461), .Y(n_504) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_492), .B(n_460), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_469), .A2(n_431), .B1(n_463), .B2(n_436), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_478), .B(n_434), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_475), .A2(n_436), .B1(n_431), .B2(n_450), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_471), .A2(n_455), .B1(n_454), .B2(n_452), .Y(n_509) );
AOI22xp5_ASAP7_75t_SL g510 ( .A1(n_466), .A2(n_445), .B1(n_454), .B2(n_452), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_487), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_470), .B(n_54), .Y(n_512) );
OAI211xp5_ASAP7_75t_SL g513 ( .A1(n_477), .A2(n_58), .B(n_59), .C(n_61), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_485), .Y(n_515) );
NOR4xp25_ASAP7_75t_SL g516 ( .A(n_503), .B(n_490), .C(n_487), .D(n_472), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_500), .B(n_470), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_493), .Y(n_518) );
NOR4xp25_ASAP7_75t_SL g519 ( .A(n_499), .B(n_487), .C(n_482), .D(n_480), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_498), .A2(n_486), .B(n_488), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g521 ( .A1(n_497), .A2(n_487), .B1(n_476), .B2(n_491), .Y(n_521) );
HB1xp67_ASAP7_75t_L g522 ( .A(n_515), .Y(n_522) );
AND3x2_ASAP7_75t_L g523 ( .A(n_511), .B(n_489), .C(n_64), .Y(n_523) );
XNOR2xp5_ASAP7_75t_L g524 ( .A(n_501), .B(n_264), .Y(n_524) );
NAND4xp25_ASAP7_75t_L g525 ( .A(n_496), .B(n_242), .C(n_234), .D(n_249), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_502), .B(n_296), .Y(n_526) );
OAI211xp5_ASAP7_75t_L g527 ( .A1(n_494), .A2(n_296), .B(n_234), .C(n_249), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_525), .A2(n_510), .B(n_508), .Y(n_528) );
OAI31xp33_ASAP7_75t_L g529 ( .A1(n_527), .A2(n_505), .A3(n_513), .B(n_495), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_518), .A2(n_504), .B1(n_506), .B2(n_514), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_520), .A2(n_509), .B(n_512), .Y(n_531) );
NAND2x1p5_ASAP7_75t_L g532 ( .A(n_518), .B(n_507), .Y(n_532) );
INVx1_ASAP7_75t_SL g533 ( .A(n_522), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_519), .A2(n_249), .B(n_261), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_531), .B(n_516), .C(n_524), .Y(n_535) );
AOI31xp33_ASAP7_75t_L g536 ( .A1(n_532), .A2(n_521), .A3(n_516), .B(n_517), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_533), .Y(n_537) );
AND3x2_ASAP7_75t_L g538 ( .A(n_529), .B(n_523), .C(n_526), .Y(n_538) );
BUFx2_ASAP7_75t_L g539 ( .A(n_532), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_534), .B(n_529), .C(n_467), .D(n_528), .Y(n_540) );
AND4x1_ASAP7_75t_L g541 ( .A(n_529), .B(n_528), .C(n_467), .D(n_531), .Y(n_541) );
AOI211xp5_ASAP7_75t_L g542 ( .A1(n_530), .A2(n_528), .B(n_531), .C(n_525), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_537), .Y(n_543) );
INVx1_ASAP7_75t_SL g544 ( .A(n_539), .Y(n_544) );
XNOR2xp5_ASAP7_75t_L g545 ( .A(n_541), .B(n_538), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_538), .Y(n_546) );
OR3x2_ASAP7_75t_L g547 ( .A(n_540), .B(n_542), .C(n_536), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_543), .Y(n_548) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_544), .Y(n_549) );
NOR2x1_ASAP7_75t_L g550 ( .A(n_546), .B(n_535), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_549), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_548), .Y(n_552) );
INVx3_ASAP7_75t_SL g553 ( .A(n_551), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_552), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_553), .A2(n_547), .B1(n_545), .B2(n_550), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_544), .B(n_554), .Y(n_556) );
endmodule