module fake_jpeg_26080_n_307 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_307);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_10;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_24),
.A2(n_12),
.B1(n_11),
.B2(n_18),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_32),
.B1(n_30),
.B2(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_20),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_20),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_52),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_46),
.B(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx2_ASAP7_75t_SL g63 ( 
.A(n_49),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_42),
.A2(n_29),
.B1(n_24),
.B2(n_32),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_53),
.B(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_33),
.Y(n_52)
);

AOI22x1_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_12),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_11),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_40),
.B2(n_35),
.Y(n_70)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_32),
.B1(n_23),
.B2(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_45),
.Y(n_90)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_76),
.B1(n_77),
.B2(n_54),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_38),
.B(n_26),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_26),
.C(n_25),
.Y(n_100)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_23),
.B(n_29),
.Y(n_73)
);

AOI32xp33_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_40),
.A3(n_57),
.B1(n_25),
.B2(n_26),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_62),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_50),
.A2(n_35),
.B1(n_36),
.B2(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_81),
.B(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_84),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_80),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_83),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_85),
.B(n_90),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_54),
.B1(n_61),
.B2(n_43),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_87),
.A2(n_98),
.B1(n_75),
.B2(n_43),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_72),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_103),
.B(n_25),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_79),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_91),
.B(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_97),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_100),
.Y(n_120)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_71),
.Y(n_99)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_26),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_94),
.A2(n_98),
.B1(n_100),
.B2(n_77),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_128),
.B1(n_96),
.B2(n_23),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_67),
.B1(n_64),
.B2(n_49),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_107),
.A2(n_115),
.B1(n_126),
.B2(n_75),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_103),
.B(n_98),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_111),
.A2(n_0),
.B(n_1),
.Y(n_137)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_114),
.B(n_28),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_67),
.B1(n_64),
.B2(n_56),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_25),
.C(n_69),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_129),
.C(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_78),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_18),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_88),
.A2(n_75),
.B1(n_76),
.B2(n_43),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_27),
.C(n_78),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_27),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_27),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_135),
.Y(n_169)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_134),
.A2(n_84),
.A3(n_101),
.B1(n_102),
.B2(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_136),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_157),
.B(n_162),
.Y(n_172)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_141),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_109),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_143),
.A2(n_151),
.B1(n_156),
.B2(n_135),
.Y(n_178)
);

NAND3xp33_ASAP7_75t_L g144 ( 
.A(n_104),
.B(n_0),
.C(n_1),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_158),
.C(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_126),
.B1(n_123),
.B2(n_127),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_145),
.A2(n_17),
.B1(n_15),
.B2(n_22),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_147),
.A2(n_150),
.B1(n_108),
.B2(n_112),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_106),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_148),
.Y(n_177)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_153),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_105),
.A2(n_96),
.B1(n_65),
.B2(n_51),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_111),
.A2(n_51),
.B1(n_10),
.B2(n_13),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_110),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_154),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_118),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_155),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_127),
.A2(n_13),
.B1(n_17),
.B2(n_15),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_125),
.B(n_31),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_125),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_120),
.B(n_28),
.C(n_13),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_116),
.C(n_117),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_107),
.B(n_31),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_28),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_16),
.B(n_21),
.Y(n_197)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_R g171 ( 
.A(n_157),
.B(n_124),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_171),
.A2(n_146),
.B(n_162),
.Y(n_200)
);

OA21x2_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_142),
.B(n_137),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_1),
.B(n_3),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_161),
.B1(n_160),
.B2(n_153),
.Y(n_201)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_159),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_120),
.B1(n_132),
.B2(n_113),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_180),
.A2(n_184),
.B1(n_194),
.B2(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_156),
.C(n_139),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_182),
.A2(n_190),
.B1(n_195),
.B2(n_162),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_165),
.A2(n_104),
.B1(n_108),
.B2(n_17),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_28),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_189),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_152),
.B(n_31),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_187),
.B(n_21),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_22),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_140),
.A2(n_16),
.B1(n_21),
.B2(n_19),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_147),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_196),
.B(n_172),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_142),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_200),
.A2(n_212),
.B(n_197),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_201),
.A2(n_202),
.B1(n_206),
.B2(n_219),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_149),
.B1(n_151),
.B2(n_146),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_182),
.B1(n_192),
.B2(n_175),
.Y(n_234)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_136),
.B1(n_168),
.B2(n_167),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_181),
.C(n_187),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_188),
.A2(n_138),
.B1(n_141),
.B2(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_213),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_138),
.Y(n_211)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_214),
.B(n_216),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_0),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_220),
.B(n_222),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_179),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_217),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_176),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_176),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_223),
.A2(n_191),
.B(n_193),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_225),
.A2(n_215),
.B(n_200),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_232),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_194),
.CI(n_178),
.CON(n_228),
.SN(n_228)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_228),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_186),
.C(n_189),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_239),
.C(n_240),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_234),
.A2(n_238),
.B1(n_242),
.B2(n_215),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_202),
.A2(n_195),
.B1(n_179),
.B2(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_21),
.C(n_4),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_3),
.C(n_4),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_205),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_206),
.Y(n_244)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_244),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_221),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_207),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_252),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_235),
.Y(n_264)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_225),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_254),
.B(n_223),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_256),
.B(n_257),
.Y(n_270)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_258),
.B(n_222),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_230),
.B1(n_250),
.B2(n_251),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_271),
.B1(n_266),
.B2(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_238),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_234),
.C(n_235),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_265),
.C(n_269),
.Y(n_280)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_253),
.C(n_255),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_232),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_268),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_210),
.C(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_274),
.A2(n_279),
.B1(n_257),
.B2(n_6),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_237),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_277),
.B(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_236),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_227),
.B1(n_236),
.B2(n_229),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_5),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_204),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_203),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_272),
.A2(n_249),
.B1(n_268),
.B2(n_221),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_285),
.B1(n_290),
.B2(n_291),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_228),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_288),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_280),
.B(n_237),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_289),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_284),
.C2(n_292),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_282),
.B(n_5),
.C(n_6),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_292),
.B(n_8),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_286),
.A2(n_276),
.B1(n_7),
.B2(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_276),
.B(n_7),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_296),
.B(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_9),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_300),
.A2(n_301),
.B(n_9),
.Y(n_302)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_299),
.B(n_9),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_305),
.A2(n_293),
.B(n_298),
.Y(n_306)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_306),
.A2(n_294),
.B(n_9),
.Y(n_307)
);


endmodule