module real_jpeg_11142_n_7 (n_5, n_4, n_36, n_0, n_39, n_37, n_40, n_1, n_41, n_2, n_38, n_6, n_3, n_7);

input n_5;
input n_4;
input n_36;
input n_0;
input n_39;
input n_37;
input n_40;
input n_1;
input n_41;
input n_2;
input n_38;
input n_6;
input n_3;

output n_7;

wire n_17;
wire n_8;
wire n_21;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_22;
wire n_18;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_15),
.C(n_31),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_26),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_17),
.C(n_25),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_4),
.B(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_5),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_5),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_14),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_27),
.C(n_28),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_21),
.C(n_22),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_36),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_37),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_38),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_39),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_40),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_41),
.Y(n_32)
);


endmodule