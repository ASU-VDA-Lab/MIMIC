module real_jpeg_31842_n_19 (n_17, n_8, n_0, n_2, n_10, n_726, n_9, n_12, n_6, n_11, n_14, n_725, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_726;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_725;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_715;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_696;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_666;
wire n_640;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_719;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_704;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_718;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_707;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_710;
wire n_110;
wire n_195;
wire n_703;
wire n_533;
wire n_592;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_689;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_697;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_716;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_712;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_714;
wire n_89;
wire n_407;
wire n_693;
wire n_721;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_711;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_698;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_635;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_686;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_699;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_720;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_708;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_723;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_701;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_695;
wire n_138;
wire n_662;
wire n_217;
wire n_709;
wire n_53;
wire n_717;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_702;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_602;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_706;
wire n_437;
wire n_268;
wire n_313;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_700;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_705;
wire n_530;
wire n_361;
wire n_694;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_722;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_690;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_713;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g253 ( 
.A(n_0),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_0),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_0),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_2),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_188),
.B1(n_189),
.B2(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_3),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_3),
.A2(n_188),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_3),
.A2(n_188),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_3),
.A2(n_188),
.B1(n_502),
.B2(n_504),
.Y(n_501)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_4),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_4),
.A2(n_51),
.B1(n_200),
.B2(n_203),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_4),
.A2(n_51),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_4),
.A2(n_51),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_5),
.A2(n_314),
.B1(n_315),
.B2(n_318),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_5),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_5),
.A2(n_105),
.B1(n_200),
.B2(n_314),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_5),
.A2(n_314),
.B1(n_552),
.B2(n_555),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_5),
.A2(n_314),
.B1(n_626),
.B2(n_630),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_6),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_6),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_6),
.A2(n_273),
.B1(n_405),
.B2(n_409),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_6),
.A2(n_273),
.B1(n_481),
.B2(n_483),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_6),
.A2(n_273),
.B1(n_580),
.B2(n_584),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_7),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g475 ( 
.A(n_7),
.Y(n_475)
);

NAND2xp33_ASAP7_75t_SL g509 ( 
.A(n_7),
.B(n_33),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_7),
.A2(n_475),
.B1(n_613),
.B2(n_614),
.Y(n_612)
);

OAI21xp33_ASAP7_75t_L g700 ( 
.A1(n_7),
.A2(n_248),
.B(n_635),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_8),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_9),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_11),
.A2(n_396),
.B1(n_397),
.B2(n_400),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_11),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_11),
.A2(n_396),
.B1(n_488),
.B2(n_492),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_11),
.A2(n_396),
.B1(n_604),
.B2(n_608),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_11),
.A2(n_396),
.B1(n_684),
.B2(n_687),
.Y(n_683)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_12),
.Y(n_141)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_12),
.Y(n_146)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_12),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_13),
.B(n_356),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_13),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_14),
.A2(n_112),
.B1(n_126),
.B2(n_130),
.Y(n_125)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_14),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_14),
.A2(n_130),
.B1(n_170),
.B2(n_175),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_14),
.A2(n_130),
.B1(n_222),
.B2(n_225),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_14),
.A2(n_130),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_15),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_15),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_16),
.A2(n_48),
.B1(n_59),
.B2(n_67),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_16),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_16),
.A2(n_67),
.B1(n_229),
.B2(n_232),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_16),
.A2(n_67),
.B1(n_288),
.B2(n_291),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_16),
.A2(n_67),
.B1(n_445),
.B2(n_447),
.Y(n_444)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_17),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_17),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_18),
.A2(n_103),
.B1(n_104),
.B2(n_110),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_18),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_18),
.A2(n_103),
.B1(n_158),
.B2(n_162),
.Y(n_157)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_18),
.A2(n_103),
.B1(n_142),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_18),
.A2(n_103),
.B1(n_349),
.B2(n_351),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_359),
.C(n_721),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_341),
.B1(n_357),
.B2(n_358),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI33xp33_ASAP7_75t_L g721 ( 
.A1(n_22),
.A2(n_361),
.A3(n_717),
.B1(n_722),
.B2(n_725),
.B3(n_726),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_207),
.B(n_339),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_23),
.B(n_718),
.Y(n_717)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_179),
.Y(n_25)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_26),
.B(n_179),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_164),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_27),
.B(n_165),
.C(n_168),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_84),
.C(n_131),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_29),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_47),
.B1(n_58),
.B2(n_68),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g345 ( 
.A1(n_31),
.A2(n_69),
.B1(n_346),
.B2(n_347),
.Y(n_345)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_32),
.A2(n_47),
.B1(n_68),
.B2(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_32),
.A2(n_58),
.B1(n_68),
.B2(n_187),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g265 ( 
.A(n_32),
.B(n_187),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_33),
.B(n_268),
.Y(n_311)
);

AO22x1_ASAP7_75t_SL g394 ( 
.A1(n_33),
.A2(n_70),
.B1(n_313),
.B2(n_395),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_33),
.B(n_395),
.Y(n_457)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_34),
.B(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_36),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_37),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_37),
.Y(n_324)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_41),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_41),
.Y(n_441)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_46),
.Y(n_412)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_50),
.Y(n_272)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_55),
.Y(n_178)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_55),
.Y(n_191)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_66),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_66),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_70),
.B(n_268),
.Y(n_267)
);

NAND2x1_ASAP7_75t_L g312 ( 
.A(n_70),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_70),
.B(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_74),
.B1(n_78),
.B2(n_81),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_81),
.Y(n_437)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_85),
.A2(n_133),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_101),
.B(n_114),
.Y(n_85)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_86),
.A2(n_402),
.B1(n_403),
.B2(n_413),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_86),
.A2(n_498),
.B(n_499),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_R g638 ( 
.A(n_86),
.B(n_475),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_87),
.Y(n_329)
);

AOI22x1_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_94),
.B2(n_97),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_90),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_91),
.A2(n_117),
.B1(n_120),
.B2(n_123),
.Y(n_116)
);

INVx5_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_93),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_99),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g558 ( 
.A(n_100),
.Y(n_558)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_109),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_109),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_109),
.Y(n_432)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_112),
.Y(n_613)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.Y(n_114)
);

OA21x2_ASAP7_75t_SL g165 ( 
.A1(n_115),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_115),
.A2(n_125),
.B1(n_166),
.B2(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_115),
.A2(n_166),
.B1(n_199),
.B2(n_228),
.Y(n_227)
);

AOI22x1_ASAP7_75t_L g320 ( 
.A1(n_115),
.A2(n_228),
.B1(n_321),
.B2(n_329),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_115),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_115),
.A2(n_166),
.B1(n_486),
.B2(n_487),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_115),
.B(n_404),
.Y(n_499)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_123),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g408 ( 
.A(n_129),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_129),
.Y(n_493)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_132),
.B(n_197),
.C(n_206),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_133),
.A2(n_184),
.B1(n_197),
.B2(n_198),
.Y(n_215)
);

OA21x2_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_147),
.B(n_157),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_134),
.A2(n_147),
.B1(n_157),
.B2(n_220),
.Y(n_219)
);

AO22x1_ASAP7_75t_L g478 ( 
.A1(n_134),
.A2(n_147),
.B1(n_479),
.B2(n_480),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_134),
.B(n_480),
.Y(n_559)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_134),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g261 ( 
.A(n_135),
.Y(n_261)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_139),
.B1(n_142),
.B2(n_145),
.Y(n_135)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_136),
.Y(n_446)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_137),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_138),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_138),
.Y(n_383)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_143),
.Y(n_634)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_144),
.Y(n_243)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_144),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_144),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_144),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_145),
.A2(n_150),
.B1(n_152),
.B2(n_154),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_146),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_147),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_147),
.A2(n_600),
.B1(n_601),
.B2(n_602),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_147),
.B(n_666),
.Y(n_665)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_148),
.A2(n_221),
.B1(n_255),
.B2(n_261),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_148),
.A2(n_255),
.B1(n_261),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_148),
.A2(n_261),
.B1(n_287),
.B2(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_148),
.A2(n_603),
.B1(n_640),
.B2(n_641),
.Y(n_639)
);

BUFx4f_ASAP7_75t_SL g650 ( 
.A(n_150),
.Y(n_650)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_156),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_156),
.Y(n_663)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_159),
.Y(n_484)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_160),
.Y(n_609)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_161),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_161),
.Y(n_576)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_163),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_169),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_174),
.Y(n_317)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_174),
.Y(n_352)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_174),
.Y(n_399)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_178),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_185),
.C(n_195),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_186),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_192),
.Y(n_474)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_202),
.Y(n_491)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_202),
.Y(n_614)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_277),
.B(n_337),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_209),
.B(n_720),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NOR2xp67_ASAP7_75t_L g338 ( 
.A(n_210),
.B(n_212),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.C(n_236),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g335 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_214),
.Y(n_336)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2x1_ASAP7_75t_L g332 ( 
.A(n_218),
.B(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_219),
.B(n_227),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g290 ( 
.A(n_226),
.Y(n_290)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_237),
.B(n_335),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_262),
.B(n_263),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_239),
.B(n_282),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_254),
.Y(n_239)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_240),
.B(n_264),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_240),
.A2(n_254),
.B1(n_262),
.B2(n_416),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_241),
.Y(n_303)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_242),
.Y(n_503)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_247),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_248),
.A2(n_294),
.B1(n_303),
.B2(n_304),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_248),
.A2(n_294),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_248),
.A2(n_444),
.B1(n_501),
.B2(n_506),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_248),
.A2(n_625),
.B(n_635),
.Y(n_624)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_249),
.A2(n_381),
.B1(n_443),
.B2(n_450),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_249),
.B(n_579),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_249),
.A2(n_678),
.B1(n_681),
.B2(n_682),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_252),
.Y(n_507)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_SL g637 ( 
.A(n_253),
.Y(n_637)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_254),
.Y(n_416)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_SL g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_261),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_267),
.B(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_334),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_279),
.B(n_334),
.Y(n_720)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.C(n_332),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_280),
.B(n_370),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_280),
.A2(n_281),
.B1(n_367),
.B2(n_370),
.Y(n_534)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_281),
.B(n_367),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_283),
.A2(n_284),
.B1(n_332),
.B2(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_309),
.B(n_330),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_285),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_293),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_286),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_293),
.B(n_464),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_296),
.Y(n_647)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_297),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_297),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_297),
.Y(n_659)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx2_ASAP7_75t_R g379 ( 
.A(n_307),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_308),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_319),
.Y(n_309)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_310),
.A2(n_319),
.B1(n_320),
.B2(n_331),
.Y(n_374)
);

NAND2x1_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_311),
.B(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_321),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_329),
.B(n_404),
.Y(n_461)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_332),
.Y(n_368)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

NAND3xp33_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_360),
.C(n_716),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_355),
.Y(n_341)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_342),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_353),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_353),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_348),
.Y(n_347)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI32xp33_ASAP7_75t_L g426 ( 
.A1(n_352),
.A2(n_427),
.A3(n_433),
.B1(n_436),
.B2(n_438),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_355),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_355),
.B(n_723),
.Y(n_722)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

NAND2x1_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_535),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_467),
.B(n_531),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_417),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_365),
.A2(n_532),
.B(n_533),
.Y(n_531)
);

NOR3xp33_ASAP7_75t_L g536 ( 
.A(n_365),
.B(n_417),
.C(n_537),
.Y(n_536)
);

AOI21x1_ASAP7_75t_L g365 ( 
.A1(n_366),
.A2(n_369),
.B(n_371),
.Y(n_365)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_367),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_371),
.B(n_534),
.Y(n_533)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_375),
.C(n_414),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_373),
.B(n_415),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_375),
.B(n_466),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_394),
.C(n_401),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_R g419 ( 
.A1(n_376),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_388),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_377),
.B(n_388),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

BUFx2_ASAP7_75t_SL g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_386),
.Y(n_586)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_387),
.Y(n_629)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_391),
.Y(n_554)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_393),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_401),
.Y(n_420)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_408),
.Y(n_574)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_413),
.A2(n_460),
.B(n_461),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g611 ( 
.A1(n_413),
.A2(n_461),
.B(n_612),
.Y(n_611)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_465),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_418),
.B(n_465),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_423),
.C(n_462),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_420),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_420),
.A2(n_421),
.B1(n_463),
.B2(n_530),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_422),
.B(n_424),
.Y(n_528)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_455),
.C(n_458),
.Y(n_424)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_442),
.Y(n_425)
);

XOR2x2_ASAP7_75t_L g494 ( 
.A(n_426),
.B(n_442),
.Y(n_494)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_431),
.Y(n_439)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_436),
.Y(n_476)
);

NAND2xp33_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

BUFx2_ASAP7_75t_SL g686 ( 
.A(n_449),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_450),
.B(n_588),
.Y(n_587)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx3_ASAP7_75t_SL g451 ( 
.A(n_452),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_455),
.A2(n_456),
.B1(n_458),
.B2(n_459),
.Y(n_520)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_460),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_463),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_523),
.C(n_526),
.Y(n_467)
);

OR2x2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_510),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_469),
.B(n_510),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_494),
.C(n_495),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_470),
.B(n_590),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_477),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_471),
.B(n_478),
.C(n_515),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_475),
.B(n_476),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_475),
.B(n_563),
.Y(n_562)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_475),
.B(n_573),
.C(n_575),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_475),
.B(n_663),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_475),
.A2(n_662),
.B(n_667),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_475),
.B(n_640),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_475),
.B(n_703),
.Y(n_702)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_485),
.Y(n_477)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_480),
.Y(n_641)
);

INVx3_ASAP7_75t_SL g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_487),
.Y(n_498)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_494),
.A2(n_495),
.B1(n_496),
.B2(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_494),
.Y(n_591)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_500),
.C(n_508),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_SL g545 ( 
.A(n_497),
.B(n_546),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_500),
.A2(n_508),
.B1(n_509),
.B2(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_500),
.Y(n_547)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_501),
.Y(n_588)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_511),
.A2(n_517),
.B(n_521),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_511),
.B(n_522),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_512),
.A2(n_513),
.B1(n_514),
.B2(n_516),
.Y(n_511)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_512),
.Y(n_516)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_514),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_516),
.Y(n_525)
);

MAJx2_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_524),
.C(n_525),
.Y(n_523)
);

INVx1_ASAP7_75t_SL g517 ( 
.A(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_518),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_523),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g526 ( 
.A(n_527),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_527),
.A2(n_538),
.B(n_539),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_529),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_540),
.Y(n_535)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_541),
.A2(n_592),
.B(n_714),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_589),
.Y(n_541)
);

INVxp67_ASAP7_75t_SL g542 ( 
.A(n_543),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_543),
.B(n_715),
.Y(n_714)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_548),
.C(n_560),
.Y(n_543)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g615 ( 
.A(n_545),
.B(n_616),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_548),
.A2(n_549),
.B1(n_560),
.B2(n_617),
.Y(n_616)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_550),
.A2(n_551),
.B(n_559),
.Y(n_549)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_551),
.Y(n_601)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_557),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_559),
.B(n_665),
.Y(n_664)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_577),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_577),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_562),
.A2(n_566),
.B(n_572),
.Y(n_561)
);

INVx4_ASAP7_75t_SL g563 ( 
.A(n_564),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_568),
.Y(n_566)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_575),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_587),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_SL g695 ( 
.A1(n_578),
.A2(n_683),
.B(n_696),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_579),
.B(n_636),
.Y(n_635)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_589),
.Y(n_715)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_593),
.A2(n_618),
.B(n_713),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_594),
.B(n_615),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g713 ( 
.A(n_594),
.B(n_615),
.Y(n_713)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_595),
.B(n_597),
.C(n_610),
.Y(n_594)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

XOR2xp5_ASAP7_75t_L g622 ( 
.A(n_599),
.B(n_611),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_603),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_619),
.B(n_673),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_620),
.A2(n_642),
.B(n_672),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_621),
.B(n_623),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_621),
.B(n_623),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_638),
.C(n_639),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_624),
.A2(n_669),
.B1(n_670),
.B2(n_671),
.Y(n_668)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_624),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_628),
.Y(n_687)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

XNOR2xp5_ASAP7_75t_L g669 ( 
.A(n_638),
.B(n_639),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_643),
.B(n_668),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_643),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_644),
.B(n_664),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g688 ( 
.A1(n_644),
.A2(n_664),
.B1(n_689),
.B2(n_690),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_644),
.Y(n_689)
);

AO221x1_ASAP7_75t_L g709 ( 
.A1(n_644),
.A2(n_664),
.B1(n_677),
.B2(n_689),
.C(n_690),
.Y(n_709)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_645),
.A2(n_648),
.B(n_656),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_651),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_652),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_654),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_657),
.A2(n_660),
.B(n_662),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_661),
.Y(n_660)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_664),
.Y(n_690)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_668),
.Y(n_711)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_669),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_672),
.B(n_674),
.C(n_710),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_675),
.A2(n_691),
.B(n_709),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_677),
.B(n_688),
.Y(n_676)
);

INVx4_ASAP7_75t_L g703 ( 
.A(n_678),
.Y(n_703)
);

INVx4_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_680),
.Y(n_679)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_685),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_686),
.Y(n_685)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_692),
.Y(n_691)
);

OAI21x1_ASAP7_75t_L g692 ( 
.A1(n_693),
.A2(n_699),
.B(n_708),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_694),
.B(n_695),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_694),
.B(n_695),
.Y(n_708)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_697),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_698),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_700),
.B(n_701),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_702),
.B(n_704),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_705),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_706),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_707),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_711),
.B(n_712),
.Y(n_710)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_717),
.Y(n_716)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_719),
.Y(n_718)
);


endmodule