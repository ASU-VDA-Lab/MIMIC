module fake_netlist_6_4748_n_183 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_183);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_183;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_78;
wire n_84;
wire n_66;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_8),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx5p33_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_6),
.Y(n_49)
);

INVxp67_ASAP7_75t_SL g50 ( 
.A(n_14),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_0),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_2),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_5),
.Y(n_72)
);

AND3x1_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_5),
.C(n_8),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AND2x4_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_52),
.Y(n_79)
);

BUFx6f_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_34),
.B1(n_37),
.B2(n_54),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_70),
.B(n_54),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_58),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_40),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_40),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_35),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_65),
.B(n_50),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_82),
.A2(n_73),
.B1(n_71),
.B2(n_68),
.Y(n_92)
);

AO21x2_ASAP7_75t_L g93 ( 
.A1(n_79),
.A2(n_71),
.B(n_57),
.Y(n_93)
);

BUFx2_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_71),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_72),
.B1(n_49),
.B2(n_51),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

NAND3x1_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_72),
.C(n_56),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_56),
.B(n_57),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_78),
.A2(n_85),
.B(n_83),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_100),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g109 ( 
.A1(n_103),
.A2(n_76),
.B(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_81),
.B1(n_59),
.B2(n_51),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_93),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_97),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g116 ( 
.A(n_110),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_115),
.B(n_108),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_117),
.Y(n_121)
);

OAI21x1_ASAP7_75t_L g122 ( 
.A1(n_113),
.A2(n_109),
.B(n_102),
.Y(n_122)
);

NOR2x1_ASAP7_75t_SL g123 ( 
.A(n_121),
.B(n_111),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_118),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_114),
.Y(n_128)
);

NAND2x1p5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_112),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_114),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_120),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_122),
.Y(n_132)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_122),
.B(n_94),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_131),
.A2(n_112),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g136 ( 
.A1(n_128),
.A2(n_110),
.B1(n_84),
.B2(n_130),
.C(n_59),
.Y(n_136)
);

AOI222xp33_ASAP7_75t_L g137 ( 
.A1(n_130),
.A2(n_116),
.B1(n_101),
.B2(n_89),
.C1(n_65),
.C2(n_75),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_131),
.B(n_88),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_80),
.B1(n_94),
.B2(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_127),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_134),
.A2(n_132),
.B(n_123),
.Y(n_143)
);

AOI221x1_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.C(n_67),
.Y(n_144)
);

O2A1O1Ixp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_58),
.B(n_61),
.C(n_66),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_123),
.B(n_133),
.Y(n_146)
);

NOR2xp67_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_125),
.Y(n_147)
);

NAND4xp25_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_62),
.C(n_63),
.D(n_55),
.Y(n_148)
);

AOI321xp33_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_63),
.A3(n_60),
.B1(n_55),
.B2(n_64),
.C(n_67),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_129),
.B1(n_96),
.B2(n_78),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_60),
.C(n_67),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_9),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_147),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_67),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_9),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_64),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_64),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_125),
.Y(n_159)
);

AOI221x1_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_60),
.B1(n_74),
.B2(n_66),
.C(n_61),
.Y(n_160)
);

AND2x2_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_149),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_153),
.B(n_158),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_126),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_155),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_60),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_163),
.A2(n_74),
.B(n_66),
.C(n_61),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_74),
.A3(n_66),
.B1(n_61),
.B2(n_58),
.C1(n_159),
.C2(n_10),
.Y(n_170)
);

OAI322xp33_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_61),
.A3(n_66),
.B1(n_74),
.B2(n_15),
.C1(n_11),
.C2(n_13),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_161),
.A2(n_74),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_22),
.C2(n_24),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g173 ( 
.A1(n_161),
.A2(n_20),
.A3(n_26),
.B1(n_28),
.B2(n_30),
.C1(n_77),
.C2(n_90),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_109),
.B1(n_77),
.B2(n_145),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_165),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_172),
.A2(n_173),
.B(n_170),
.Y(n_178)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_166),
.B1(n_177),
.B2(n_178),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_178),
.A2(n_166),
.B1(n_171),
.B2(n_174),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_180),
.B1(n_181),
.B2(n_164),
.Y(n_183)
);


endmodule