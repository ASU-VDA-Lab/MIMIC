module fake_netlist_5_159_n_2130 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2130);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2130;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1581;
wire n_1463;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_604;
wire n_314;
wire n_433;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_968;
wire n_912;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_336;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_1138;
wire n_364;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_64),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_89),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_73),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_121),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_125),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_153),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_197),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_69),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_164),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_48),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_200),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_13),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_92),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_44),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_51),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_13),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_182),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_49),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_102),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_39),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_191),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_143),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_183),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_90),
.Y(n_261)
);

BUFx10_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_85),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_6),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_220),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_55),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_60),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_165),
.Y(n_269)
);

BUFx8_ASAP7_75t_SL g270 ( 
.A(n_145),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_208),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_62),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_146),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_187),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_141),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_203),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_128),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_202),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_84),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_150),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_77),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_224),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_22),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_194),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_27),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_86),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_46),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_61),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_94),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_98),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_135),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_148),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_171),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_5),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_30),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_87),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_49),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_2),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_185),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_38),
.Y(n_302)
);

INVxp33_ASAP7_75t_SL g303 ( 
.A(n_178),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_122),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_168),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_174),
.Y(n_307)
);

INVx2_ASAP7_75t_SL g308 ( 
.A(n_79),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_88),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_108),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_151),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_100),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_110),
.Y(n_314)
);

BUFx8_ASAP7_75t_SL g315 ( 
.A(n_207),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_8),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_149),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_15),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_206),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_75),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_37),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_45),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_25),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_28),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_19),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_105),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

BUFx2_ASAP7_75t_L g328 ( 
.A(n_219),
.Y(n_328)
);

BUFx2_ASAP7_75t_SL g329 ( 
.A(n_50),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_160),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_114),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_190),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_212),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_68),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_152),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_126),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_196),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_69),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_184),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_60),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_166),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_36),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_115),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_218),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_18),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_14),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_65),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_64),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_27),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_37),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_119),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_188),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_161),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_91),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_111),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_154),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_116),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_62),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_97),
.Y(n_361)
);

BUFx2_ASAP7_75t_R g362 ( 
.A(n_82),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_106),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_107),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_42),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_221),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_50),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_186),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_2),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_65),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_101),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_142),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_19),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_83),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_71),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_21),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_8),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_140),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_170),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_20),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_129),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_155),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_109),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_12),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_104),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_0),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_130),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_38),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_78),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_204),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_10),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_44),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_40),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_56),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_11),
.Y(n_395)
);

BUFx5_ASAP7_75t_L g396 ( 
.A(n_56),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_43),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_31),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_70),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_29),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_53),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_63),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_138),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_9),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_205),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_80),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_22),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_58),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_113),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_34),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_29),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_17),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_81),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_58),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_179),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_35),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_99),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_93),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_144),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_117),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_198),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_40),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_3),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_177),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_216),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_211),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_59),
.Y(n_427)
);

BUFx5_ASAP7_75t_L g428 ( 
.A(n_193),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_59),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_76),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_54),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_137),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_74),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_68),
.Y(n_434)
);

BUFx8_ASAP7_75t_SL g435 ( 
.A(n_118),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_181),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_167),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_95),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_131),
.Y(n_439)
);

CKINVDCx14_ASAP7_75t_R g440 ( 
.A(n_31),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_127),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_45),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_30),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_139),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_328),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_396),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_396),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_396),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_440),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_396),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_349),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_226),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_323),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_250),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_266),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_228),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_346),
.Y(n_461)
);

INVxp67_ASAP7_75t_SL g462 ( 
.A(n_382),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_322),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_228),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_259),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_382),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_322),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_259),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_322),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_268),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_272),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_430),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_322),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_322),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_367),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_367),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_231),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_367),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_367),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_367),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_286),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_428),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_257),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_257),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_369),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_369),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_400),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_400),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_235),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_288),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_442),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_241),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_264),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_280),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_289),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_316),
.Y(n_498)
);

BUFx2_ASAP7_75t_SL g499 ( 
.A(n_276),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_295),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_428),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_321),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_348),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_276),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_354),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_296),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_298),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_227),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_365),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_384),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_299),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_335),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_388),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_335),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_394),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_339),
.Y(n_517)
);

INVxp67_ASAP7_75t_SL g518 ( 
.A(n_232),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_339),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_305),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_399),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_410),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_422),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_347),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_242),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_429),
.Y(n_528)
);

INVxp33_ASAP7_75t_L g529 ( 
.A(n_270),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_237),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_240),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_251),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_310),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_254),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_256),
.Y(n_535)
);

INVxp33_ASAP7_75t_SL g536 ( 
.A(n_242),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_245),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_245),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_229),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_229),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_425),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_425),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_324),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_265),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_243),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_437),
.Y(n_546)
);

INVx1_ASAP7_75t_SL g547 ( 
.A(n_347),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_269),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_325),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_334),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_428),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_428),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_271),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_347),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_329),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_437),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_338),
.Y(n_558)
);

INVxp67_ASAP7_75t_SL g559 ( 
.A(n_274),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_341),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_428),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_277),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_279),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_343),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_281),
.Y(n_565)
);

CKINVDCx14_ASAP7_75t_R g566 ( 
.A(n_379),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_477),
.B(n_294),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_L g568 ( 
.A(n_449),
.B(n_455),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_508),
.B(n_294),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_463),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_454),
.B(n_233),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_518),
.B(n_308),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_L g573 ( 
.A(n_449),
.B(n_243),
.Y(n_573)
);

OAI21x1_ASAP7_75t_L g574 ( 
.A1(n_454),
.A2(n_293),
.B(n_290),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_463),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_483),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_475),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_475),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_447),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_448),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_451),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_491),
.B(n_358),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_308),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_450),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_499),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_530),
.B(n_313),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_452),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_499),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_453),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_467),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_470),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_451),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_455),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_446),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_446),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_474),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_462),
.B(n_438),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_474),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_476),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_531),
.B(n_313),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_539),
.A2(n_311),
.B(n_304),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_473),
.B(n_262),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_479),
.Y(n_606)
);

AND2x4_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_371),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_483),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_480),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_480),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_481),
.Y(n_612)
);

OA21x2_ASAP7_75t_L g613 ( 
.A1(n_539),
.A2(n_327),
.B(n_326),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_SL g614 ( 
.A1(n_460),
.A2(n_249),
.B1(n_300),
.B2(n_284),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_481),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_540),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_466),
.B(n_262),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_464),
.B(n_249),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_534),
.B(n_535),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_466),
.B(n_262),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_544),
.B(n_371),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_548),
.B(n_244),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_501),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_459),
.B(n_247),
.Y(n_624)
);

CKINVDCx20_ASAP7_75t_R g625 ( 
.A(n_465),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_540),
.Y(n_626)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_469),
.A2(n_300),
.B1(n_302),
.B2(n_284),
.Y(n_627)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_459),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_468),
.B(n_456),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_553),
.B(n_562),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_501),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_541),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_551),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_551),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_541),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_552),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_457),
.A2(n_373),
.B1(n_401),
.B2(n_302),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_468),
.B(n_273),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_547),
.B(n_273),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_542),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_552),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_542),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_SL g643 ( 
.A1(n_504),
.A2(n_401),
.B1(n_373),
.B2(n_247),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_458),
.B(n_273),
.Y(n_644)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_526),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_562),
.B(n_244),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_555),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_563),
.B(n_331),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_546),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_557),
.Y(n_653)
);

CKINVDCx8_ASAP7_75t_R g654 ( 
.A(n_471),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_557),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_494),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_484),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_484),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_485),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_563),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_485),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_575),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_583),
.B(n_566),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_631),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_637),
.A2(n_445),
.B1(n_554),
.B2(n_318),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_631),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_583),
.B(n_565),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_R g669 ( 
.A(n_595),
.B(n_512),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_575),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_629),
.B(n_565),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_631),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_631),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_597),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_622),
.B(n_545),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_575),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_577),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_586),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_596),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_596),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_622),
.B(n_461),
.Y(n_681)
);

INVx3_ASAP7_75t_L g682 ( 
.A(n_631),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_577),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_631),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_629),
.B(n_495),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_589),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_577),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_645),
.B(n_536),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_599),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_599),
.B(n_471),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_596),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_633),
.Y(n_692)
);

NAND2xp33_ASAP7_75t_SL g693 ( 
.A(n_605),
.B(n_415),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_597),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_472),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_605),
.B(n_472),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_654),
.B(n_482),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_624),
.B(n_482),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_598),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_597),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_569),
.B(n_492),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_597),
.Y(n_702)
);

INVx5_ASAP7_75t_L g703 ( 
.A(n_571),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_579),
.Y(n_704)
);

NAND2xp33_ASAP7_75t_L g705 ( 
.A(n_571),
.B(n_233),
.Y(n_705)
);

AND3x4_ASAP7_75t_L g706 ( 
.A(n_643),
.B(n_517),
.C(n_514),
.Y(n_706)
);

INVx5_ASAP7_75t_L g707 ( 
.A(n_571),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_579),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_579),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_606),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_580),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_580),
.Y(n_713)
);

NAND3xp33_ASAP7_75t_L g714 ( 
.A(n_646),
.B(n_556),
.C(n_497),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_580),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_569),
.B(n_492),
.Y(n_716)
);

INVx4_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_606),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_584),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_606),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_623),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_633),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_567),
.B(n_497),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_SL g724 ( 
.A(n_654),
.B(n_362),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_584),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_633),
.Y(n_726)
);

INVx1_ASAP7_75t_SL g727 ( 
.A(n_618),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_623),
.Y(n_728)
);

NAND3xp33_ASAP7_75t_L g729 ( 
.A(n_646),
.B(n_572),
.C(n_506),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_623),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_567),
.B(n_500),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_636),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_584),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_654),
.B(n_500),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_639),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_588),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_588),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_617),
.B(n_506),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_588),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_636),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_636),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_633),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_572),
.B(n_507),
.Y(n_743)
);

BUFx6f_ASAP7_75t_SL g744 ( 
.A(n_619),
.Y(n_744)
);

INVx6_ASAP7_75t_L g745 ( 
.A(n_576),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_590),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_581),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_590),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_617),
.B(n_537),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_576),
.B(n_511),
.Y(n_750)
);

XNOR2xp5_ASAP7_75t_L g751 ( 
.A(n_614),
.B(n_519),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_620),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_590),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_647),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_587),
.B(n_486),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_576),
.B(n_511),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_571),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_587),
.B(n_486),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_633),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_647),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_647),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_656),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_656),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_656),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_628),
.A2(n_267),
.B1(n_351),
.B2(n_350),
.Y(n_765)
);

INVxp33_ASAP7_75t_L g766 ( 
.A(n_637),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_578),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_608),
.Y(n_768)
);

INVx3_ASAP7_75t_L g769 ( 
.A(n_634),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_620),
.B(n_520),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_571),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_608),
.Y(n_772)
);

AOI22x1_ASAP7_75t_L g773 ( 
.A1(n_587),
.A2(n_538),
.B1(n_537),
.B2(n_533),
.Y(n_773)
);

INVxp33_ASAP7_75t_L g774 ( 
.A(n_614),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_625),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_634),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_638),
.B(n_644),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_608),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_578),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_648),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_634),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_578),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_648),
.Y(n_783)
);

BUFx4f_ASAP7_75t_L g784 ( 
.A(n_604),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_578),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_638),
.B(n_520),
.Y(n_786)
);

BUFx10_ASAP7_75t_L g787 ( 
.A(n_593),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_585),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_587),
.B(n_487),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_585),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_648),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_573),
.B(n_543),
.C(n_533),
.Y(n_792)
);

AND3x2_ASAP7_75t_L g793 ( 
.A(n_644),
.B(n_525),
.C(n_342),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_591),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_634),
.Y(n_795)
);

AND3x2_ASAP7_75t_L g796 ( 
.A(n_607),
.B(n_345),
.C(n_336),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_649),
.A2(n_303),
.B1(n_498),
.B2(n_496),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_591),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_582),
.B(n_543),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_648),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_592),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_634),
.Y(n_802)
);

NAND2xp33_ASAP7_75t_SL g803 ( 
.A(n_603),
.B(n_252),
.Y(n_803)
);

OAI22xp33_ASAP7_75t_L g804 ( 
.A1(n_603),
.A2(n_370),
.B1(n_376),
.B2(n_360),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_592),
.Y(n_805)
);

OAI22xp33_ASAP7_75t_L g806 ( 
.A1(n_621),
.A2(n_380),
.B1(n_386),
.B2(n_377),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_643),
.Y(n_807)
);

BUFx3_ASAP7_75t_L g808 ( 
.A(n_619),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_594),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_634),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_594),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_619),
.B(n_549),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_619),
.B(n_549),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_661),
.B(n_550),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_601),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_607),
.B(n_550),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_607),
.B(n_558),
.Y(n_817)
);

INVx5_ASAP7_75t_L g818 ( 
.A(n_571),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_784),
.A2(n_613),
.B1(n_604),
.B2(n_607),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_671),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_671),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_689),
.B(n_558),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_669),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_811),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_685),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_723),
.B(n_560),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_731),
.B(n_560),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_701),
.B(n_661),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_716),
.B(n_564),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_743),
.B(n_661),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_752),
.B(n_564),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_681),
.B(n_627),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_L g833 ( 
.A(n_695),
.B(n_568),
.Y(n_833)
);

BUFx6f_ASAP7_75t_SL g834 ( 
.A(n_787),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_767),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_784),
.A2(n_613),
.B1(n_604),
.B2(n_649),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_752),
.B(n_303),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_811),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_668),
.B(n_814),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_815),
.Y(n_840)
);

OAI21xp33_ASAP7_75t_L g841 ( 
.A1(n_675),
.A2(n_478),
.B(n_502),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_815),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_689),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_710),
.B(n_627),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_808),
.B(n_657),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_750),
.B(n_649),
.Y(n_846)
);

OAI22xp33_ASAP7_75t_L g847 ( 
.A1(n_766),
.A2(n_621),
.B1(n_255),
.B2(n_423),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_729),
.B(n_307),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_792),
.B(n_657),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_779),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_784),
.A2(n_604),
.B1(n_613),
.B2(n_649),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_756),
.B(n_641),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_694),
.B(n_641),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_685),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_808),
.A2(n_375),
.B1(n_390),
.B2(n_353),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_782),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_694),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_685),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_700),
.B(n_641),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_700),
.B(n_641),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_745),
.B(n_641),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_745),
.B(n_641),
.Y(n_862)
);

BUFx5_ASAP7_75t_L g863 ( 
.A(n_674),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_745),
.B(n_650),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_745),
.B(n_702),
.Y(n_865)
);

INVxp67_ASAP7_75t_L g866 ( 
.A(n_681),
.Y(n_866)
);

NOR3xp33_ASAP7_75t_L g867 ( 
.A(n_693),
.B(n_630),
.C(n_357),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_782),
.Y(n_868)
);

INVx8_ASAP7_75t_L g869 ( 
.A(n_744),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_698),
.B(n_246),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_786),
.B(n_246),
.Y(n_871)
);

AOI22xp5_ASAP7_75t_SL g872 ( 
.A1(n_774),
.A2(n_252),
.B1(n_423),
.B2(n_255),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_755),
.B(n_758),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_747),
.B(n_538),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_788),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_675),
.B(n_248),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_790),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_688),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_785),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_790),
.Y(n_880)
);

INVx8_ASAP7_75t_L g881 ( 
.A(n_744),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_794),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_794),
.B(n_602),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_798),
.Y(n_884)
);

AND2x4_ASAP7_75t_SL g885 ( 
.A(n_787),
.B(n_301),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_664),
.A2(n_378),
.B1(n_383),
.B2(n_356),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_798),
.B(n_602),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_801),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_801),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_805),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_747),
.B(n_529),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_805),
.B(n_609),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_749),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_809),
.B(n_609),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_714),
.B(n_248),
.Y(n_895)
);

AO22x2_ASAP7_75t_L g896 ( 
.A1(n_706),
.A2(n_690),
.B1(n_735),
.B2(n_696),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_809),
.B(n_610),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_777),
.A2(n_230),
.B1(n_234),
.B2(n_225),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_755),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_802),
.B(n_610),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_785),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_749),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_678),
.B(n_253),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_758),
.B(n_611),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_738),
.B(n_253),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_678),
.B(n_258),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_789),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_789),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_665),
.B(n_611),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_793),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_777),
.A2(n_337),
.B1(n_332),
.B2(n_330),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_665),
.B(n_615),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_686),
.B(n_258),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_749),
.Y(n_914)
);

CKINVDCx20_ASAP7_75t_R g915 ( 
.A(n_775),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_770),
.B(n_426),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_768),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_773),
.B(n_428),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_787),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_721),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_SL g921 ( 
.A(n_797),
.B(n_432),
.C(n_426),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_777),
.A2(n_333),
.B1(n_319),
.B2(n_314),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_777),
.A2(n_749),
.B1(n_817),
.B2(n_816),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_812),
.B(n_432),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_686),
.B(n_804),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_813),
.B(n_433),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_803),
.A2(n_340),
.B1(n_309),
.B2(n_306),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_667),
.B(n_659),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_806),
.B(n_433),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_803),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_768),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_772),
.Y(n_932)
);

INVx8_ASAP7_75t_L g933 ( 
.A(n_744),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_705),
.A2(n_630),
.B(n_524),
.C(n_523),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_799),
.A2(n_409),
.B1(n_417),
.B2(n_418),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_728),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_667),
.B(n_659),
.Y(n_937)
);

AOI22xp5_ASAP7_75t_L g938 ( 
.A1(n_697),
.A2(n_385),
.B1(n_278),
.B2(n_275),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_773),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_734),
.B(n_441),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_778),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_666),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_765),
.B(n_441),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_728),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_730),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_667),
.B(n_659),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_672),
.B(n_659),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_778),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_724),
.B(n_236),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_727),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_818),
.B(n_238),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_796),
.B(n_503),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_780),
.B(n_391),
.Y(n_953)
);

AOI22xp33_ASAP7_75t_L g954 ( 
.A1(n_666),
.A2(n_613),
.B1(n_574),
.B2(n_374),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_783),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_703),
.B(n_239),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_783),
.B(n_505),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_730),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_666),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_672),
.B(n_600),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_704),
.A2(n_312),
.B1(n_261),
.B2(n_263),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_666),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_708),
.B(n_616),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_663),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_672),
.B(n_600),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_807),
.B(n_393),
.C(n_392),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_732),
.Y(n_967)
);

INVx1_ASAP7_75t_SL g968 ( 
.A(n_751),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_706),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_709),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_791),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_712),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_732),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_807),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_791),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_869),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_880),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_917),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_857),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_931),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_839),
.B(n_679),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_833),
.B(n_703),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_861),
.A2(n_726),
.B(n_717),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_932),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_873),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_823),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_821),
.B(n_679),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_833),
.A2(n_829),
.B1(n_826),
.B2(n_827),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_869),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_821),
.B(n_680),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_828),
.B(n_703),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_915),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_964),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_829),
.B(n_680),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_964),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_969),
.Y(n_996)
);

AND2x2_ASAP7_75t_L g997 ( 
.A(n_866),
.B(n_751),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_843),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_830),
.B(n_691),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_875),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_941),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_948),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_874),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_826),
.B(n_691),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_910),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_873),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_846),
.B(n_703),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_827),
.B(n_800),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_845),
.B(n_673),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_893),
.B(n_703),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_824),
.B(n_800),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_822),
.B(n_509),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_838),
.B(n_673),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_874),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_955),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_971),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_857),
.B(n_707),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_840),
.B(n_673),
.Y(n_1018)
);

AOI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_848),
.A2(n_684),
.B1(n_692),
.B2(n_682),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_847),
.B(n_434),
.C(n_431),
.Y(n_1020)
);

BUFx4f_ASAP7_75t_L g1021 ( 
.A(n_869),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_878),
.B(n_682),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_842),
.B(n_845),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_SL g1024 ( 
.A1(n_968),
.A2(n_443),
.B1(n_397),
.B2(n_402),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_877),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_820),
.B(n_682),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_874),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_975),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_878),
.B(n_684),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_857),
.B(n_707),
.Y(n_1030)
);

AOI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_921),
.A2(n_719),
.B1(n_736),
.B2(n_725),
.Y(n_1031)
);

INVxp67_ASAP7_75t_L g1032 ( 
.A(n_891),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_893),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_848),
.A2(n_692),
.B1(n_722),
.B2(n_684),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_881),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_919),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_847),
.B(n_443),
.C(n_404),
.Y(n_1037)
);

AOI22xp33_ASAP7_75t_L g1038 ( 
.A1(n_921),
.A2(n_753),
.B1(n_739),
.B2(n_737),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_952),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_882),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_884),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_888),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_862),
.A2(n_726),
.B(n_717),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_889),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_899),
.A2(n_692),
.B1(n_810),
.B2(n_795),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_907),
.B(n_722),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_908),
.B(n_841),
.Y(n_1047)
);

OAI22xp5_ASAP7_75t_L g1048 ( 
.A1(n_819),
.A2(n_769),
.B1(n_810),
.B2(n_795),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_890),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_864),
.A2(n_726),
.B(n_717),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_957),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_957),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_819),
.A2(n_742),
.B1(n_810),
.B2(n_795),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_904),
.B(n_722),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_939),
.B(n_742),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_893),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_930),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_970),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_854),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_876),
.B(n_510),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_858),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_972),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_883),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_887),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_881),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_893),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_892),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_953),
.B(n_769),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_835),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_905),
.B(n_916),
.Y(n_1070)
);

INVx2_ASAP7_75t_SL g1071 ( 
.A(n_952),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_852),
.A2(n_781),
.B(n_759),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_825),
.B(n_776),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_849),
.B(n_776),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_834),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_836),
.A2(n_574),
.B(n_719),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_737),
.B1(n_739),
.B2(n_736),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_920),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_836),
.B(n_851),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_905),
.B(n_513),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_902),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_881),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_950),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_974),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_851),
.B(n_776),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_894),
.Y(n_1086)
);

AND2x6_ASAP7_75t_SL g1087 ( 
.A(n_844),
.B(n_515),
.Y(n_1087)
);

AND3x1_ASAP7_75t_L g1088 ( 
.A(n_867),
.B(n_521),
.C(n_516),
.Y(n_1088)
);

AND2x6_ASAP7_75t_L g1089 ( 
.A(n_902),
.B(n_725),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_954),
.A2(n_753),
.B1(n_574),
.B2(n_233),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_954),
.A2(n_233),
.B1(n_374),
.B2(n_260),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_930),
.B(n_713),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_924),
.B(n_715),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_897),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_936),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_850),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_856),
.Y(n_1097)
);

CKINVDCx20_ASAP7_75t_R g1098 ( 
.A(n_974),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_914),
.B(n_616),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_868),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_924),
.B(n_733),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_863),
.B(n_923),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_944),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_902),
.Y(n_1104)
);

INVx8_ASAP7_75t_L g1105 ( 
.A(n_933),
.Y(n_1105)
);

AND2x6_ASAP7_75t_SL g1106 ( 
.A(n_844),
.B(n_522),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_885),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_902),
.B(n_757),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_832),
.B(n_527),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_959),
.B(n_746),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_831),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_933),
.Y(n_1112)
);

INVxp67_ASAP7_75t_SL g1113 ( 
.A(n_853),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_925),
.B(n_748),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_933),
.Y(n_1115)
);

AND3x1_ASAP7_75t_SL g1116 ( 
.A(n_872),
.B(n_528),
.C(n_494),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_879),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_901),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_945),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_926),
.A2(n_421),
.B1(n_439),
.B2(n_436),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_916),
.Y(n_1121)
);

INVx2_ASAP7_75t_SL g1122 ( 
.A(n_837),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_940),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_958),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_942),
.B(n_626),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_962),
.B(n_903),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_926),
.B(n_763),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_870),
.B(n_763),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_962),
.B(n_759),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_895),
.B(n_759),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_967),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_844),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_834),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_973),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_963),
.B(n_764),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_867),
.B(n_764),
.Y(n_1136)
);

BUFx4f_ASAP7_75t_L g1137 ( 
.A(n_966),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_896),
.A2(n_374),
.B1(n_372),
.B2(n_260),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_898),
.B(n_626),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_859),
.Y(n_1140)
);

AND2x4_ASAP7_75t_L g1141 ( 
.A(n_911),
.B(n_632),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_860),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_909),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_912),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_928),
.Y(n_1145)
);

AO22x1_ASAP7_75t_L g1146 ( 
.A1(n_895),
.A2(n_416),
.B1(n_395),
.B2(n_407),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_922),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_SL g1148 ( 
.A(n_865),
.B(n_757),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_896),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_937),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_983),
.A2(n_965),
.B(n_960),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_993),
.Y(n_1152)
);

NOR3xp33_ASAP7_75t_SL g1153 ( 
.A(n_992),
.B(n_949),
.C(n_913),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1079),
.A2(n_1076),
.B(n_1113),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1085),
.A2(n_1102),
.B(n_1072),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1102),
.A2(n_781),
.B(n_900),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_988),
.B(n_1070),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_985),
.B(n_871),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_1121),
.B(n_906),
.Y(n_1159)
);

NAND3xp33_ASAP7_75t_L g1160 ( 
.A(n_1120),
.B(n_935),
.C(n_929),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_993),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_1112),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_1109),
.A2(n_943),
.B(n_886),
.C(n_855),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_978),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_998),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_986),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_980),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_995),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_984),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_986),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1084),
.B(n_938),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_SL g1172 ( 
.A(n_1058),
.B(n_927),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1063),
.B(n_896),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1064),
.B(n_961),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_R g1175 ( 
.A(n_992),
.B(n_1036),
.Y(n_1175)
);

CKINVDCx8_ASAP7_75t_R g1176 ( 
.A(n_1112),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_995),
.Y(n_1177)
);

BUFx10_ASAP7_75t_L g1178 ( 
.A(n_1112),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_999),
.A2(n_947),
.B(n_946),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_981),
.A2(n_771),
.B(n_757),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_1024),
.B(n_412),
.C(n_411),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_985),
.B(n_632),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1114),
.A2(n_1091),
.B(n_1130),
.C(n_1067),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1001),
.Y(n_1184)
);

AOI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1149),
.A2(n_419),
.B1(n_424),
.B2(n_368),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1007),
.A2(n_771),
.B(n_757),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1007),
.A2(n_818),
.B(n_771),
.Y(n_1187)
);

AND2x6_ASAP7_75t_L g1188 ( 
.A(n_1056),
.B(n_260),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1086),
.B(n_740),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1006),
.B(n_635),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1004),
.A2(n_934),
.B(n_956),
.C(n_951),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_996),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1112),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1012),
.B(n_487),
.Y(n_1194)
);

AOI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1114),
.A2(n_287),
.B1(n_285),
.B2(n_283),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1094),
.B(n_740),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1078),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1091),
.A2(n_1138),
.B1(n_1090),
.B2(n_990),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_SL g1199 ( 
.A1(n_982),
.A2(n_490),
.B(n_488),
.C(n_493),
.Y(n_1199)
);

AND2x6_ASAP7_75t_L g1200 ( 
.A(n_1056),
.B(n_260),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1002),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_1083),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1095),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1056),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_SL g1205 ( 
.A(n_1058),
.B(n_771),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1080),
.B(n_741),
.Y(n_1206)
);

OAI22xp5_ASAP7_75t_SL g1207 ( 
.A1(n_1098),
.A2(n_414),
.B1(n_282),
.B2(n_292),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1138),
.A2(n_934),
.B1(n_655),
.B2(n_653),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1068),
.A2(n_818),
.B(n_705),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1009),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1143),
.B(n_741),
.Y(n_1211)
);

BUFx12f_ASAP7_75t_L g1212 ( 
.A(n_1075),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1130),
.A2(n_818),
.B(n_760),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_SL g1214 ( 
.A(n_1062),
.B(n_291),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1098),
.A2(n_387),
.B1(n_381),
.B2(n_444),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1056),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1043),
.A2(n_1050),
.B(n_987),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_1057),
.B(n_315),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_994),
.B(n_754),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_976),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1055),
.A2(n_762),
.B(n_761),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1008),
.B(n_762),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1003),
.Y(n_1223)
);

AOI21x1_ASAP7_75t_L g1224 ( 
.A1(n_991),
.A2(n_720),
.B(n_718),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1144),
.B(n_761),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1090),
.A2(n_640),
.B1(n_653),
.B2(n_652),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1147),
.A2(n_260),
.B1(n_374),
.B2(n_372),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1032),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1139),
.A2(n_635),
.B(n_640),
.C(n_642),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1081),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1009),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1062),
.B(n_1006),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1048),
.A2(n_720),
.B(n_718),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1054),
.A2(n_711),
.B(n_699),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1081),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1137),
.B(n_297),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1014),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1095),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1081),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1009),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1137),
.B(n_317),
.Y(n_1241)
);

NOR2xp33_ASAP7_75t_L g1242 ( 
.A(n_997),
.B(n_1122),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1147),
.A2(n_374),
.B1(n_372),
.B2(n_301),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1081),
.Y(n_1244)
);

OAI22xp5_ASAP7_75t_L g1245 ( 
.A1(n_1126),
.A2(n_652),
.B1(n_655),
.B2(n_651),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_R g1246 ( 
.A(n_996),
.B(n_320),
.Y(n_1246)
);

AOI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1139),
.A2(n_352),
.B1(n_361),
.B2(n_363),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1111),
.B(n_435),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_SL g1249 ( 
.A1(n_1108),
.A2(n_687),
.B(n_683),
.C(n_677),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1103),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1023),
.B(n_344),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1053),
.A2(n_676),
.B(n_670),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1092),
.B(n_651),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1139),
.A2(n_420),
.B1(n_355),
.B2(n_359),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_SL g1255 ( 
.A1(n_1092),
.A2(n_670),
.B(n_663),
.C(n_662),
.Y(n_1255)
);

CKINVDCx16_ASAP7_75t_R g1256 ( 
.A(n_976),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1105),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1103),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1022),
.B(n_658),
.Y(n_1259)
);

AND2x4_ASAP7_75t_L g1260 ( 
.A(n_989),
.B(n_489),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1015),
.Y(n_1261)
);

BUFx6f_ASAP7_75t_L g1262 ( 
.A(n_1105),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1029),
.A2(n_493),
.B(n_490),
.C(n_489),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1022),
.B(n_658),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1027),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1127),
.A2(n_372),
.B1(n_660),
.B2(n_658),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1000),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1123),
.B(n_364),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1060),
.B(n_301),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1136),
.A2(n_662),
.B(n_660),
.C(n_5),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1047),
.B(n_660),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1125),
.Y(n_1272)
);

A2O1A1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_1141),
.A2(n_1101),
.B(n_1093),
.C(n_1051),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1141),
.B(n_366),
.Y(n_1274)
);

AOI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1141),
.A2(n_413),
.B1(n_403),
.B2(n_405),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1104),
.Y(n_1276)
);

INVx1_ASAP7_75t_SL g1277 ( 
.A(n_1099),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1133),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1133),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1148),
.A2(n_406),
.B(n_389),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1140),
.B(n_662),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1016),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_1052),
.A2(n_1059),
.B(n_1061),
.C(n_1028),
.Y(n_1283)
);

AO22x1_ASAP7_75t_L g1284 ( 
.A1(n_1132),
.A2(n_571),
.B1(n_4),
.B2(n_6),
.Y(n_1284)
);

AND2x2_ASAP7_75t_SL g1285 ( 
.A(n_1021),
.B(n_1),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1035),
.B(n_96),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1142),
.A2(n_612),
.B(n_600),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1099),
.B(n_1039),
.Y(n_1288)
);

AO21x2_ASAP7_75t_L g1289 ( 
.A1(n_1155),
.A2(n_1034),
.B(n_1019),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1164),
.Y(n_1290)
);

OAI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1154),
.A2(n_1038),
.B(n_1031),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1217),
.A2(n_1135),
.B(n_1142),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1221),
.A2(n_1252),
.B(n_1233),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1202),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1165),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1269),
.B(n_1242),
.Y(n_1296)
);

NOR2xp67_ASAP7_75t_L g1297 ( 
.A(n_1210),
.B(n_1033),
.Y(n_1297)
);

AO21x2_ASAP7_75t_L g1298 ( 
.A1(n_1183),
.A2(n_1074),
.B(n_1110),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1156),
.A2(n_1128),
.B(n_1011),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1210),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1159),
.B(n_1021),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1160),
.B(n_1037),
.C(n_1020),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1167),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1157),
.A2(n_1116),
.B1(n_1088),
.B2(n_1099),
.Y(n_1304)
);

AO31x2_ASAP7_75t_L g1305 ( 
.A1(n_1266),
.A2(n_1110),
.A3(n_1129),
.B(n_1044),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1176),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1169),
.Y(n_1307)
);

NOR2xp67_ASAP7_75t_L g1308 ( 
.A(n_1231),
.B(n_1033),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_SL g1309 ( 
.A1(n_1173),
.A2(n_1031),
.B(n_1038),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1273),
.A2(n_1108),
.B(n_1018),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1198),
.A2(n_1129),
.B1(n_1033),
.B2(n_1066),
.Y(n_1311)
);

BUFx10_ASAP7_75t_L g1312 ( 
.A(n_1166),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1194),
.B(n_1146),
.Y(n_1313)
);

A2O1A1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1163),
.A2(n_1049),
.B(n_1041),
.C(n_1040),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1224),
.A2(n_1145),
.B(n_1077),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1184),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1220),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1151),
.A2(n_1145),
.B(n_1077),
.Y(n_1318)
);

AO32x2_ASAP7_75t_L g1319 ( 
.A1(n_1198),
.A2(n_1066),
.A3(n_1116),
.B1(n_1071),
.B2(n_1107),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1231),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1192),
.Y(n_1321)
);

NOR3xp33_ASAP7_75t_L g1322 ( 
.A(n_1274),
.B(n_1066),
.C(n_1026),
.Y(n_1322)
);

OR2x2_ASAP7_75t_L g1323 ( 
.A(n_1272),
.B(n_1025),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1179),
.A2(n_1013),
.B(n_1046),
.Y(n_1324)
);

AND2x6_ASAP7_75t_L g1325 ( 
.A(n_1204),
.B(n_1035),
.Y(n_1325)
);

OAI22x1_ASAP7_75t_L g1326 ( 
.A1(n_1185),
.A2(n_1106),
.B1(n_1087),
.B2(n_1042),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1266),
.A2(n_1025),
.A3(n_1044),
.B(n_1042),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1227),
.A2(n_1045),
.B(n_979),
.Y(n_1329)
);

AOI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1259),
.A2(n_1118),
.B(n_1100),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1264),
.A2(n_1097),
.B(n_1096),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1272),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1191),
.A2(n_979),
.B(n_1030),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1234),
.A2(n_1117),
.B(n_1134),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1257),
.B(n_1065),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1206),
.A2(n_1219),
.B(n_1222),
.Y(n_1336)
);

AOI221x1_ASAP7_75t_L g1337 ( 
.A1(n_1160),
.A2(n_1119),
.B1(n_1124),
.B2(n_977),
.C(n_1069),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1255),
.A2(n_1017),
.B(n_1073),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1201),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_SL g1340 ( 
.A(n_1204),
.B(n_1150),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1277),
.B(n_1150),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1174),
.A2(n_1010),
.B(n_1115),
.Y(n_1342)
);

NOR2x1_ASAP7_75t_SL g1343 ( 
.A(n_1204),
.B(n_1065),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1253),
.B(n_1073),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1257),
.B(n_1082),
.Y(n_1345)
);

AO21x1_ASAP7_75t_L g1346 ( 
.A1(n_1270),
.A2(n_1172),
.B(n_1208),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_1175),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1213),
.A2(n_1073),
.B(n_1089),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1208),
.A2(n_1089),
.A3(n_1131),
.B(n_1010),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1281),
.A2(n_1105),
.B(n_1115),
.Y(n_1350)
);

OR2x6_ASAP7_75t_L g1351 ( 
.A(n_1262),
.B(n_1286),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1209),
.A2(n_1082),
.B(n_1089),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1228),
.B(n_1005),
.Y(n_1353)
);

INVxp67_ASAP7_75t_L g1354 ( 
.A(n_1223),
.Y(n_1354)
);

CKINVDCx6p67_ASAP7_75t_R g1355 ( 
.A(n_1212),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_L g1356 ( 
.A(n_1262),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1261),
.B(n_1089),
.Y(n_1357)
);

AOI221x1_ASAP7_75t_L g1358 ( 
.A1(n_1207),
.A2(n_570),
.B1(n_612),
.B2(n_9),
.C(n_10),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1271),
.A2(n_570),
.B(n_612),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1229),
.A2(n_571),
.A3(n_7),
.B(n_11),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1171),
.B(n_1),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1282),
.B(n_7),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1287),
.A2(n_159),
.B(n_223),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1247),
.A2(n_612),
.B1(n_14),
.B2(n_16),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1162),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1288),
.B(n_12),
.Y(n_1366)
);

INVx5_ASAP7_75t_L g1367 ( 
.A(n_1216),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1182),
.B(n_17),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1182),
.B(n_18),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1170),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1199),
.A2(n_217),
.B(n_215),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1162),
.Y(n_1372)
);

OAI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1243),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1211),
.A2(n_214),
.B(n_213),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1158),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1375)
);

AOI21x1_ASAP7_75t_L g1376 ( 
.A1(n_1251),
.A2(n_209),
.B(n_195),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1267),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1226),
.A2(n_26),
.A3(n_28),
.B(n_32),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1268),
.B(n_1218),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1190),
.B(n_26),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1211),
.A2(n_1189),
.B(n_1196),
.Y(n_1381)
);

O2A1O1Ixp5_ASAP7_75t_SL g1382 ( 
.A1(n_1236),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1190),
.B(n_33),
.Y(n_1383)
);

AO21x1_ASAP7_75t_L g1384 ( 
.A1(n_1226),
.A2(n_36),
.B(n_39),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1278),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1158),
.B(n_41),
.Y(n_1386)
);

BUFx10_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1225),
.A2(n_112),
.B(n_189),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1180),
.A2(n_1186),
.B(n_1187),
.Y(n_1389)
);

AO221x2_ASAP7_75t_L g1390 ( 
.A1(n_1284),
.A2(n_41),
.B1(n_43),
.B2(n_46),
.C(n_47),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1283),
.B(n_47),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1247),
.B(n_48),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1254),
.B(n_1275),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_SL g1394 ( 
.A1(n_1185),
.A2(n_123),
.B(n_180),
.Y(n_1394)
);

O2A1O1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1241),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1240),
.B(n_192),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1254),
.B(n_52),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1249),
.A2(n_124),
.B(n_157),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1205),
.A2(n_120),
.B(n_156),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1214),
.A2(n_103),
.B(n_147),
.Y(n_1400)
);

NAND2xp33_ASAP7_75t_SL g1401 ( 
.A(n_1153),
.B(n_57),
.Y(n_1401)
);

CKINVDCx6p67_ASAP7_75t_R g1402 ( 
.A(n_1279),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1265),
.B(n_57),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1275),
.B(n_63),
.Y(n_1404)
);

AOI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1280),
.A2(n_169),
.B(n_133),
.Y(n_1405)
);

O2A1O1Ixp33_ASAP7_75t_SL g1406 ( 
.A1(n_1232),
.A2(n_134),
.B(n_136),
.C(n_70),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1195),
.A2(n_66),
.B(n_67),
.C(n_1181),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1240),
.A2(n_66),
.B(n_67),
.Y(n_1408)
);

AO31x2_ASAP7_75t_L g1409 ( 
.A1(n_1245),
.A2(n_1152),
.A3(n_1161),
.B(n_1177),
.Y(n_1409)
);

AOI211x1_ASAP7_75t_L g1410 ( 
.A1(n_1245),
.A2(n_1285),
.B(n_1207),
.C(n_1215),
.Y(n_1410)
);

OAI21xp5_ASAP7_75t_L g1411 ( 
.A1(n_1263),
.A2(n_1258),
.B(n_1250),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1197),
.A2(n_1238),
.B(n_1203),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1168),
.A2(n_1276),
.B(n_1195),
.Y(n_1413)
);

INVx1_ASAP7_75t_SL g1414 ( 
.A(n_1237),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1286),
.B(n_1260),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_SL g1416 ( 
.A(n_1216),
.B(n_1230),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1260),
.B(n_1230),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1246),
.Y(n_1418)
);

BUFx8_ASAP7_75t_L g1419 ( 
.A(n_1162),
.Y(n_1419)
);

AOI21xp33_ASAP7_75t_L g1420 ( 
.A1(n_1215),
.A2(n_1235),
.B(n_1244),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1239),
.B(n_1193),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1239),
.B(n_1193),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1256),
.A2(n_1188),
.B1(n_1200),
.B2(n_1193),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1188),
.Y(n_1424)
);

BUFx2_ASAP7_75t_L g1425 ( 
.A(n_1188),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1178),
.B(n_988),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1221),
.A2(n_1252),
.B(n_1233),
.Y(n_1427)
);

OA21x2_ASAP7_75t_L g1428 ( 
.A1(n_1155),
.A2(n_1154),
.B(n_1221),
.Y(n_1428)
);

NOR4xp25_ASAP7_75t_L g1429 ( 
.A(n_1270),
.B(n_1070),
.C(n_1138),
.D(n_1183),
.Y(n_1429)
);

AND2x4_ASAP7_75t_L g1430 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1157),
.B(n_988),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1217),
.A2(n_1154),
.B(n_1079),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1269),
.B(n_997),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1221),
.A2(n_1252),
.B(n_1233),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1163),
.A2(n_988),
.B(n_1070),
.C(n_829),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1164),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1257),
.B(n_1262),
.Y(n_1437)
);

O2A1O1Ixp5_ASAP7_75t_L g1438 ( 
.A1(n_1183),
.A2(n_829),
.B(n_1070),
.C(n_870),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1290),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1440)
);

AND2x6_ASAP7_75t_L g1441 ( 
.A(n_1423),
.B(n_1424),
.Y(n_1441)
);

AOI221x1_ASAP7_75t_L g1442 ( 
.A1(n_1435),
.A2(n_1364),
.B1(n_1393),
.B2(n_1302),
.C(n_1407),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1370),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1432),
.A2(n_1337),
.B(n_1291),
.Y(n_1444)
);

AO21x2_ASAP7_75t_L g1445 ( 
.A1(n_1291),
.A2(n_1346),
.B(n_1292),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1303),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1385),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_L g1448 ( 
.A1(n_1392),
.A2(n_1404),
.B(n_1397),
.C(n_1361),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1433),
.B(n_1296),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1390),
.A2(n_1302),
.B1(n_1431),
.B2(n_1384),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1390),
.A2(n_1373),
.B1(n_1375),
.B2(n_1379),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1438),
.A2(n_1310),
.B(n_1336),
.Y(n_1452)
);

NAND2xp33_ASAP7_75t_L g1453 ( 
.A(n_1325),
.B(n_1322),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1332),
.Y(n_1454)
);

AO21x2_ASAP7_75t_L g1455 ( 
.A1(n_1429),
.A2(n_1333),
.B(n_1324),
.Y(n_1455)
);

BUFx2_ASAP7_75t_R g1456 ( 
.A(n_1418),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1409),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1409),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1318),
.A2(n_1324),
.B(n_1299),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1307),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1334),
.Y(n_1461)
);

AO21x2_ASAP7_75t_L g1462 ( 
.A1(n_1429),
.A2(n_1309),
.B(n_1330),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1315),
.A2(n_1371),
.B(n_1331),
.Y(n_1463)
);

BUFx2_ASAP7_75t_L g1464 ( 
.A(n_1354),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1304),
.B(n_1323),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1321),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1415),
.B(n_1304),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1426),
.B(n_1313),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1316),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1339),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1341),
.B(n_1295),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1359),
.A2(n_1381),
.B(n_1358),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1366),
.B(n_1368),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1344),
.B(n_1414),
.Y(n_1474)
);

OAI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1314),
.A2(n_1329),
.B(n_1413),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1391),
.A2(n_1373),
.B(n_1357),
.C(n_1395),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1311),
.Y(n_1477)
);

OA21x2_ASAP7_75t_L g1478 ( 
.A1(n_1411),
.A2(n_1374),
.B(n_1363),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1298),
.A2(n_1289),
.B(n_1311),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1401),
.A2(n_1326),
.B1(n_1408),
.B2(n_1386),
.Y(n_1480)
);

OR2x6_ASAP7_75t_L g1481 ( 
.A(n_1350),
.B(n_1410),
.Y(n_1481)
);

OAI21x1_ASAP7_75t_L g1482 ( 
.A1(n_1405),
.A2(n_1428),
.B(n_1348),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1347),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1428),
.A2(n_1348),
.B(n_1334),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1414),
.B(n_1377),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1349),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1436),
.Y(n_1487)
);

AOI22xp33_ASAP7_75t_SL g1488 ( 
.A1(n_1410),
.A2(n_1403),
.B1(n_1394),
.B2(n_1362),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1319),
.A2(n_1412),
.A3(n_1327),
.B(n_1340),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1376),
.A2(n_1411),
.B(n_1388),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1399),
.A2(n_1400),
.B(n_1382),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1329),
.A2(n_1301),
.B(n_1380),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1317),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_L g1494 ( 
.A(n_1325),
.B(n_1423),
.Y(n_1494)
);

OAI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1417),
.A2(n_1345),
.B1(n_1383),
.B2(n_1369),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1349),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1300),
.B(n_1320),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1297),
.B(n_1308),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1421),
.A2(n_1422),
.B(n_1297),
.Y(n_1499)
);

INVx3_ASAP7_75t_SL g1500 ( 
.A(n_1306),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1387),
.A2(n_1420),
.B1(n_1312),
.B2(n_1306),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1353),
.A2(n_1387),
.B1(n_1294),
.B2(n_1306),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1378),
.Y(n_1503)
);

OAI21x1_ASAP7_75t_L g1504 ( 
.A1(n_1398),
.A2(n_1327),
.B(n_1349),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1327),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1378),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1378),
.Y(n_1507)
);

OAI21x1_ASAP7_75t_L g1508 ( 
.A1(n_1338),
.A2(n_1319),
.B(n_1305),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1355),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1338),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1367),
.Y(n_1511)
);

NAND2x1p5_ASAP7_75t_L g1512 ( 
.A(n_1367),
.B(n_1437),
.Y(n_1512)
);

INVx2_ASAP7_75t_L g1513 ( 
.A(n_1305),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1305),
.A2(n_1319),
.B(n_1425),
.Y(n_1514)
);

INVx6_ASAP7_75t_L g1515 ( 
.A(n_1419),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1416),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1335),
.B(n_1437),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1360),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1360),
.Y(n_1519)
);

OAI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1328),
.A2(n_1430),
.B1(n_1367),
.B2(n_1356),
.Y(n_1520)
);

OAI21x1_ASAP7_75t_L g1521 ( 
.A1(n_1406),
.A2(n_1343),
.B(n_1325),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1365),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1402),
.A2(n_1325),
.B1(n_1419),
.B2(n_1328),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1365),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1356),
.A2(n_988),
.B1(n_1393),
.B2(n_1358),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1372),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1430),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1372),
.A2(n_1427),
.B(n_1293),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1431),
.B(n_1157),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1431),
.B(n_1157),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1431),
.B(n_1157),
.Y(n_1531)
);

OA21x2_ASAP7_75t_L g1532 ( 
.A1(n_1432),
.A2(n_1337),
.B(n_1291),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_SL g1533 ( 
.A(n_1370),
.B(n_1166),
.Y(n_1533)
);

NOR2x1_ASAP7_75t_R g1534 ( 
.A(n_1370),
.B(n_1166),
.Y(n_1534)
);

OAI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1535)
);

OAI21x1_ASAP7_75t_SL g1536 ( 
.A1(n_1394),
.A2(n_1384),
.B(n_1346),
.Y(n_1536)
);

BUFx8_ASAP7_75t_L g1537 ( 
.A(n_1306),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1290),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_SL g1539 ( 
.A1(n_1435),
.A2(n_1183),
.B(n_1198),
.C(n_1393),
.Y(n_1539)
);

BUFx2_ASAP7_75t_L g1540 ( 
.A(n_1332),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1409),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1390),
.A2(n_1070),
.B1(n_988),
.B2(n_1393),
.Y(n_1543)
);

OR2x6_ASAP7_75t_L g1544 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1390),
.A2(n_1070),
.B1(n_988),
.B2(n_1393),
.Y(n_1545)
);

NAND2x1p5_ASAP7_75t_L g1546 ( 
.A(n_1367),
.B(n_1033),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1390),
.A2(n_1070),
.B1(n_988),
.B2(n_1393),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1549)
);

AO21x2_ASAP7_75t_L g1550 ( 
.A1(n_1432),
.A2(n_1291),
.B(n_1389),
.Y(n_1550)
);

NAND2x1p5_ASAP7_75t_L g1551 ( 
.A(n_1367),
.B(n_1033),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1552)
);

NOR2xp67_ASAP7_75t_L g1553 ( 
.A(n_1370),
.B(n_1083),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1431),
.B(n_1157),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1393),
.A2(n_988),
.B1(n_1358),
.B2(n_1198),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1396),
.B(n_1351),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_L g1557 ( 
.A1(n_1390),
.A2(n_1070),
.B1(n_988),
.B2(n_1393),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1393),
.A2(n_988),
.B1(n_829),
.B2(n_1070),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1290),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_1321),
.Y(n_1561)
);

OAI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1431),
.B(n_988),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1290),
.Y(n_1565)
);

AOI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1330),
.A2(n_1331),
.B(n_1352),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1409),
.Y(n_1567)
);

OAI21x1_ASAP7_75t_L g1568 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1379),
.A2(n_988),
.B1(n_829),
.B2(n_1393),
.Y(n_1569)
);

AO21x2_ASAP7_75t_L g1570 ( 
.A1(n_1432),
.A2(n_1291),
.B(n_1389),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1370),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1419),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1370),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1433),
.B(n_1296),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1396),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_SL g1576 ( 
.A1(n_1394),
.A2(n_1384),
.B(n_1346),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1432),
.A2(n_1337),
.B(n_1291),
.Y(n_1577)
);

XOR2x2_ASAP7_75t_L g1578 ( 
.A(n_1410),
.B(n_706),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1432),
.A2(n_1337),
.B(n_1291),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1396),
.B(n_1351),
.Y(n_1580)
);

OA21x2_ASAP7_75t_L g1581 ( 
.A1(n_1432),
.A2(n_1337),
.B(n_1291),
.Y(n_1581)
);

AOI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1379),
.A2(n_988),
.B1(n_829),
.B2(n_1393),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1433),
.B(n_1296),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1396),
.B(n_1351),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_SL g1585 ( 
.A1(n_1390),
.A2(n_464),
.B1(n_465),
.B2(n_460),
.Y(n_1585)
);

BUFx3_ASAP7_75t_L g1586 ( 
.A(n_1419),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1419),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1323),
.B(n_1431),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1393),
.A2(n_988),
.B1(n_829),
.B2(n_1070),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_R g1590 ( 
.A(n_1370),
.B(n_1166),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1317),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1396),
.B(n_1351),
.Y(n_1592)
);

OAI211xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1435),
.A2(n_988),
.B(n_878),
.C(n_1121),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_L g1594 ( 
.A1(n_1293),
.A2(n_1434),
.B(n_1427),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1564),
.B(n_1574),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1585),
.A2(n_1582),
.B1(n_1569),
.B2(n_1451),
.Y(n_1597)
);

INVx1_ASAP7_75t_SL g1598 ( 
.A(n_1583),
.Y(n_1598)
);

OA21x2_ASAP7_75t_L g1599 ( 
.A1(n_1504),
.A2(n_1475),
.B(n_1452),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1585),
.A2(n_1451),
.B1(n_1557),
.B2(n_1547),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1588),
.B(n_1467),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1517),
.B(n_1474),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1485),
.B(n_1465),
.Y(n_1604)
);

NAND2x1_ASAP7_75t_L g1605 ( 
.A(n_1440),
.B(n_1542),
.Y(n_1605)
);

A2O1A1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1448),
.A2(n_1589),
.B(n_1559),
.C(n_1557),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_SL g1607 ( 
.A1(n_1546),
.A2(n_1551),
.B(n_1531),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1543),
.A2(n_1547),
.B1(n_1545),
.B2(n_1450),
.Y(n_1608)
);

OA22x2_ASAP7_75t_L g1609 ( 
.A1(n_1481),
.A2(n_1442),
.B1(n_1468),
.B2(n_1492),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_1443),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1468),
.B(n_1454),
.Y(n_1611)
);

INVx2_ASAP7_75t_SL g1612 ( 
.A(n_1537),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1471),
.B(n_1540),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1593),
.A2(n_1555),
.B(n_1525),
.C(n_1545),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1543),
.A2(n_1488),
.B1(n_1530),
.B2(n_1554),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1446),
.B(n_1460),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1488),
.A2(n_1501),
.B1(n_1525),
.B2(n_1480),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1477),
.B(n_1539),
.Y(n_1618)
);

O2A1O1Ixp33_ASAP7_75t_L g1619 ( 
.A1(n_1593),
.A2(n_1539),
.B(n_1476),
.C(n_1576),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1477),
.B(n_1441),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_SL g1621 ( 
.A1(n_1546),
.A2(n_1551),
.B(n_1511),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1441),
.B(n_1469),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1482),
.A2(n_1484),
.B(n_1508),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1441),
.B(n_1470),
.Y(n_1624)
);

O2A1O1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1476),
.A2(n_1536),
.B(n_1480),
.C(n_1495),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1522),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1556),
.B(n_1580),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1505),
.A2(n_1496),
.B(n_1486),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1487),
.B(n_1538),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1584),
.B(n_1592),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1550),
.A2(n_1570),
.B(n_1453),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1501),
.A2(n_1502),
.B1(n_1515),
.B2(n_1565),
.Y(n_1632)
);

AOI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1445),
.A2(n_1453),
.B(n_1581),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_SL g1634 ( 
.A1(n_1511),
.A2(n_1590),
.B(n_1534),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1443),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1494),
.A2(n_1491),
.B(n_1490),
.C(n_1575),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1441),
.B(n_1560),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1445),
.A2(n_1581),
.B(n_1532),
.Y(n_1638)
);

O2A1O1Ixp5_ASAP7_75t_L g1639 ( 
.A1(n_1503),
.A2(n_1506),
.B(n_1507),
.C(n_1518),
.Y(n_1639)
);

O2A1O1Ixp33_ASAP7_75t_L g1640 ( 
.A1(n_1481),
.A2(n_1494),
.B(n_1500),
.C(n_1440),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1441),
.B(n_1462),
.Y(n_1641)
);

NOR2xp67_ASAP7_75t_L g1642 ( 
.A(n_1553),
.B(n_1447),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_SL g1643 ( 
.A(n_1575),
.B(n_1497),
.Y(n_1643)
);

BUFx12f_ASAP7_75t_L g1644 ( 
.A(n_1466),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1527),
.B(n_1526),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1526),
.B(n_1481),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1466),
.B(n_1561),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1464),
.B(n_1462),
.Y(n_1648)
);

OAI22xp5_ASAP7_75t_L g1649 ( 
.A1(n_1515),
.A2(n_1523),
.B1(n_1500),
.B2(n_1586),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1440),
.B(n_1542),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_SL g1651 ( 
.A1(n_1511),
.A2(n_1542),
.B(n_1544),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1447),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1499),
.Y(n_1653)
);

NOR2xp67_ASAP7_75t_L g1654 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1455),
.B(n_1513),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1455),
.B(n_1513),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1537),
.Y(n_1657)
);

O2A1O1Ixp5_ASAP7_75t_L g1658 ( 
.A1(n_1519),
.A2(n_1566),
.B(n_1516),
.C(n_1510),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1444),
.B(n_1532),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1515),
.A2(n_1523),
.B1(n_1572),
.B2(n_1586),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1544),
.B(n_1572),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1444),
.B(n_1532),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1578),
.B(n_1524),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_L g1664 ( 
.A(n_1571),
.B(n_1573),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1444),
.B(n_1581),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1578),
.B(n_1512),
.Y(n_1666)
);

AOI31xp33_ASAP7_75t_L g1667 ( 
.A1(n_1512),
.A2(n_1483),
.A3(n_1520),
.B(n_1591),
.Y(n_1667)
);

INVx3_ASAP7_75t_L g1668 ( 
.A(n_1498),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1537),
.Y(n_1669)
);

INVx6_ASAP7_75t_L g1670 ( 
.A(n_1587),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1493),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1533),
.B(n_1587),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1509),
.A2(n_1472),
.B1(n_1514),
.B2(n_1577),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1509),
.A2(n_1472),
.B1(n_1514),
.B2(n_1577),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1577),
.B(n_1579),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1579),
.A2(n_1472),
.B(n_1483),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1514),
.B(n_1479),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1579),
.B(n_1479),
.Y(n_1678)
);

O2A1O1Ixp5_ASAP7_75t_L g1679 ( 
.A1(n_1510),
.A2(n_1567),
.B(n_1457),
.C(n_1458),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_SL g1680 ( 
.A1(n_1478),
.A2(n_1459),
.B(n_1463),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1489),
.B(n_1521),
.Y(n_1681)
);

OAI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1458),
.A2(n_1541),
.B1(n_1567),
.B2(n_1456),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1489),
.B(n_1491),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1461),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1463),
.A2(n_1563),
.B(n_1535),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1463),
.B(n_1528),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1528),
.B(n_1548),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1594),
.A2(n_1549),
.B(n_1552),
.C(n_1558),
.Y(n_1688)
);

AND2x4_ASAP7_75t_L g1689 ( 
.A(n_1562),
.B(n_1568),
.Y(n_1689)
);

AOI21xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1569),
.A2(n_1183),
.B(n_1435),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1585),
.A2(n_1091),
.B1(n_1582),
.B2(n_1569),
.Y(n_1692)
);

CKINVDCx20_ASAP7_75t_R g1693 ( 
.A(n_1561),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1694)
);

NOR2xp67_ASAP7_75t_L g1695 ( 
.A(n_1553),
.B(n_1370),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1452),
.A2(n_1198),
.B(n_1183),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1449),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1537),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1564),
.B(n_1529),
.Y(n_1699)
);

CKINVDCx5p33_ASAP7_75t_R g1700 ( 
.A(n_1443),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1588),
.B(n_1465),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1585),
.A2(n_1091),
.B1(n_1582),
.B2(n_1569),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1703)
);

O2A1O1Ixp33_ASAP7_75t_L g1704 ( 
.A1(n_1559),
.A2(n_1435),
.B(n_829),
.C(n_1589),
.Y(n_1704)
);

OA21x2_ASAP7_75t_L g1705 ( 
.A1(n_1504),
.A2(n_1475),
.B(n_1452),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1454),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1473),
.B(n_1449),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1559),
.A2(n_1435),
.B(n_829),
.C(n_1589),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1585),
.A2(n_1091),
.B1(n_1582),
.B2(n_1569),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1588),
.B(n_1465),
.Y(n_1710)
);

INVx3_ASAP7_75t_SL g1711 ( 
.A(n_1443),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1588),
.B(n_1465),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1588),
.B(n_1465),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1564),
.B(n_775),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1588),
.B(n_1465),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1439),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_SL g1717 ( 
.A1(n_1569),
.A2(n_1183),
.B(n_1435),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1569),
.A2(n_1183),
.B(n_1435),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1511),
.Y(n_1719)
);

OA22x2_ASAP7_75t_L g1720 ( 
.A1(n_1569),
.A2(n_1582),
.B1(n_1358),
.B2(n_706),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_SL g1721 ( 
.A1(n_1569),
.A2(n_1183),
.B(n_1435),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1439),
.Y(n_1722)
);

INVxp33_ASAP7_75t_L g1723 ( 
.A(n_1449),
.Y(n_1723)
);

CKINVDCx12_ASAP7_75t_R g1724 ( 
.A(n_1534),
.Y(n_1724)
);

O2A1O1Ixp33_ASAP7_75t_L g1725 ( 
.A1(n_1559),
.A2(n_1435),
.B(n_829),
.C(n_1589),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1704),
.A2(n_1725),
.B(n_1708),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1604),
.B(n_1600),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1648),
.B(n_1641),
.Y(n_1728)
);

OR2x2_ASAP7_75t_SL g1729 ( 
.A(n_1622),
.B(n_1624),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1639),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1602),
.B(n_1646),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1606),
.A2(n_1702),
.B(n_1692),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1714),
.B(n_1600),
.Y(n_1733)
);

OAI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1692),
.A2(n_1709),
.B(n_1702),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1641),
.B(n_1655),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1684),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1653),
.Y(n_1737)
);

NOR2x1_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1651),
.Y(n_1738)
);

BUFx6f_ASAP7_75t_L g1739 ( 
.A(n_1605),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1683),
.B(n_1681),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1655),
.B(n_1656),
.Y(n_1741)
);

AOI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1638),
.A2(n_1633),
.B(n_1685),
.Y(n_1742)
);

OR2x6_ASAP7_75t_L g1743 ( 
.A(n_1640),
.B(n_1631),
.Y(n_1743)
);

INVx2_ASAP7_75t_SL g1744 ( 
.A(n_1616),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1691),
.B(n_1694),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1716),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1722),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1620),
.B(n_1673),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1622),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1691),
.B(n_1694),
.Y(n_1750)
);

NAND3xp33_ASAP7_75t_L g1751 ( 
.A(n_1709),
.B(n_1601),
.C(n_1617),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1597),
.A2(n_1601),
.B1(n_1720),
.B2(n_1608),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1679),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1650),
.B(n_1636),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1629),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1689),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1617),
.A2(n_1720),
.B(n_1614),
.Y(n_1757)
);

NAND2x1_ASAP7_75t_L g1758 ( 
.A(n_1650),
.B(n_1607),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1673),
.B(n_1674),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1699),
.B(n_1701),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1656),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1623),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1611),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1689),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1706),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1699),
.B(n_1710),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1690),
.B(n_1717),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1674),
.B(n_1712),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1624),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1661),
.Y(n_1770)
);

AND2x4_ASAP7_75t_L g1771 ( 
.A(n_1668),
.B(n_1687),
.Y(n_1771)
);

INVx3_ASAP7_75t_L g1772 ( 
.A(n_1686),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1658),
.Y(n_1773)
);

AO21x2_ASAP7_75t_L g1774 ( 
.A1(n_1678),
.A2(n_1680),
.B(n_1696),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1613),
.Y(n_1775)
);

OA21x2_ASAP7_75t_L g1776 ( 
.A1(n_1659),
.A2(n_1662),
.B(n_1665),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1626),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1637),
.B(n_1677),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1693),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1659),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1675),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1609),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1609),
.B(n_1596),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1618),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1595),
.B(n_1703),
.Y(n_1785)
);

CKINVDCx5p33_ASAP7_75t_R g1786 ( 
.A(n_1610),
.Y(n_1786)
);

AO21x2_ASAP7_75t_L g1787 ( 
.A1(n_1688),
.A2(n_1721),
.B(n_1718),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1635),
.Y(n_1788)
);

HB1xp67_ASAP7_75t_L g1789 ( 
.A(n_1713),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1608),
.A2(n_1615),
.B1(n_1632),
.B2(n_1667),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1670),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1715),
.B(n_1603),
.Y(n_1792)
);

AO21x2_ASAP7_75t_L g1793 ( 
.A1(n_1682),
.A2(n_1615),
.B(n_1619),
.Y(n_1793)
);

INVxp67_ASAP7_75t_L g1794 ( 
.A(n_1707),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1599),
.Y(n_1795)
);

BUFx2_ASAP7_75t_L g1796 ( 
.A(n_1599),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1652),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1705),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1746),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1734),
.A2(n_1625),
.B1(n_1632),
.B2(n_1697),
.C(n_1598),
.Y(n_1800)
);

INVx3_ASAP7_75t_L g1801 ( 
.A(n_1756),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1746),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1747),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_1762),
.Y(n_1804)
);

OAI221xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1752),
.A2(n_1666),
.B1(n_1634),
.B2(n_1663),
.C(n_1672),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1778),
.B(n_1630),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1735),
.B(n_1649),
.Y(n_1807)
);

AO21x2_ASAP7_75t_L g1808 ( 
.A1(n_1742),
.A2(n_1649),
.B(n_1660),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1740),
.B(n_1723),
.Y(n_1809)
);

INVxp67_ASAP7_75t_R g1810 ( 
.A(n_1759),
.Y(n_1810)
);

AND2x2_ASAP7_75t_L g1811 ( 
.A(n_1748),
.B(n_1627),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1737),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1748),
.B(n_1645),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1759),
.B(n_1660),
.Y(n_1814)
);

AOI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1767),
.A2(n_1732),
.B(n_1726),
.Y(n_1815)
);

NOR2xp33_ASAP7_75t_L g1816 ( 
.A(n_1751),
.B(n_1643),
.Y(n_1816)
);

INVxp67_ASAP7_75t_SL g1817 ( 
.A(n_1730),
.Y(n_1817)
);

INVxp67_ASAP7_75t_L g1818 ( 
.A(n_1728),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1764),
.B(n_1719),
.Y(n_1819)
);

INVxp67_ASAP7_75t_SL g1820 ( 
.A(n_1730),
.Y(n_1820)
);

OR2x6_ASAP7_75t_L g1821 ( 
.A(n_1743),
.B(n_1621),
.Y(n_1821)
);

AOI31xp33_ASAP7_75t_L g1822 ( 
.A1(n_1751),
.A2(n_1669),
.A3(n_1612),
.B(n_1647),
.Y(n_1822)
);

CKINVDCx6p67_ASAP7_75t_R g1823 ( 
.A(n_1743),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1728),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1735),
.B(n_1776),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1739),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1772),
.B(n_1628),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1784),
.B(n_1671),
.Y(n_1828)
);

BUFx2_ASAP7_75t_L g1829 ( 
.A(n_1771),
.Y(n_1829)
);

AND2x2_ASAP7_75t_L g1830 ( 
.A(n_1774),
.B(n_1776),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1771),
.B(n_1698),
.Y(n_1831)
);

AOI33xp33_ASAP7_75t_L g1832 ( 
.A1(n_1800),
.A2(n_1783),
.A3(n_1782),
.B1(n_1773),
.B2(n_1757),
.B3(n_1753),
.Y(n_1832)
);

OR2x2_ASAP7_75t_L g1833 ( 
.A(n_1824),
.B(n_1825),
.Y(n_1833)
);

OAI31xp33_ASAP7_75t_L g1834 ( 
.A1(n_1815),
.A2(n_1790),
.A3(n_1783),
.B(n_1782),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1815),
.A2(n_1757),
.B1(n_1767),
.B2(n_1738),
.Y(n_1835)
);

OAI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1822),
.A2(n_1743),
.B1(n_1758),
.B2(n_1768),
.Y(n_1836)
);

OAI221xp5_ASAP7_75t_L g1837 ( 
.A1(n_1805),
.A2(n_1733),
.B1(n_1758),
.B2(n_1760),
.C(n_1766),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1799),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1799),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1824),
.B(n_1768),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1802),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1826),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1802),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1816),
.A2(n_1793),
.B1(n_1787),
.B2(n_1800),
.Y(n_1844)
);

BUFx2_ASAP7_75t_L g1845 ( 
.A(n_1819),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1816),
.A2(n_1745),
.B1(n_1750),
.B2(n_1775),
.C(n_1794),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1803),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1819),
.Y(n_1848)
);

NOR4xp25_ASAP7_75t_SL g1849 ( 
.A(n_1805),
.B(n_1796),
.C(n_1773),
.D(n_1737),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_1831),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1814),
.A2(n_1793),
.B1(n_1787),
.B2(n_1754),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1829),
.B(n_1810),
.Y(n_1852)
);

AND2x4_ASAP7_75t_SL g1853 ( 
.A(n_1821),
.B(n_1739),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1809),
.B(n_1789),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1801),
.B(n_1754),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_1812),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1819),
.Y(n_1857)
);

NAND4xp25_ASAP7_75t_L g1858 ( 
.A(n_1828),
.B(n_1784),
.C(n_1727),
.D(n_1749),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_R g1859 ( 
.A(n_1823),
.B(n_1788),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1804),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1818),
.Y(n_1861)
);

INVx2_ASAP7_75t_SL g1862 ( 
.A(n_1831),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1810),
.B(n_1771),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_L g1864 ( 
.A1(n_1823),
.A2(n_1743),
.B1(n_1749),
.B2(n_1769),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1813),
.B(n_1769),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1818),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1813),
.B(n_1763),
.Y(n_1867)
);

AOI222xp33_ASAP7_75t_L g1868 ( 
.A1(n_1809),
.A2(n_1765),
.B1(n_1779),
.B2(n_1792),
.C1(n_1785),
.C2(n_1644),
.Y(n_1868)
);

INVx2_ASAP7_75t_SL g1869 ( 
.A(n_1831),
.Y(n_1869)
);

OAI321xp33_ASAP7_75t_L g1870 ( 
.A1(n_1821),
.A2(n_1753),
.A3(n_1742),
.B1(n_1796),
.B2(n_1795),
.C(n_1798),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1809),
.B(n_1731),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1822),
.A2(n_1729),
.B1(n_1736),
.B2(n_1670),
.Y(n_1872)
);

AOI33xp33_ASAP7_75t_L g1873 ( 
.A1(n_1830),
.A2(n_1744),
.A3(n_1761),
.B1(n_1785),
.B2(n_1780),
.B3(n_1781),
.Y(n_1873)
);

BUFx3_ASAP7_75t_L g1874 ( 
.A(n_1831),
.Y(n_1874)
);

NAND4xp25_ASAP7_75t_L g1875 ( 
.A(n_1828),
.B(n_1741),
.C(n_1642),
.D(n_1761),
.Y(n_1875)
);

AOI221xp5_ASAP7_75t_L g1876 ( 
.A1(n_1817),
.A2(n_1777),
.B1(n_1744),
.B2(n_1731),
.C(n_1755),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1817),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1813),
.B(n_1806),
.Y(n_1879)
);

OAI22xp5_ASAP7_75t_L g1880 ( 
.A1(n_1823),
.A2(n_1729),
.B1(n_1670),
.B2(n_1770),
.Y(n_1880)
);

INVxp67_ASAP7_75t_SL g1881 ( 
.A(n_1820),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_SL g1882 ( 
.A(n_1849),
.B(n_1830),
.C(n_1807),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1856),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1856),
.Y(n_1884)
);

OAI21xp5_ASAP7_75t_L g1885 ( 
.A1(n_1835),
.A2(n_1844),
.B(n_1832),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1838),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1852),
.B(n_1830),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_SL g1888 ( 
.A(n_1836),
.B(n_1786),
.C(n_1700),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1870),
.A2(n_1808),
.B(n_1821),
.Y(n_1889)
);

INVx1_ASAP7_75t_SL g1890 ( 
.A(n_1859),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_L g1891 ( 
.A(n_1858),
.B(n_1811),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1855),
.Y(n_1892)
);

INVx5_ASAP7_75t_L g1893 ( 
.A(n_1842),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1852),
.B(n_1825),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1839),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1860),
.Y(n_1896)
);

INVx4_ASAP7_75t_L g1897 ( 
.A(n_1853),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1877),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1841),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1843),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1847),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1873),
.B(n_1820),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1833),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1842),
.Y(n_1904)
);

INVx1_ASAP7_75t_SL g1905 ( 
.A(n_1859),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1840),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1840),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1861),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1845),
.B(n_1808),
.Y(n_1909)
);

INVx1_ASAP7_75t_SL g1910 ( 
.A(n_1842),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1866),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_SL g1912 ( 
.A(n_1873),
.B(n_1739),
.Y(n_1912)
);

NOR3xp33_ASAP7_75t_L g1913 ( 
.A(n_1832),
.B(n_1695),
.C(n_1654),
.Y(n_1913)
);

AND2x4_ASAP7_75t_L g1914 ( 
.A(n_1855),
.B(n_1801),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1881),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1867),
.B(n_1827),
.Y(n_1916)
);

INVx1_ASAP7_75t_SL g1917 ( 
.A(n_1863),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1865),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1896),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1891),
.B(n_1846),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1891),
.B(n_1876),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1892),
.B(n_1917),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1885),
.B(n_1867),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1885),
.B(n_1865),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1886),
.Y(n_1925)
);

INVx4_ASAP7_75t_L g1926 ( 
.A(n_1893),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1893),
.B(n_1853),
.Y(n_1927)
);

HB1xp67_ASAP7_75t_L g1928 ( 
.A(n_1883),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1902),
.B(n_1879),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1883),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1892),
.B(n_1855),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1908),
.B(n_1834),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_SL g1933 ( 
.A(n_1890),
.B(n_1872),
.Y(n_1933)
);

INVx2_ASAP7_75t_SL g1934 ( 
.A(n_1893),
.Y(n_1934)
);

INVxp67_ASAP7_75t_SL g1935 ( 
.A(n_1906),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1917),
.B(n_1862),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1902),
.B(n_1854),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1908),
.B(n_1806),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1886),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1895),
.Y(n_1940)
);

NOR3xp33_ASAP7_75t_L g1941 ( 
.A(n_1882),
.B(n_1837),
.C(n_1875),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1897),
.B(n_1862),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1907),
.B(n_1871),
.Y(n_1943)
);

NOR2xp33_ASAP7_75t_L g1944 ( 
.A(n_1890),
.B(n_1905),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1896),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1905),
.B(n_1711),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1895),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1897),
.B(n_1869),
.Y(n_1948)
);

NAND2xp33_ASAP7_75t_R g1949 ( 
.A(n_1888),
.B(n_1850),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1897),
.B(n_1869),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1897),
.B(n_1848),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1899),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1897),
.B(n_1857),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1907),
.B(n_1807),
.Y(n_1954)
);

OR2x2_ASAP7_75t_L g1955 ( 
.A(n_1907),
.B(n_1807),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1899),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1900),
.Y(n_1957)
);

AND2x4_ASAP7_75t_L g1958 ( 
.A(n_1893),
.B(n_1874),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1900),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1901),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1914),
.B(n_1906),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1914),
.B(n_1863),
.Y(n_1962)
);

HB1xp67_ASAP7_75t_L g1963 ( 
.A(n_1884),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1901),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1893),
.B(n_1878),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1923),
.B(n_1911),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1944),
.B(n_1916),
.Y(n_1967)
);

OR2x6_ASAP7_75t_L g1968 ( 
.A(n_1926),
.B(n_1934),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1920),
.B(n_1916),
.Y(n_1969)
);

NAND2x1_ASAP7_75t_SL g1970 ( 
.A(n_1926),
.B(n_1884),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1924),
.B(n_1918),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1925),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1942),
.B(n_1914),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1922),
.Y(n_1974)
);

INVxp67_ASAP7_75t_L g1975 ( 
.A(n_1932),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1942),
.B(n_1887),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1921),
.B(n_1918),
.Y(n_1977)
);

AND2x4_ASAP7_75t_L g1978 ( 
.A(n_1926),
.B(n_1893),
.Y(n_1978)
);

AOI221xp5_ASAP7_75t_L g1979 ( 
.A1(n_1941),
.A2(n_1882),
.B1(n_1889),
.B2(n_1912),
.C(n_1913),
.Y(n_1979)
);

NAND2xp33_ASAP7_75t_L g1980 ( 
.A(n_1928),
.B(n_1913),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1948),
.B(n_1887),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1948),
.B(n_1887),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1950),
.B(n_1894),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1925),
.Y(n_1984)
);

OAI21xp33_ASAP7_75t_L g1985 ( 
.A1(n_1937),
.A2(n_1889),
.B(n_1851),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1935),
.B(n_1912),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1937),
.B(n_1929),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1939),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1950),
.B(n_1894),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1939),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1940),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1940),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1947),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1947),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1930),
.Y(n_1995)
);

INVxp67_ASAP7_75t_SL g1996 ( 
.A(n_1963),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1954),
.B(n_1903),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1952),
.Y(n_1998)
);

INVxp67_ASAP7_75t_SL g1999 ( 
.A(n_1934),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1952),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1956),
.Y(n_2001)
);

NOR2x1_ASAP7_75t_L g2002 ( 
.A(n_1926),
.B(n_1797),
.Y(n_2002)
);

INVx3_ASAP7_75t_SL g2003 ( 
.A(n_1927),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1927),
.B(n_1894),
.Y(n_2004)
);

AOI21xp33_ASAP7_75t_SL g2005 ( 
.A1(n_1949),
.A2(n_1868),
.B(n_1880),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1956),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_2003),
.B(n_1961),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1975),
.B(n_1929),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1970),
.Y(n_2009)
);

INVx1_ASAP7_75t_SL g2010 ( 
.A(n_2003),
.Y(n_2010)
);

NOR2xp67_ASAP7_75t_SL g2011 ( 
.A(n_1995),
.B(n_1657),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_2000),
.Y(n_2012)
);

NOR2xp33_ASAP7_75t_L g2013 ( 
.A(n_1969),
.B(n_1946),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_2000),
.Y(n_2014)
);

OR2x2_ASAP7_75t_L g2015 ( 
.A(n_1996),
.B(n_1954),
.Y(n_2015)
);

INVx1_ASAP7_75t_SL g2016 ( 
.A(n_2002),
.Y(n_2016)
);

AOI22xp5_ASAP7_75t_L g2017 ( 
.A1(n_1980),
.A2(n_1933),
.B1(n_1927),
.B2(n_1953),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1979),
.B(n_1977),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1972),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_2006),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1970),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1984),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1988),
.Y(n_2023)
);

AOI22xp33_ASAP7_75t_L g2024 ( 
.A1(n_1980),
.A2(n_1927),
.B1(n_1821),
.B2(n_1943),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1967),
.B(n_1938),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2004),
.B(n_1961),
.Y(n_2026)
);

INVxp67_ASAP7_75t_L g2027 ( 
.A(n_1966),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_2004),
.B(n_1951),
.Y(n_2028)
);

INVx4_ASAP7_75t_L g2029 ( 
.A(n_1968),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1968),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1986),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1990),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1991),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1992),
.Y(n_2034)
);

AND2x4_ASAP7_75t_L g2035 ( 
.A(n_1968),
.B(n_1958),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1973),
.B(n_1951),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2012),
.Y(n_2037)
);

OAI21xp33_ASAP7_75t_SL g2038 ( 
.A1(n_2017),
.A2(n_1968),
.B(n_1999),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2012),
.Y(n_2039)
);

AOI221xp5_ASAP7_75t_L g2040 ( 
.A1(n_2018),
.A2(n_1985),
.B1(n_2005),
.B2(n_1987),
.C(n_1971),
.Y(n_2040)
);

NOR2xp67_ASAP7_75t_L g2041 ( 
.A(n_2021),
.B(n_1974),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_2014),
.Y(n_2042)
);

AOI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_2016),
.A2(n_1974),
.B1(n_1953),
.B2(n_1978),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_2029),
.B(n_2010),
.Y(n_2044)
);

HB1xp67_ASAP7_75t_L g2045 ( 
.A(n_2009),
.Y(n_2045)
);

OAI31xp33_ASAP7_75t_L g2046 ( 
.A1(n_2009),
.A2(n_1978),
.A3(n_1898),
.B(n_1909),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_2015),
.B(n_1997),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_2013),
.B(n_1978),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2031),
.B(n_1983),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_2026),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_L g2051 ( 
.A(n_2029),
.B(n_2030),
.C(n_2008),
.Y(n_2051)
);

NAND2x1p5_ASAP7_75t_L g2052 ( 
.A(n_2029),
.B(n_1664),
.Y(n_2052)
);

OAI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2024),
.A2(n_1888),
.B1(n_1898),
.B2(n_1864),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_2014),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_2028),
.B(n_1973),
.Y(n_2055)
);

AOI211x1_ASAP7_75t_L g2056 ( 
.A1(n_2011),
.A2(n_1976),
.B(n_1982),
.C(n_1981),
.Y(n_2056)
);

AOI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_2011),
.A2(n_1965),
.B1(n_1958),
.B2(n_1989),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2032),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2032),
.Y(n_2059)
);

OR2x2_ASAP7_75t_L g2060 ( 
.A(n_2047),
.B(n_2015),
.Y(n_2060)
);

BUFx2_ASAP7_75t_L g2061 ( 
.A(n_2044),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2055),
.B(n_2028),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2050),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_L g2064 ( 
.A(n_2045),
.B(n_2027),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2044),
.B(n_2030),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2051),
.B(n_2026),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_2048),
.B(n_2021),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2037),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2043),
.B(n_2036),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2039),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2042),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2049),
.B(n_2025),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_2038),
.B(n_2007),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_2056),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2054),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2061),
.B(n_2040),
.Y(n_2076)
);

INVxp67_ASAP7_75t_SL g2077 ( 
.A(n_2073),
.Y(n_2077)
);

NAND3xp33_ASAP7_75t_SL g2078 ( 
.A(n_2073),
.B(n_2046),
.C(n_2052),
.Y(n_2078)
);

OAI221xp5_ASAP7_75t_SL g2079 ( 
.A1(n_2074),
.A2(n_2046),
.B1(n_2057),
.B2(n_2007),
.C(n_2058),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_2062),
.B(n_2041),
.Y(n_2080)
);

AOI21xp33_ASAP7_75t_SL g2081 ( 
.A1(n_2060),
.A2(n_2052),
.B(n_2053),
.Y(n_2081)
);

O2A1O1Ixp33_ASAP7_75t_L g2082 ( 
.A1(n_2074),
.A2(n_2059),
.B(n_2053),
.C(n_2019),
.Y(n_2082)
);

AOI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2066),
.A2(n_2065),
.B(n_2064),
.Y(n_2083)
);

O2A1O1Ixp33_ASAP7_75t_L g2084 ( 
.A1(n_2067),
.A2(n_2020),
.B(n_2034),
.C(n_2023),
.Y(n_2084)
);

AOI21xp5_ASAP7_75t_L g2085 ( 
.A1(n_2067),
.A2(n_2035),
.B(n_2022),
.Y(n_2085)
);

AOI21xp5_ASAP7_75t_SL g2086 ( 
.A1(n_2068),
.A2(n_2035),
.B(n_2033),
.Y(n_2086)
);

AOI221xp5_ASAP7_75t_SL g2087 ( 
.A1(n_2069),
.A2(n_2033),
.B1(n_2036),
.B2(n_1993),
.C(n_2001),
.Y(n_2087)
);

AOI22xp5_ASAP7_75t_L g2088 ( 
.A1(n_2062),
.A2(n_2035),
.B1(n_1965),
.B2(n_1958),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_2081),
.B(n_2072),
.Y(n_2089)
);

AND2x2_ASAP7_75t_L g2090 ( 
.A(n_2077),
.B(n_2063),
.Y(n_2090)
);

NOR2x1_ASAP7_75t_SL g2091 ( 
.A(n_2078),
.B(n_2070),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_2080),
.B(n_2071),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2082),
.A2(n_2075),
.B(n_1997),
.Y(n_2093)
);

NOR2xp33_ASAP7_75t_L g2094 ( 
.A(n_2076),
.B(n_1994),
.Y(n_2094)
);

OAI221xp5_ASAP7_75t_L g2095 ( 
.A1(n_2079),
.A2(n_1998),
.B1(n_1922),
.B2(n_1981),
.C(n_1982),
.Y(n_2095)
);

OAI21xp33_ASAP7_75t_L g2096 ( 
.A1(n_2088),
.A2(n_1989),
.B(n_1983),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2090),
.Y(n_2097)
);

AND2x2_ASAP7_75t_L g2098 ( 
.A(n_2091),
.B(n_2083),
.Y(n_2098)
);

INVx3_ASAP7_75t_L g2099 ( 
.A(n_2096),
.Y(n_2099)
);

NOR2xp33_ASAP7_75t_R g2100 ( 
.A(n_2092),
.B(n_1724),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2089),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2094),
.Y(n_2102)
);

INVxp67_ASAP7_75t_L g2103 ( 
.A(n_2093),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2095),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_2097),
.Y(n_2105)
);

OAI21xp5_ASAP7_75t_SL g2106 ( 
.A1(n_2103),
.A2(n_2098),
.B(n_2101),
.Y(n_2106)
);

NOR2x1p5_ASAP7_75t_L g2107 ( 
.A(n_2099),
.B(n_2086),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_L g2108 ( 
.A(n_2099),
.B(n_2085),
.Y(n_2108)
);

AND2x4_ASAP7_75t_L g2109 ( 
.A(n_2102),
.B(n_1976),
.Y(n_2109)
);

OAI22xp5_ASAP7_75t_SL g2110 ( 
.A1(n_2103),
.A2(n_2084),
.B1(n_1958),
.B2(n_1965),
.Y(n_2110)
);

NOR3xp33_ASAP7_75t_L g2111 ( 
.A(n_2106),
.B(n_2104),
.C(n_2100),
.Y(n_2111)
);

NAND3xp33_ASAP7_75t_L g2112 ( 
.A(n_2108),
.B(n_2087),
.C(n_1893),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2109),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_2107),
.Y(n_2114)
);

NOR2x1_ASAP7_75t_L g2115 ( 
.A(n_2113),
.B(n_2105),
.Y(n_2115)
);

AND3x1_ASAP7_75t_L g2116 ( 
.A(n_2111),
.B(n_2110),
.C(n_1931),
.Y(n_2116)
);

AOI322xp5_ASAP7_75t_L g2117 ( 
.A1(n_2115),
.A2(n_2114),
.A3(n_2112),
.B1(n_1936),
.B2(n_1965),
.C1(n_1909),
.C2(n_1910),
.Y(n_2117)
);

NAND3xp33_ASAP7_75t_SL g2118 ( 
.A(n_2116),
.B(n_1955),
.C(n_1910),
.Y(n_2118)
);

OR2x2_ASAP7_75t_L g2119 ( 
.A(n_2118),
.B(n_1955),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2117),
.Y(n_2120)
);

OR2x2_ASAP7_75t_L g2121 ( 
.A(n_2119),
.B(n_1943),
.Y(n_2121)
);

HB1xp67_ASAP7_75t_L g2122 ( 
.A(n_2120),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2122),
.B(n_1957),
.Y(n_2123)
);

OAI22xp5_ASAP7_75t_SL g2124 ( 
.A1(n_2121),
.A2(n_1893),
.B1(n_1964),
.B2(n_1957),
.Y(n_2124)
);

OAI221xp5_ASAP7_75t_L g2125 ( 
.A1(n_2123),
.A2(n_1964),
.B1(n_1960),
.B2(n_1959),
.C(n_1945),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2125),
.A2(n_2124),
.B1(n_1904),
.B2(n_1945),
.Y(n_2126)
);

NAND2x1p5_ASAP7_75t_L g2127 ( 
.A(n_2126),
.B(n_1791),
.Y(n_2127)
);

AOI22xp5_ASAP7_75t_L g2128 ( 
.A1(n_2127),
.A2(n_1931),
.B1(n_1960),
.B2(n_1959),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2128),
.A2(n_1919),
.B1(n_1936),
.B2(n_1904),
.Y(n_2129)
);

AOI211xp5_ASAP7_75t_L g2130 ( 
.A1(n_2129),
.A2(n_1919),
.B(n_1915),
.C(n_1962),
.Y(n_2130)
);


endmodule