module fake_ariane_2695_n_2097 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2097);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2097;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_365;
wire n_238;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_2016;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1252;
wire n_1129;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_1),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_213),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_124),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_60),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_113),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_133),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_61),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_112),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_18),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_16),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_103),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_58),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_115),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

BUFx2_ASAP7_75t_L g233 ( 
.A(n_126),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_67),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_84),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_97),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_155),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_19),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_8),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_72),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_147),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_38),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_70),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_69),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_61),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_164),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_10),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_78),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_171),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_191),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_44),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_111),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_120),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_30),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_185),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_59),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_106),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

BUFx2_ASAP7_75t_SL g268 ( 
.A(n_33),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_16),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_136),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_21),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_47),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_35),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_138),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_192),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_142),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_63),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_95),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_22),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_157),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_98),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_143),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_159),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_104),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_199),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_43),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_214),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_123),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_54),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_205),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_73),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_208),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_166),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_109),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_30),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_86),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_13),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_144),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_117),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_11),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_176),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_160),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_128),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_196),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_19),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_0),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_74),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g312 ( 
.A(n_209),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_56),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_183),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_195),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_184),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_188),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_156),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_63),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_22),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_6),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_131),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g324 ( 
.A(n_85),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_25),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_5),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_81),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_150),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_204),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_99),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_114),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_193),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_26),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_1),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_119),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_49),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_3),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_139),
.Y(n_339)
);

BUFx5_ASAP7_75t_L g340 ( 
.A(n_47),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_145),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_168),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_174),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_178),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_2),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_141),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_64),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_42),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_38),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_53),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_194),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_212),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_67),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_59),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_88),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_130),
.Y(n_356)
);

INVxp33_ASAP7_75t_SL g357 ( 
.A(n_167),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_170),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_121),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_181),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_152),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_137),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_9),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_4),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_189),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_108),
.Y(n_366)
);

BUFx8_ASAP7_75t_SL g367 ( 
.A(n_34),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_45),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_46),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_202),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_58),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_40),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_82),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_25),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_29),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_29),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_55),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_92),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_148),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_70),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_206),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_52),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_40),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_66),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_107),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_27),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_163),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_53),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_132),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_125),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_72),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_68),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_27),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_26),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_23),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_101),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_71),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_56),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_127),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_134),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_94),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_89),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_211),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_161),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_200),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_71),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_41),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_210),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_12),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_2),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_77),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_17),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_51),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_54),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_18),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_165),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_62),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_7),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_122),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_179),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_65),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_116),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_32),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_93),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_226),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_226),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_376),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_250),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_250),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_340),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_415),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_234),
.B(n_0),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g439 ( 
.A(n_234),
.B(n_3),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_340),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_367),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_358),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_264),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_340),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_295),
.Y(n_446)
);

INVxp67_ASAP7_75t_SL g447 ( 
.A(n_263),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_233),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_340),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_328),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_263),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_340),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_263),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_340),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_283),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_330),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_299),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_381),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_222),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_263),
.Y(n_460)
);

INVxp67_ASAP7_75t_SL g461 ( 
.A(n_263),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_276),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_268),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_276),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_229),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_232),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_222),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_240),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g469 ( 
.A(n_217),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_241),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_228),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_245),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_259),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_228),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_276),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_359),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_294),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_404),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_265),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_217),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_269),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_320),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_272),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_231),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_274),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_300),
.B(n_6),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_276),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_321),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_281),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_370),
.B(n_7),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_286),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_289),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_231),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_235),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_380),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_247),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_296),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_426),
.B(n_219),
.Y(n_498)
);

OR2x2_ASAP7_75t_L g499 ( 
.A(n_414),
.B(n_8),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_235),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_237),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_304),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_392),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_237),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_309),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_316),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_247),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_243),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_243),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_335),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_337),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_350),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_252),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_368),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_374),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_276),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_365),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_252),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_256),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_382),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_365),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_236),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_220),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_236),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_262),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_220),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_223),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_218),
.Y(n_529)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_223),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_384),
.Y(n_531)
);

BUFx2_ASAP7_75t_SL g532 ( 
.A(n_218),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_258),
.B(n_9),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_390),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_393),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_256),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_325),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_435),
.Y(n_538)
);

OA21x2_ASAP7_75t_L g539 ( 
.A1(n_437),
.A2(n_225),
.B(n_224),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_435),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_447),
.B(n_230),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_452),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_262),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_433),
.B(n_408),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_454),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_475),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_516),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_477),
.B(n_357),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_460),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_258),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_460),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_433),
.B(n_417),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_533),
.B(n_261),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_427),
.B(n_420),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_451),
.B(n_239),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_469),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_516),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_477),
.B(n_357),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_507),
.B(n_293),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_462),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_499),
.B(n_425),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_464),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_523),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_523),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_496),
.B(n_261),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_525),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_431),
.B(n_324),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_445),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_453),
.B(n_249),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_527),
.A2(n_338),
.B1(n_396),
.B2(n_227),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_525),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_526),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_532),
.B(n_307),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_526),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_522),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_532),
.B(n_355),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_461),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_496),
.B(n_324),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_487),
.B(n_257),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_499),
.A2(n_305),
.B(n_293),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_522),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_429),
.Y(n_591)
);

INVx6_ASAP7_75t_L g592 ( 
.A(n_529),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_465),
.Y(n_593)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_457),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_498),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_432),
.B(n_260),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_466),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_469),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_468),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_434),
.B(n_266),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_470),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_443),
.B(n_315),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_473),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g606 ( 
.A(n_488),
.B(n_227),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_481),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_459),
.B(n_305),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_483),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_485),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_491),
.A2(n_331),
.B(n_327),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_497),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_502),
.B(n_267),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_463),
.B(n_402),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_506),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_510),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_511),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_512),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_515),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_531),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_568),
.B(n_489),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_538),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_538),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_540),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_555),
.B(n_559),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_555),
.B(n_327),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_593),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_538),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g633 ( 
.A(n_576),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_595),
.B(n_459),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_567),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_568),
.B(n_520),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_567),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_567),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_573),
.Y(n_640)
);

INVx2_ASAP7_75t_SL g641 ( 
.A(n_576),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_595),
.B(n_467),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_582),
.B(n_467),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_594),
.B(n_537),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_573),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_573),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_592),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_577),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_552),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_577),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_582),
.B(n_471),
.Y(n_652)
);

AOI22xp33_ASAP7_75t_L g653 ( 
.A1(n_555),
.A2(n_490),
.B1(n_486),
.B2(n_430),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_555),
.A2(n_430),
.B1(n_530),
.B2(n_524),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_608),
.B(n_529),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_543),
.Y(n_656)
);

INVxp67_ASAP7_75t_SL g657 ( 
.A(n_543),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_552),
.B(n_471),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

OAI22xp33_ASAP7_75t_L g660 ( 
.A1(n_568),
.A2(n_448),
.B1(n_458),
.B2(n_455),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_554),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_585),
.B(n_474),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_554),
.Y(n_663)
);

OR2x2_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_482),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_576),
.Y(n_665)
);

BUFx10_ASAP7_75t_L g666 ( 
.A(n_564),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_556),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_543),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_543),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_540),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g671 ( 
.A(n_598),
.B(n_436),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_555),
.A2(n_530),
.B1(n_455),
.B2(n_458),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_564),
.B(n_474),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_547),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_585),
.B(n_484),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_559),
.A2(n_448),
.B1(n_438),
.B2(n_439),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_565),
.B(n_484),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_608),
.B(n_493),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_562),
.B(n_493),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_618),
.B(n_534),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_618),
.B(n_535),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_559),
.A2(n_546),
.B1(n_568),
.B2(n_539),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_606),
.Y(n_683)
);

INVxp67_ASAP7_75t_SL g684 ( 
.A(n_547),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_568),
.A2(n_494),
.B1(n_501),
.B2(n_500),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_606),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_559),
.B(n_331),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_592),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_568),
.A2(n_500),
.B1(n_501),
.B2(n_494),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_547),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_556),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_547),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_592),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_547),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_558),
.Y(n_695)
);

INVxp33_ASAP7_75t_L g696 ( 
.A(n_598),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_562),
.B(n_504),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_586),
.B(n_559),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_540),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_544),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_565),
.B(n_504),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_614),
.B(n_508),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_586),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_544),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_545),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_540),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_603),
.B(n_508),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_545),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_617),
.B(n_509),
.Y(n_709)
);

INVx3_ASAP7_75t_L g710 ( 
.A(n_540),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_617),
.B(n_509),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_574),
.B(n_513),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_558),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_614),
.B(n_480),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_549),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_541),
.B(n_513),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_566),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_574),
.B(n_518),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_622),
.B(n_517),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_549),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_540),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_546),
.A2(n_529),
.B1(n_521),
.B2(n_528),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_593),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_546),
.A2(n_536),
.B1(n_519),
.B2(n_518),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_553),
.Y(n_725)
);

INVx5_ASAP7_75t_L g726 ( 
.A(n_546),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_566),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_592),
.B(n_442),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_579),
.B(n_519),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_574),
.B(n_536),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_553),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_574),
.B(n_287),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_540),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_593),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_574),
.B(n_405),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_569),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_542),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_542),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_569),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_542),
.Y(n_740)
);

OR2x6_ASAP7_75t_L g741 ( 
.A(n_560),
.B(n_402),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_550),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_546),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_550),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_592),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_579),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_550),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_587),
.B(n_560),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_546),
.A2(n_428),
.B1(n_406),
.B2(n_326),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_551),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_548),
.A2(n_255),
.B1(n_254),
.B2(n_253),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_551),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_587),
.B(n_315),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_587),
.B(n_387),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_592),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_570),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_551),
.Y(n_757)
);

INVx4_ASAP7_75t_L g758 ( 
.A(n_546),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_546),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_570),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_584),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_587),
.B(n_387),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_563),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_589),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_622),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_560),
.B(n_406),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_589),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_539),
.A2(n_622),
.B1(n_587),
.B2(n_613),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_589),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_611),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_618),
.B(n_238),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_596),
.B(n_271),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_548),
.B(n_557),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_584),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_548),
.B(n_442),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_541),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_584),
.Y(n_777)
);

NAND3xp33_ASAP7_75t_SL g778 ( 
.A(n_557),
.B(n_242),
.C(n_238),
.Y(n_778)
);

NAND2x1p5_ASAP7_75t_L g779 ( 
.A(n_758),
.B(n_618),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_776),
.B(n_618),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_626),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_766),
.B(n_557),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_716),
.B(n_623),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_635),
.B(n_623),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_626),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_L g786 ( 
.A(n_642),
.B(n_578),
.C(n_561),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_633),
.B(n_623),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_633),
.B(n_623),
.Y(n_788)
);

NAND2x1p5_ASAP7_75t_L g789 ( 
.A(n_758),
.B(n_623),
.Y(n_789)
);

AOI221xp5_ASAP7_75t_L g790 ( 
.A1(n_660),
.A2(n_419),
.B1(n_255),
.B2(n_254),
.C(n_253),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_632),
.Y(n_791)
);

NOR3xp33_ASAP7_75t_L g792 ( 
.A(n_685),
.B(n_599),
.C(n_597),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_641),
.B(n_561),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_664),
.B(n_591),
.Y(n_794)
);

INVx8_ASAP7_75t_L g795 ( 
.A(n_629),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_641),
.B(n_578),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_664),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_665),
.B(n_588),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_643),
.B(n_588),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_652),
.B(n_591),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_662),
.B(n_675),
.Y(n_801)
);

AOI22xp5_ASAP7_75t_L g802 ( 
.A1(n_687),
.A2(n_599),
.B1(n_601),
.B2(n_597),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_632),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_758),
.B(n_605),
.Y(n_804)
);

NOR2x1p5_ASAP7_75t_L g805 ( 
.A(n_671),
.B(n_601),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_687),
.A2(n_682),
.B1(n_766),
.B2(n_630),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_700),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_661),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_677),
.B(n_591),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_700),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_634),
.B(n_605),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_719),
.Y(n_812)
);

NOR2xp67_ASAP7_75t_L g813 ( 
.A(n_671),
.B(n_602),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_634),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_665),
.B(n_605),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_625),
.B(n_602),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_711),
.B(n_605),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_625),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_629),
.B(n_605),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_634),
.B(n_605),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_704),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_765),
.B(n_605),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_704),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_669),
.Y(n_824)
);

INVxp33_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_701),
.B(n_604),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_663),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_629),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_709),
.B(n_604),
.Y(n_829)
);

BUFx8_ASAP7_75t_L g830 ( 
.A(n_719),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_658),
.B(n_607),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_625),
.B(n_612),
.Y(n_832)
);

AND2x4_ASAP7_75t_L g833 ( 
.A(n_637),
.B(n_607),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_629),
.B(n_612),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_L g835 ( 
.A(n_672),
.B(n_619),
.C(n_612),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_637),
.B(n_612),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_689),
.B(n_616),
.C(n_609),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_637),
.B(n_765),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_743),
.B(n_612),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_629),
.B(n_612),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_705),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_663),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_743),
.B(n_612),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_714),
.B(n_609),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_708),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_708),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_653),
.A2(n_400),
.B1(n_244),
.B2(n_246),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_683),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_629),
.B(n_619),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_667),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_715),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_703),
.B(n_619),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_703),
.B(n_619),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_720),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_667),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_771),
.B(n_619),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_771),
.B(n_619),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_714),
.B(n_696),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_669),
.A2(n_611),
.B(n_615),
.C(n_616),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_720),
.Y(n_860)
);

OAI22x1_ASAP7_75t_L g861 ( 
.A1(n_729),
.A2(n_495),
.B1(n_503),
.B2(n_450),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_725),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_691),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_691),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_695),
.Y(n_865)
);

NOR2xp67_ASAP7_75t_L g866 ( 
.A(n_724),
.B(n_610),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_680),
.B(n_619),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_628),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_695),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_759),
.B(n_391),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_SL g871 ( 
.A(n_746),
.B(n_444),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_731),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_683),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_630),
.A2(n_624),
.B1(n_621),
.B2(n_620),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_673),
.B(n_596),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_766),
.B(n_610),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_669),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_713),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_SL g879 ( 
.A(n_729),
.B(n_446),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_713),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_SL g881 ( 
.A(n_728),
.B(n_242),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_680),
.B(n_610),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_681),
.B(n_772),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_649),
.B(n_615),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_654),
.A2(n_423),
.B1(n_251),
.B2(n_399),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_717),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_678),
.B(n_600),
.Y(n_887)
);

OAI221xp5_ASAP7_75t_L g888 ( 
.A1(n_676),
.A2(n_600),
.B1(n_388),
.B2(n_394),
.C(n_395),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_731),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_719),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_649),
.B(n_613),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_686),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_681),
.B(n_613),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_772),
.B(n_620),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_759),
.B(n_391),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_772),
.B(n_698),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_772),
.B(n_620),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_748),
.B(n_621),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_649),
.B(n_621),
.Y(n_899)
);

INVx2_ASAP7_75t_SL g900 ( 
.A(n_775),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_766),
.A2(n_539),
.B1(n_624),
.B2(n_580),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_657),
.B(n_624),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_684),
.B(n_571),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_737),
.Y(n_904)
);

BUFx5_ASAP7_75t_L g905 ( 
.A(n_764),
.Y(n_905)
);

NAND2x1_ASAP7_75t_L g906 ( 
.A(n_647),
.B(n_539),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_674),
.B(n_403),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_727),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_732),
.B(n_735),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_674),
.B(n_403),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_674),
.B(n_407),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_666),
.B(n_571),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_727),
.Y(n_913)
);

NOR2x1p5_ASAP7_75t_L g914 ( 
.A(n_775),
.B(n_244),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_726),
.B(n_407),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_712),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_726),
.B(n_410),
.Y(n_917)
);

NOR2x1p5_ASAP7_75t_L g918 ( 
.A(n_778),
.B(n_246),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_628),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_666),
.B(n_456),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_656),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_730),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_630),
.B(n_572),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_666),
.B(n_476),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_726),
.B(n_410),
.Y(n_925)
);

AND2x2_ASAP7_75t_SL g926 ( 
.A(n_722),
.B(n_539),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_707),
.A2(n_248),
.B1(n_251),
.B2(n_388),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_630),
.B(n_572),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_741),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_630),
.B(n_575),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_718),
.B(n_575),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_630),
.B(n_580),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_773),
.B(n_478),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_726),
.Y(n_934)
);

NOR3xp33_ASAP7_75t_L g935 ( 
.A(n_679),
.B(n_394),
.C(n_248),
.Y(n_935)
);

AND2x6_ASAP7_75t_L g936 ( 
.A(n_764),
.B(n_580),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_738),
.Y(n_937)
);

NAND2x1_ASAP7_75t_L g938 ( 
.A(n_647),
.B(n_581),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_736),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_768),
.B(n_581),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_739),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_741),
.B(n_581),
.Y(n_942)
);

OR2x6_ASAP7_75t_L g943 ( 
.A(n_741),
.B(n_590),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_741),
.B(n_583),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_783),
.A2(n_769),
.B(n_767),
.Y(n_945)
);

HB1xp67_ASAP7_75t_L g946 ( 
.A(n_797),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_818),
.A2(n_697),
.B1(n_702),
.B2(n_655),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_808),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_817),
.A2(n_769),
.B(n_767),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_SL g950 ( 
.A1(n_826),
.A2(n_754),
.B(n_753),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_799),
.B(n_749),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_827),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_848),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_799),
.B(n_762),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_801),
.B(n_631),
.Y(n_955)
);

OAI21xp5_ASAP7_75t_L g956 ( 
.A1(n_859),
.A2(n_659),
.B(n_656),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_801),
.B(n_723),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_816),
.B(n_833),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_797),
.B(n_751),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_826),
.B(n_734),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_784),
.A2(n_706),
.B(n_668),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_856),
.A2(n_668),
.B(n_659),
.Y(n_962)
);

AO21x1_ASAP7_75t_L g963 ( 
.A1(n_891),
.A2(n_899),
.B(n_809),
.Y(n_963)
);

INVx4_ASAP7_75t_L g964 ( 
.A(n_795),
.Y(n_964)
);

BUFx4f_ASAP7_75t_L g965 ( 
.A(n_943),
.Y(n_965)
);

INVx11_ASAP7_75t_L g966 ( 
.A(n_830),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_829),
.A2(n_690),
.B(n_694),
.C(n_692),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_829),
.B(n_638),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_867),
.A2(n_692),
.B(n_690),
.Y(n_969)
);

OAI22xp5_ASAP7_75t_L g970 ( 
.A1(n_806),
.A2(n_694),
.B1(n_756),
.B2(n_739),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_921),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_857),
.A2(n_721),
.B(n_710),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_795),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_875),
.B(n_638),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_921),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_916),
.A2(n_756),
.B(n_760),
.C(n_645),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_781),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_916),
.A2(n_760),
.B(n_648),
.C(n_639),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_780),
.A2(n_688),
.B(n_647),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_816),
.B(n_726),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_922),
.B(n_900),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_922),
.B(n_686),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_842),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_875),
.B(n_639),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_804),
.A2(n_693),
.B(n_688),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_804),
.A2(n_693),
.B(n_688),
.Y(n_986)
);

CKINVDCx8_ASAP7_75t_R g987 ( 
.A(n_873),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_830),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_809),
.B(n_640),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_858),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_902),
.A2(n_745),
.B(n_693),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_811),
.A2(n_755),
.B(n_745),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_811),
.A2(n_820),
.B(n_882),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_805),
.B(n_590),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_912),
.B(n_640),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_820),
.A2(n_893),
.B(n_891),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_785),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_791),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_912),
.B(n_899),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_828),
.B(n_655),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_903),
.A2(n_755),
.B(n_745),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_884),
.A2(n_755),
.B(n_721),
.Y(n_1002)
);

OAI21xp33_ASAP7_75t_L g1003 ( 
.A1(n_927),
.A2(n_399),
.B(n_395),
.Y(n_1003)
);

BUFx3_ASAP7_75t_L g1004 ( 
.A(n_892),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_L g1005 ( 
.A(n_838),
.B(n_710),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_800),
.A2(n_906),
.B(n_938),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_838),
.B(n_710),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_803),
.Y(n_1008)
);

OAI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_819),
.A2(n_770),
.B(n_648),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_834),
.A2(n_770),
.B(n_645),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_793),
.B(n_627),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_840),
.A2(n_646),
.B(n_636),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_812),
.B(n_818),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_800),
.A2(n_733),
.B(n_721),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_796),
.B(n_627),
.Y(n_1015)
);

NOR2xp67_ASAP7_75t_L g1016 ( 
.A(n_786),
.B(n_920),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_806),
.A2(n_761),
.B1(n_733),
.B2(n_636),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_887),
.A2(n_651),
.B(n_650),
.C(n_646),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_904),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_828),
.B(n_833),
.Y(n_1020)
);

CKINVDCx10_ASAP7_75t_R g1021 ( 
.A(n_782),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_795),
.B(n_774),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_849),
.A2(n_733),
.B(n_761),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_933),
.B(n_590),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_887),
.A2(n_651),
.B(n_650),
.C(n_761),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_782),
.A2(n_813),
.B1(n_836),
.B2(n_832),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_822),
.A2(n_670),
.B(n_628),
.Y(n_1027)
);

NOR2x1_ASAP7_75t_L g1028 ( 
.A(n_794),
.B(n_583),
.Y(n_1028)
);

AOI21x1_ASAP7_75t_L g1029 ( 
.A1(n_839),
.A2(n_740),
.B(n_738),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_815),
.A2(n_670),
.B(n_628),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_890),
.B(n_628),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_782),
.A2(n_777),
.B1(n_774),
.B2(n_699),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_787),
.A2(n_699),
.B(n_670),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_924),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_798),
.B(n_740),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_831),
.A2(n_611),
.B(n_752),
.C(n_763),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_909),
.B(n_742),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_788),
.A2(n_699),
.B(n_670),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_L g1039 ( 
.A(n_790),
.B(n_409),
.C(n_400),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_850),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_943),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_831),
.B(n_742),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_844),
.B(n_583),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_866),
.A2(n_747),
.B(n_744),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_855),
.A2(n_699),
.B(n_670),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_926),
.A2(n_752),
.B1(n_744),
.B2(n_763),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_802),
.B(n_931),
.Y(n_1047)
);

AO21x1_ASAP7_75t_L g1048 ( 
.A1(n_870),
.A2(n_303),
.B(n_275),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_863),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_931),
.B(n_792),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_929),
.B(n_879),
.Y(n_1051)
);

OAI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_847),
.A2(n_411),
.B(n_409),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_883),
.B(n_774),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_937),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_943),
.B(n_699),
.Y(n_1055)
);

AO21x1_ASAP7_75t_L g1056 ( 
.A1(n_870),
.A2(n_314),
.B(n_311),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_868),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_839),
.A2(n_750),
.B(n_747),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_888),
.B(n_774),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_792),
.B(n_750),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_896),
.A2(n_865),
.B(n_869),
.C(n_864),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_914),
.B(n_411),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_878),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_807),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_876),
.B(n_757),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_876),
.B(n_757),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_880),
.A2(n_777),
.B(n_774),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_886),
.A2(n_777),
.B(n_333),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_843),
.A2(n_341),
.B(n_332),
.Y(n_1069)
);

INVx5_ASAP7_75t_L g1070 ( 
.A(n_814),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_837),
.B(n_777),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_868),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_843),
.A2(n_343),
.B(n_342),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_837),
.B(n_777),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_810),
.A2(n_823),
.B(n_821),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_908),
.A2(n_351),
.B(n_344),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_942),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_913),
.A2(n_360),
.B(n_361),
.C(n_424),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_939),
.Y(n_1079)
);

INVx11_ASAP7_75t_L g1080 ( 
.A(n_936),
.Y(n_1080)
);

OR2x6_ASAP7_75t_SL g1081 ( 
.A(n_885),
.B(n_412),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_861),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_814),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_825),
.B(n_412),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_941),
.A2(n_389),
.B(n_362),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_944),
.B(n_416),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_852),
.A2(n_398),
.B(n_397),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_853),
.A2(n_401),
.B(n_413),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_898),
.B(n_584),
.Y(n_1089)
);

NAND2x1_ASAP7_75t_L g1090 ( 
.A(n_814),
.B(n_584),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_907),
.A2(n_563),
.B(n_418),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_814),
.B(n_563),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_824),
.B(n_416),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_935),
.A2(n_418),
.B1(n_422),
.B2(n_421),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_907),
.A2(n_421),
.B(n_422),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_868),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_910),
.A2(n_322),
.B(n_273),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_910),
.A2(n_369),
.B(n_348),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_911),
.A2(n_877),
.B(n_824),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_911),
.A2(n_310),
.B(n_349),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_877),
.A2(n_845),
.B(n_841),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_871),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_935),
.A2(n_423),
.B(n_419),
.C(n_386),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_846),
.A2(n_279),
.B(n_383),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_894),
.B(n_292),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_851),
.A2(n_301),
.B(n_313),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_835),
.A2(n_334),
.B1(n_345),
.B2(n_347),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_897),
.B(n_353),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_779),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_854),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_934),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_918),
.B(n_354),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_860),
.A2(n_363),
.B(n_364),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_862),
.A2(n_375),
.B(n_377),
.Y(n_1114)
);

BUFx4f_ASAP7_75t_L g1115 ( 
.A(n_936),
.Y(n_1115)
);

OAI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_901),
.A2(n_789),
.B1(n_779),
.B2(n_926),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_872),
.B(n_216),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_889),
.A2(n_385),
.B(n_379),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_895),
.B(n_270),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_895),
.A2(n_378),
.B(n_373),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_881),
.A2(n_306),
.B1(n_356),
.B2(n_352),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_901),
.B(n_940),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_789),
.A2(n_298),
.B1(n_346),
.B2(n_339),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_923),
.A2(n_930),
.B(n_928),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_874),
.B(n_277),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_919),
.A2(n_297),
.B(n_336),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_932),
.B(n_278),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_915),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_955),
.A2(n_919),
.B(n_905),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_999),
.A2(n_919),
.B1(n_905),
.B2(n_925),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_954),
.A2(n_1050),
.B(n_967),
.C(n_957),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_982),
.B(n_14),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_946),
.B(n_15),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_959),
.B(n_15),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_981),
.B(n_919),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_980),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_958),
.B(n_905),
.Y(n_1137)
);

INVxp33_ASAP7_75t_L g1138 ( 
.A(n_1084),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_960),
.A2(n_905),
.B(n_925),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_965),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1043),
.B(n_936),
.Y(n_1141)
);

AND2x2_ASAP7_75t_L g1142 ( 
.A(n_958),
.B(n_20),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_965),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_990),
.B(n_915),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1024),
.B(n_936),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_964),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1047),
.B(n_936),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_968),
.A2(n_905),
.B(n_917),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_964),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1013),
.B(n_905),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_L g1151 ( 
.A(n_973),
.B(n_934),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_966),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_989),
.A2(n_302),
.B(n_329),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_949),
.A2(n_290),
.B(n_323),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_SL g1155 ( 
.A1(n_1094),
.A2(n_280),
.B1(n_282),
.B2(n_284),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1077),
.B(n_20),
.Y(n_1156)
);

AOI221xp5_ASAP7_75t_L g1157 ( 
.A1(n_1052),
.A2(n_285),
.B1(n_319),
.B2(n_318),
.C(n_317),
.Y(n_1157)
);

NAND2x1p5_ASAP7_75t_L g1158 ( 
.A(n_980),
.B(n_366),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_948),
.Y(n_1159)
);

INVx1_ASAP7_75t_SL g1160 ( 
.A(n_1021),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_994),
.B(n_23),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1103),
.A2(n_1003),
.B(n_1061),
.C(n_950),
.Y(n_1162)
);

NOR3xp33_ASAP7_75t_SL g1163 ( 
.A(n_953),
.B(n_1039),
.C(n_1097),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_SL g1164 ( 
.A1(n_956),
.A2(n_24),
.B(n_28),
.C(n_31),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_974),
.B(n_24),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_R g1166 ( 
.A(n_987),
.B(n_1004),
.Y(n_1166)
);

AO22x1_ASAP7_75t_L g1167 ( 
.A1(n_988),
.A2(n_1051),
.B1(n_1102),
.B2(n_1082),
.Y(n_1167)
);

BUFx12f_ASAP7_75t_L g1168 ( 
.A(n_1034),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_SL g1169 ( 
.A(n_1016),
.B(n_288),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1080),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_976),
.A2(n_366),
.B(n_308),
.C(n_221),
.Y(n_1171)
);

AND2x4_ASAP7_75t_L g1172 ( 
.A(n_973),
.B(n_1041),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_1057),
.B(n_90),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_1020),
.B(n_1026),
.Y(n_1174)
);

AOI222xp33_ASAP7_75t_L g1175 ( 
.A1(n_1081),
.A2(n_366),
.B1(n_308),
.B2(n_221),
.C1(n_34),
.C2(n_35),
.Y(n_1175)
);

AOI22xp5_ASAP7_75t_L g1176 ( 
.A1(n_963),
.A2(n_312),
.B1(n_291),
.B2(n_308),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_L g1177 ( 
.A1(n_947),
.A2(n_1063),
.B1(n_952),
.B2(n_1040),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_949),
.A2(n_945),
.B(n_1001),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_1070),
.Y(n_1179)
);

OR2x6_ASAP7_75t_SL g1180 ( 
.A(n_1062),
.B(n_28),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_995),
.A2(n_31),
.B(n_32),
.C(n_36),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_984),
.A2(n_366),
.B1(n_308),
.B2(n_221),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_983),
.B(n_36),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_945),
.A2(n_366),
.B(n_308),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1049),
.B(n_37),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1078),
.A2(n_37),
.B(n_39),
.C(n_41),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_979),
.A2(n_221),
.B(n_102),
.Y(n_1187)
);

O2A1O1Ixp5_ASAP7_75t_L g1188 ( 
.A1(n_1006),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1079),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1011),
.B(n_1015),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_991),
.A2(n_221),
.B(n_110),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_996),
.A2(n_291),
.B(n_312),
.Y(n_1192)
);

A2O1A1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1059),
.A2(n_312),
.B(n_291),
.C(n_50),
.Y(n_1193)
);

NOR3xp33_ASAP7_75t_L g1194 ( 
.A(n_1112),
.B(n_46),
.C(n_48),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1070),
.B(n_118),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_993),
.A2(n_291),
.B(n_312),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_1070),
.B(n_105),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1014),
.A2(n_129),
.B(n_215),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1037),
.B(n_48),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1070),
.B(n_1109),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1057),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_SL g1202 ( 
.A1(n_1071),
.A2(n_1074),
.B(n_1000),
.C(n_1025),
.Y(n_1202)
);

AND2x2_ASAP7_75t_SL g1203 ( 
.A(n_1115),
.B(n_50),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1033),
.A2(n_135),
.B(n_201),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1086),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1033),
.A2(n_100),
.B(n_197),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1115),
.B(n_312),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1055),
.Y(n_1208)
);

HB1xp67_ASAP7_75t_L g1209 ( 
.A(n_971),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_970),
.A2(n_51),
.B1(n_52),
.B2(n_55),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1038),
.A2(n_140),
.B(n_190),
.Y(n_1211)
);

OR2x6_ASAP7_75t_L g1212 ( 
.A(n_1116),
.B(n_57),
.Y(n_1212)
);

NAND2xp33_ASAP7_75t_R g1213 ( 
.A(n_1119),
.B(n_1083),
.Y(n_1213)
);

AO21x2_ASAP7_75t_L g1214 ( 
.A1(n_1036),
.A2(n_312),
.B(n_291),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1110),
.A2(n_312),
.B1(n_291),
.B2(n_62),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1057),
.Y(n_1216)
);

AND2x6_ASAP7_75t_L g1217 ( 
.A(n_1083),
.B(n_312),
.Y(n_1217)
);

A2O1A1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_978),
.A2(n_291),
.B(n_60),
.C(n_64),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1093),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_1032),
.B(n_291),
.Y(n_1220)
);

OR2x2_ASAP7_75t_SL g1221 ( 
.A(n_1105),
.B(n_57),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1108),
.B(n_65),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1005),
.A2(n_66),
.B1(n_68),
.B2(n_75),
.Y(n_1223)
);

O2A1O1Ixp5_ASAP7_75t_SL g1224 ( 
.A1(n_1053),
.A2(n_76),
.B(n_79),
.C(n_83),
.Y(n_1224)
);

INVxp67_ASAP7_75t_L g1225 ( 
.A(n_1104),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1128),
.A2(n_91),
.B(n_96),
.C(n_146),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1072),
.Y(n_1227)
);

A2O1A1Ixp33_ASAP7_75t_L g1228 ( 
.A1(n_1076),
.A2(n_149),
.B(n_151),
.C(n_153),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1107),
.B(n_154),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1076),
.A2(n_162),
.B(n_173),
.C(n_180),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1007),
.A2(n_186),
.B1(n_187),
.B2(n_1060),
.Y(n_1231)
);

NOR3xp33_ASAP7_75t_L g1232 ( 
.A(n_1097),
.B(n_1100),
.C(n_1098),
.Y(n_1232)
);

NOR3xp33_ASAP7_75t_SL g1233 ( 
.A(n_1098),
.B(n_1100),
.C(n_1095),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1035),
.B(n_1042),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_975),
.B(n_1121),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_SL g1236 ( 
.A(n_1096),
.B(n_1122),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1028),
.B(n_1085),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1065),
.B(n_1066),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_SL g1239 ( 
.A1(n_1044),
.A2(n_1010),
.B(n_1009),
.C(n_1075),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1104),
.A2(n_1106),
.B(n_1113),
.C(n_1114),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1085),
.A2(n_1069),
.B(n_1073),
.C(n_1099),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1096),
.B(n_1072),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_977),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1099),
.A2(n_1072),
.B1(n_1095),
.B2(n_1031),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1106),
.B(n_1113),
.Y(n_1245)
);

HB1xp67_ASAP7_75t_L g1246 ( 
.A(n_997),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1111),
.B(n_1092),
.Y(n_1247)
);

OAI22x1_ASAP7_75t_L g1248 ( 
.A1(n_998),
.A2(n_1054),
.B1(n_1008),
.B2(n_1019),
.Y(n_1248)
);

BUFx6f_ASAP7_75t_L g1249 ( 
.A(n_1092),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1017),
.A2(n_1125),
.B1(n_1124),
.B2(n_1117),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1123),
.B(n_1111),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1068),
.A2(n_1091),
.B(n_1101),
.C(n_1088),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1038),
.A2(n_1030),
.B(n_961),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1068),
.B(n_1022),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_969),
.B(n_1018),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1012),
.B(n_962),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1090),
.Y(n_1257)
);

CKINVDCx8_ASAP7_75t_R g1258 ( 
.A(n_1048),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1030),
.A2(n_961),
.B(n_1045),
.Y(n_1259)
);

OR2x6_ASAP7_75t_L g1260 ( 
.A(n_1101),
.B(n_1091),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1127),
.B(n_1120),
.Y(n_1261)
);

AND2x4_ASAP7_75t_L g1262 ( 
.A(n_1058),
.B(n_1046),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1056),
.B(n_1118),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1045),
.A2(n_972),
.B(n_1067),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_969),
.A2(n_972),
.B1(n_1067),
.B2(n_1120),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_1029),
.Y(n_1266)
);

OAI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1023),
.A2(n_1002),
.B1(n_1118),
.B2(n_1089),
.Y(n_1267)
);

INVx4_ASAP7_75t_L g1268 ( 
.A(n_1126),
.Y(n_1268)
);

CKINVDCx11_ASAP7_75t_R g1269 ( 
.A(n_1126),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1087),
.A2(n_1088),
.B(n_992),
.C(n_1027),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1087),
.B(n_985),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_986),
.B(n_958),
.Y(n_1272)
);

BUFx4f_ASAP7_75t_L g1273 ( 
.A(n_958),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_982),
.A2(n_746),
.B1(n_933),
.B2(n_729),
.Y(n_1274)
);

BUFx8_ASAP7_75t_L g1275 ( 
.A(n_1004),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_955),
.A2(n_957),
.B(n_960),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_L g1277 ( 
.A(n_1050),
.B(n_564),
.C(n_552),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_964),
.Y(n_1278)
);

AOI22x1_ASAP7_75t_L g1279 ( 
.A1(n_1006),
.A2(n_1099),
.B1(n_961),
.B2(n_969),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_1050),
.A2(n_801),
.B(n_951),
.C(n_826),
.Y(n_1280)
);

INVx2_ASAP7_75t_L g1281 ( 
.A(n_1064),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_955),
.A2(n_957),
.B(n_960),
.Y(n_1282)
);

OAI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1212),
.A2(n_1180),
.B1(n_1258),
.B2(n_1175),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1159),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1277),
.B(n_1138),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1273),
.Y(n_1287)
);

AO21x1_ASAP7_75t_L g1288 ( 
.A1(n_1250),
.A2(n_1162),
.B(n_1276),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1280),
.A2(n_1212),
.B(n_1190),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1140),
.B(n_1143),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1205),
.Y(n_1291)
);

AO31x2_ASAP7_75t_L g1292 ( 
.A1(n_1253),
.A2(n_1264),
.A3(n_1267),
.B(n_1178),
.Y(n_1292)
);

BUFx6f_ASAP7_75t_L g1293 ( 
.A(n_1273),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1274),
.B(n_1142),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1134),
.B(n_1208),
.Y(n_1295)
);

AO21x2_ASAP7_75t_L g1296 ( 
.A1(n_1176),
.A2(n_1261),
.B(n_1214),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1212),
.A2(n_1282),
.B1(n_1203),
.B2(n_1222),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1155),
.A2(n_1269),
.B1(n_1132),
.B2(n_1174),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1165),
.A2(n_1210),
.B1(n_1155),
.B2(n_1221),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1279),
.A2(n_1255),
.B(n_1184),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1189),
.B(n_1219),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1275),
.Y(n_1302)
);

AOI221x1_ASAP7_75t_L g1303 ( 
.A1(n_1193),
.A2(n_1232),
.B1(n_1223),
.B2(n_1218),
.C(n_1194),
.Y(n_1303)
);

NOR2xp67_ASAP7_75t_L g1304 ( 
.A(n_1179),
.B(n_1146),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1196),
.A2(n_1270),
.B(n_1192),
.Y(n_1305)
);

OAI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1239),
.A2(n_1241),
.B(n_1147),
.Y(n_1306)
);

INVx3_ASAP7_75t_L g1307 ( 
.A(n_1179),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1129),
.A2(n_1191),
.B(n_1271),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1131),
.A2(n_1164),
.B(n_1181),
.C(n_1186),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1176),
.A2(n_1225),
.B(n_1139),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1136),
.B(n_1140),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1187),
.A2(n_1148),
.B(n_1244),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1150),
.A2(n_1234),
.B(n_1130),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1171),
.A2(n_1256),
.B(n_1245),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1160),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1246),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_SL g1317 ( 
.A(n_1136),
.B(n_1229),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1263),
.A2(n_1248),
.A3(n_1268),
.B(n_1177),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1133),
.B(n_1160),
.Y(n_1319)
);

AO32x2_ASAP7_75t_L g1320 ( 
.A1(n_1268),
.A2(n_1182),
.A3(n_1231),
.B1(n_1214),
.B2(n_1233),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_SL g1321 ( 
.A1(n_1200),
.A2(n_1262),
.B(n_1256),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1243),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1144),
.B(n_1136),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1135),
.B(n_1140),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1202),
.A2(n_1236),
.B(n_1251),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1236),
.A2(n_1272),
.B(n_1137),
.Y(n_1326)
);

O2A1O1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1240),
.A2(n_1226),
.B(n_1183),
.C(n_1185),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1143),
.B(n_1172),
.Y(n_1328)
);

NOR2xp67_ASAP7_75t_L g1329 ( 
.A(n_1146),
.B(n_1278),
.Y(n_1329)
);

BUFx6f_ASAP7_75t_L g1330 ( 
.A(n_1143),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1204),
.A2(n_1206),
.B(n_1211),
.Y(n_1331)
);

BUFx2_ASAP7_75t_SL g1332 ( 
.A(n_1152),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1198),
.A2(n_1199),
.B(n_1260),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1260),
.A2(n_1141),
.B(n_1262),
.Y(n_1334)
);

AOI221x1_ASAP7_75t_L g1335 ( 
.A1(n_1228),
.A2(n_1230),
.B1(n_1235),
.B2(n_1237),
.C(n_1145),
.Y(n_1335)
);

OAI22x1_ASAP7_75t_L g1336 ( 
.A1(n_1174),
.A2(n_1156),
.B1(n_1169),
.B2(n_1209),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1260),
.A2(n_1254),
.B(n_1153),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1224),
.A2(n_1220),
.B(n_1188),
.Y(n_1338)
);

BUFx2_ASAP7_75t_SL g1339 ( 
.A(n_1170),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1281),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1254),
.A2(n_1207),
.B(n_1154),
.Y(n_1341)
);

O2A1O1Ixp5_ASAP7_75t_L g1342 ( 
.A1(n_1161),
.A2(n_1278),
.B(n_1149),
.C(n_1247),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1254),
.A2(n_1238),
.B(n_1200),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1195),
.A2(n_1242),
.B(n_1158),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1149),
.A2(n_1247),
.B(n_1197),
.Y(n_1345)
);

AOI221x1_ASAP7_75t_L g1346 ( 
.A1(n_1249),
.A2(n_1257),
.B1(n_1201),
.B2(n_1172),
.C(n_1213),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1166),
.B(n_1227),
.Y(n_1347)
);

NOR2x1_ASAP7_75t_SL g1348 ( 
.A(n_1201),
.B(n_1216),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_SL g1349 ( 
.A(n_1249),
.B(n_1201),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1215),
.A2(n_1197),
.B(n_1163),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1170),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1173),
.A2(n_1151),
.B(n_1217),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1167),
.B(n_1249),
.Y(n_1353)
);

INVx5_ASAP7_75t_L g1354 ( 
.A(n_1168),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1275),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1157),
.B(n_1217),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1217),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_1217),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1151),
.A2(n_1282),
.B(n_1276),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1257),
.B(n_797),
.Y(n_1360)
);

OR2x2_ASAP7_75t_L g1361 ( 
.A(n_1274),
.B(n_797),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1133),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1274),
.B(n_797),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1277),
.B(n_797),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_1273),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_SL g1369 ( 
.A(n_1175),
.B(n_1277),
.C(n_564),
.Y(n_1369)
);

NOR2xp67_ASAP7_75t_SL g1370 ( 
.A(n_1152),
.B(n_987),
.Y(n_1370)
);

BUFx10_ASAP7_75t_L g1371 ( 
.A(n_1152),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1166),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1277),
.B(n_797),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1166),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1253),
.A2(n_1178),
.B(n_1259),
.Y(n_1376)
);

INVx2_ASAP7_75t_SL g1377 ( 
.A(n_1275),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1277),
.B(n_797),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1277),
.B(n_797),
.Y(n_1381)
);

O2A1O1Ixp33_ASAP7_75t_SL g1382 ( 
.A1(n_1280),
.A2(n_999),
.B(n_1050),
.C(n_954),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1275),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1275),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1136),
.B(n_965),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1273),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_L g1388 ( 
.A(n_1277),
.B(n_982),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1280),
.B(n_1190),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1274),
.B(n_797),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1280),
.B(n_1190),
.Y(n_1393)
);

OAI22xp5_ASAP7_75t_L g1394 ( 
.A1(n_1280),
.A2(n_1212),
.B1(n_1050),
.B2(n_1047),
.Y(n_1394)
);

AO31x2_ASAP7_75t_L g1395 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1136),
.B(n_1140),
.Y(n_1396)
);

AO31x2_ASAP7_75t_L g1397 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1274),
.B(n_797),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1280),
.A2(n_801),
.B(n_826),
.C(n_1222),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1277),
.B(n_797),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1277),
.B(n_797),
.Y(n_1401)
);

BUFx4_ASAP7_75t_SL g1402 ( 
.A(n_1227),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1205),
.Y(n_1403)
);

A2O1A1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1280),
.A2(n_801),
.B(n_826),
.C(n_1222),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1275),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1407)
);

AOI221xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1210),
.A2(n_1280),
.B1(n_1218),
.B2(n_1181),
.C(n_1162),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1277),
.B(n_982),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1410)
);

O2A1O1Ixp5_ASAP7_75t_SL g1411 ( 
.A1(n_1261),
.A2(n_1192),
.B(n_1265),
.C(n_1196),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1277),
.B(n_797),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1136),
.B(n_1140),
.Y(n_1414)
);

NOR4xp25_ASAP7_75t_L g1415 ( 
.A(n_1280),
.B(n_1162),
.C(n_1050),
.D(n_1210),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1417)
);

OAI21xp5_ASAP7_75t_SL g1418 ( 
.A1(n_1175),
.A2(n_564),
.B(n_552),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1419)
);

A2O1A1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1280),
.A2(n_801),
.B(n_826),
.C(n_1222),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1280),
.A2(n_1050),
.B(n_999),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1159),
.Y(n_1424)
);

BUFx10_ASAP7_75t_L g1425 ( 
.A(n_1152),
.Y(n_1425)
);

AO31x2_ASAP7_75t_L g1426 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1280),
.B(n_1190),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1208),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1430)
);

OAI21xp33_ASAP7_75t_L g1431 ( 
.A1(n_1280),
.A2(n_1277),
.B(n_801),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1432)
);

A2O1A1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1280),
.A2(n_801),
.B(n_826),
.C(n_1222),
.Y(n_1433)
);

AOI21xp5_ASAP7_75t_L g1434 ( 
.A1(n_1276),
.A2(n_1282),
.B(n_1280),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1277),
.B(n_797),
.Y(n_1435)
);

AO31x2_ASAP7_75t_L g1436 ( 
.A1(n_1265),
.A2(n_1266),
.A3(n_1252),
.B(n_1259),
.Y(n_1436)
);

BUFx2_ASAP7_75t_R g1437 ( 
.A(n_1227),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1280),
.A2(n_801),
.B(n_826),
.C(n_1222),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1259),
.A2(n_1264),
.B(n_1253),
.Y(n_1439)
);

AOI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1162),
.A2(n_1050),
.B(n_1175),
.Y(n_1440)
);

O2A1O1Ixp5_ASAP7_75t_SL g1441 ( 
.A1(n_1261),
.A2(n_1192),
.B(n_1265),
.C(n_1196),
.Y(n_1441)
);

INVxp67_ASAP7_75t_L g1442 ( 
.A(n_1133),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1175),
.A2(n_1277),
.B1(n_1050),
.B2(n_552),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1274),
.B(n_797),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1437),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1315),
.Y(n_1446)
);

CKINVDCx11_ASAP7_75t_R g1447 ( 
.A(n_1302),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1371),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1285),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1287),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1371),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1283),
.A2(n_1369),
.B1(n_1440),
.B2(n_1443),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1440),
.B1(n_1443),
.B2(n_1299),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1402),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1418),
.A2(n_1409),
.B1(n_1420),
.B2(n_1399),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1299),
.A2(n_1297),
.B1(n_1398),
.B2(n_1392),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1425),
.Y(n_1458)
);

CKINVDCx11_ASAP7_75t_R g1459 ( 
.A(n_1425),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1418),
.A2(n_1404),
.B1(n_1438),
.B2(n_1433),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1297),
.A2(n_1444),
.B1(n_1364),
.B2(n_1294),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1387),
.Y(n_1462)
);

OAI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1394),
.A2(n_1431),
.B1(n_1381),
.B2(n_1435),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1394),
.A2(n_1431),
.B1(n_1380),
.B2(n_1412),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1287),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1361),
.A2(n_1298),
.B1(n_1317),
.B2(n_1422),
.Y(n_1466)
);

INVx5_ASAP7_75t_L g1467 ( 
.A(n_1287),
.Y(n_1467)
);

CKINVDCx11_ASAP7_75t_R g1468 ( 
.A(n_1355),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1372),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1317),
.A2(n_1356),
.B1(n_1422),
.B2(n_1350),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1424),
.Y(n_1471)
);

CKINVDCx11_ASAP7_75t_R g1472 ( 
.A(n_1383),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1293),
.Y(n_1473)
);

CKINVDCx11_ASAP7_75t_R g1474 ( 
.A(n_1385),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1286),
.A2(n_1442),
.B1(n_1363),
.B2(n_1387),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1429),
.B(n_1367),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1389),
.A2(n_1393),
.B1(n_1428),
.B2(n_1288),
.Y(n_1477)
);

BUFx8_ASAP7_75t_SL g1478 ( 
.A(n_1375),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1285),
.Y(n_1479)
);

NAND2x1p5_ASAP7_75t_L g1480 ( 
.A(n_1293),
.B(n_1368),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1374),
.B(n_1400),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1293),
.B(n_1368),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1322),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1301),
.A2(n_1353),
.B1(n_1393),
.B2(n_1428),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1330),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1340),
.Y(n_1486)
);

BUFx2_ASAP7_75t_L g1487 ( 
.A(n_1360),
.Y(n_1487)
);

BUFx2_ASAP7_75t_SL g1488 ( 
.A(n_1354),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1316),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1389),
.A2(n_1350),
.B1(n_1401),
.B2(n_1336),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1324),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1358),
.A2(n_1289),
.B1(n_1352),
.B2(n_1314),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1330),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1323),
.A2(n_1403),
.B1(n_1291),
.B2(n_1384),
.Y(n_1494)
);

INVx2_ASAP7_75t_SL g1495 ( 
.A(n_1347),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1346),
.Y(n_1496)
);

INVx1_ASAP7_75t_SL g1497 ( 
.A(n_1332),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1337),
.A2(n_1325),
.B(n_1359),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1408),
.A2(n_1319),
.B1(n_1368),
.B2(n_1415),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1408),
.A2(n_1415),
.B1(n_1370),
.B2(n_1290),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1318),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1349),
.Y(n_1502)
);

INVx2_ASAP7_75t_SL g1503 ( 
.A(n_1354),
.Y(n_1503)
);

OR2x2_ASAP7_75t_L g1504 ( 
.A(n_1328),
.B(n_1321),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1334),
.A2(n_1391),
.B1(n_1379),
.B2(n_1434),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1382),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1342),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1343),
.Y(n_1508)
);

OAI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1303),
.A2(n_1335),
.B1(n_1365),
.B2(n_1432),
.Y(n_1509)
);

AOI21xp33_ASAP7_75t_L g1510 ( 
.A1(n_1327),
.A2(n_1309),
.B(n_1296),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1348),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1358),
.A2(n_1352),
.B1(n_1314),
.B2(n_1310),
.Y(n_1512)
);

BUFx10_ASAP7_75t_L g1513 ( 
.A(n_1377),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1306),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1362),
.A2(n_1423),
.B1(n_1373),
.B2(n_1430),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1311),
.B(n_1396),
.Y(n_1516)
);

BUFx6f_ASAP7_75t_L g1517 ( 
.A(n_1386),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1306),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1378),
.A2(n_1410),
.B1(n_1421),
.B2(n_1419),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1413),
.A2(n_1310),
.B1(n_1354),
.B2(n_1396),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1311),
.A2(n_1414),
.B1(n_1290),
.B2(n_1313),
.Y(n_1521)
);

INVx4_ASAP7_75t_L g1522 ( 
.A(n_1351),
.Y(n_1522)
);

INVx4_ASAP7_75t_SL g1523 ( 
.A(n_1357),
.Y(n_1523)
);

INVx1_ASAP7_75t_SL g1524 ( 
.A(n_1414),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1339),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1329),
.A2(n_1351),
.B1(n_1333),
.B2(n_1304),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_SL g1527 ( 
.A1(n_1296),
.A2(n_1406),
.B1(n_1386),
.B2(n_1305),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_SL g1528 ( 
.A1(n_1326),
.A2(n_1338),
.B1(n_1331),
.B2(n_1345),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1307),
.Y(n_1529)
);

BUFx8_ASAP7_75t_L g1530 ( 
.A(n_1320),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1329),
.A2(n_1344),
.B1(n_1300),
.B2(n_1376),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1376),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_SL g1533 ( 
.A1(n_1312),
.A2(n_1441),
.B1(n_1411),
.B2(n_1320),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1534)
);

OAI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1341),
.A2(n_1308),
.B(n_1407),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1320),
.A2(n_1416),
.B1(n_1436),
.B2(n_1426),
.Y(n_1536)
);

CKINVDCx6p67_ASAP7_75t_R g1537 ( 
.A(n_1397),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1416),
.B(n_1436),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1366),
.A2(n_1417),
.B1(n_1390),
.B2(n_1405),
.Y(n_1539)
);

BUFx8_ASAP7_75t_L g1540 ( 
.A(n_1416),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1426),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1436),
.Y(n_1542)
);

CKINVDCx11_ASAP7_75t_R g1543 ( 
.A(n_1292),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1292),
.A2(n_1443),
.B1(n_1418),
.B2(n_1409),
.Y(n_1544)
);

INVx4_ASAP7_75t_L g1545 ( 
.A(n_1292),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1427),
.A2(n_1283),
.B1(n_1317),
.B2(n_1297),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1439),
.A2(n_1283),
.B1(n_1175),
.B2(n_1369),
.Y(n_1547)
);

CKINVDCx11_ASAP7_75t_R g1548 ( 
.A(n_1315),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1418),
.A2(n_1443),
.B1(n_1283),
.B2(n_1369),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1284),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1284),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1443),
.A2(n_1418),
.B1(n_1409),
.B2(n_1388),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_SL g1553 ( 
.A1(n_1283),
.A2(n_1317),
.B1(n_1297),
.B2(n_1299),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1284),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_1402),
.Y(n_1555)
);

CKINVDCx16_ASAP7_75t_R g1556 ( 
.A(n_1302),
.Y(n_1556)
);

INVx4_ASAP7_75t_L g1557 ( 
.A(n_1372),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1399),
.A2(n_1420),
.B(n_1404),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1559)
);

BUFx12f_ASAP7_75t_L g1560 ( 
.A(n_1315),
.Y(n_1560)
);

BUFx8_ASAP7_75t_SL g1561 ( 
.A(n_1302),
.Y(n_1561)
);

CKINVDCx6p67_ASAP7_75t_R g1562 ( 
.A(n_1302),
.Y(n_1562)
);

BUFx6f_ASAP7_75t_SL g1563 ( 
.A(n_1355),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1283),
.A2(n_1317),
.B1(n_1297),
.B2(n_1299),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1567)
);

INVx11_ASAP7_75t_L g1568 ( 
.A(n_1402),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_SL g1569 ( 
.A1(n_1298),
.A2(n_1388),
.B1(n_1409),
.B2(n_1221),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1284),
.Y(n_1570)
);

OAI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1418),
.A2(n_1443),
.B1(n_1212),
.B2(n_1369),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1372),
.Y(n_1572)
);

AOI22xp33_ASAP7_75t_L g1573 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1284),
.Y(n_1575)
);

BUFx10_ASAP7_75t_L g1576 ( 
.A(n_1377),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1364),
.B(n_1392),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_SL g1579 ( 
.A1(n_1283),
.A2(n_1317),
.B1(n_1297),
.B2(n_1299),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1284),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1429),
.B(n_1388),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1284),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1315),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1364),
.B(n_1392),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1284),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1372),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1588)
);

AOI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1399),
.A2(n_1420),
.B(n_1404),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1284),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1283),
.A2(n_1175),
.B1(n_1369),
.B2(n_1440),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1295),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1545),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1508),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1540),
.Y(n_1595)
);

AO21x1_ASAP7_75t_L g1596 ( 
.A1(n_1571),
.A2(n_1544),
.B(n_1460),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_1450),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1514),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1518),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1501),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1510),
.A2(n_1536),
.B(n_1509),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1592),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1532),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1481),
.B(n_1476),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1540),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1498),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1537),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1538),
.B(n_1577),
.Y(n_1608)
);

NOR2x1_ASAP7_75t_R g1609 ( 
.A(n_1446),
.B(n_1548),
.Y(n_1609)
);

BUFx12f_ASAP7_75t_L g1610 ( 
.A(n_1447),
.Y(n_1610)
);

HB1xp67_ASAP7_75t_L g1611 ( 
.A(n_1494),
.Y(n_1611)
);

AND2x4_ASAP7_75t_L g1612 ( 
.A(n_1523),
.B(n_1541),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1471),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1550),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1551),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1554),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1561),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1570),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1575),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1559),
.A2(n_1591),
.B1(n_1565),
.B2(n_1588),
.C(n_1567),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1580),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1553),
.A2(n_1579),
.B1(n_1566),
.B2(n_1565),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1463),
.B(n_1464),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1450),
.Y(n_1624)
);

CKINVDCx6p67_ASAP7_75t_R g1625 ( 
.A(n_1563),
.Y(n_1625)
);

INVx3_ASAP7_75t_L g1626 ( 
.A(n_1507),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1558),
.A2(n_1589),
.B(n_1456),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1529),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1479),
.Y(n_1630)
);

NOR2xp33_ASAP7_75t_L g1631 ( 
.A(n_1449),
.B(n_1564),
.Y(n_1631)
);

CKINVDCx20_ASAP7_75t_R g1632 ( 
.A(n_1584),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1583),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1586),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1585),
.B(n_1457),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1523),
.B(n_1479),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1487),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1535),
.A2(n_1519),
.B(n_1515),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1457),
.B(n_1543),
.Y(n_1639)
);

AO21x2_ASAP7_75t_L g1640 ( 
.A1(n_1536),
.A2(n_1509),
.B(n_1534),
.Y(n_1640)
);

INVx2_ASAP7_75t_SL g1641 ( 
.A(n_1590),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1483),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1486),
.Y(n_1643)
);

BUFx6f_ASAP7_75t_L g1644 ( 
.A(n_1542),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1489),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1461),
.B(n_1477),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1530),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1461),
.B(n_1477),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1469),
.Y(n_1649)
);

INVx3_ASAP7_75t_L g1650 ( 
.A(n_1506),
.Y(n_1650)
);

OA21x2_ASAP7_75t_L g1651 ( 
.A1(n_1515),
.A2(n_1505),
.B(n_1539),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1530),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1582),
.B(n_1552),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1505),
.A2(n_1539),
.B(n_1531),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1484),
.Y(n_1655)
);

BUFx3_ASAP7_75t_L g1656 ( 
.A(n_1572),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1512),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1502),
.Y(n_1658)
);

OAI21x1_ASAP7_75t_L g1659 ( 
.A1(n_1531),
.A2(n_1520),
.B(n_1526),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1512),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1454),
.B(n_1453),
.C(n_1549),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1470),
.B(n_1553),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1491),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1523),
.B(n_1520),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1466),
.B(n_1454),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1490),
.A2(n_1547),
.B(n_1466),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1490),
.A2(n_1521),
.B(n_1500),
.Y(n_1667)
);

BUFx3_ASAP7_75t_L g1668 ( 
.A(n_1572),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1527),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_1447),
.Y(n_1670)
);

BUFx3_ASAP7_75t_L g1671 ( 
.A(n_1587),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1527),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1470),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1492),
.Y(n_1674)
);

BUFx3_ASAP7_75t_L g1675 ( 
.A(n_1587),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1492),
.Y(n_1676)
);

OAI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1453),
.A2(n_1591),
.B1(n_1588),
.B2(n_1581),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1566),
.B(n_1579),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1546),
.B(n_1499),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1533),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1571),
.A2(n_1533),
.B(n_1516),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1546),
.B(n_1547),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1559),
.A2(n_1573),
.B(n_1581),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1528),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1462),
.A2(n_1528),
.B(n_1482),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1475),
.B(n_1578),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1567),
.A2(n_1573),
.B1(n_1578),
.B2(n_1574),
.Y(n_1688)
);

OA21x2_ASAP7_75t_L g1689 ( 
.A1(n_1574),
.A2(n_1511),
.B(n_1524),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1495),
.B(n_1485),
.Y(n_1690)
);

OAI21x1_ASAP7_75t_L g1691 ( 
.A1(n_1462),
.A2(n_1480),
.B(n_1482),
.Y(n_1691)
);

BUFx12f_ASAP7_75t_L g1692 ( 
.A(n_1468),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1485),
.B(n_1493),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1569),
.A2(n_1517),
.B1(n_1488),
.B2(n_1445),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1557),
.B(n_1497),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1557),
.B(n_1525),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1503),
.A2(n_1458),
.B(n_1522),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1568),
.Y(n_1698)
);

INVx4_ASAP7_75t_L g1699 ( 
.A(n_1467),
.Y(n_1699)
);

CKINVDCx20_ASAP7_75t_R g1700 ( 
.A(n_1556),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1467),
.Y(n_1701)
);

AND2x4_ASAP7_75t_L g1702 ( 
.A(n_1467),
.B(n_1555),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1563),
.A2(n_1451),
.B1(n_1473),
.B2(n_1465),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1562),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_SL g1705 ( 
.A1(n_1448),
.A2(n_1452),
.B(n_1459),
.Y(n_1705)
);

INVx3_ASAP7_75t_L g1706 ( 
.A(n_1513),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1513),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1576),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1620),
.A2(n_1455),
.B(n_1468),
.C(n_1478),
.Y(n_1709)
);

AOI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1678),
.A2(n_1472),
.B1(n_1474),
.B2(n_1560),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1622),
.A2(n_1688),
.B1(n_1623),
.B2(n_1653),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1637),
.B(n_1608),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1653),
.A2(n_1661),
.B1(n_1677),
.B2(n_1665),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1637),
.B(n_1656),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1602),
.B(n_1641),
.Y(n_1715)
);

AND2x4_ASAP7_75t_L g1716 ( 
.A(n_1656),
.B(n_1668),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1678),
.A2(n_1683),
.B(n_1662),
.C(n_1665),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1611),
.A2(n_1684),
.B(n_1662),
.Y(n_1718)
);

NAND4xp25_ASAP7_75t_L g1719 ( 
.A(n_1687),
.B(n_1694),
.C(n_1680),
.D(n_1683),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1668),
.B(n_1671),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1671),
.B(n_1675),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1684),
.A2(n_1687),
.B(n_1679),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_SL g1723 ( 
.A1(n_1632),
.A2(n_1700),
.B(n_1704),
.C(n_1708),
.Y(n_1723)
);

OAI21x1_ASAP7_75t_L g1724 ( 
.A1(n_1638),
.A2(n_1606),
.B(n_1686),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1684),
.A2(n_1679),
.B(n_1667),
.Y(n_1725)
);

AOI21xp33_ASAP7_75t_L g1726 ( 
.A1(n_1596),
.A2(n_1684),
.B(n_1628),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1667),
.A2(n_1680),
.B(n_1648),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1628),
.A2(n_1596),
.B(n_1601),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1671),
.B(n_1675),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1695),
.B(n_1696),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1639),
.A2(n_1646),
.B1(n_1648),
.B2(n_1666),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1598),
.B(n_1599),
.Y(n_1732)
);

AOI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1655),
.A2(n_1646),
.B1(n_1673),
.B2(n_1685),
.C(n_1631),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1639),
.A2(n_1673),
.B(n_1685),
.C(n_1655),
.Y(n_1734)
);

AOI221xp5_ASAP7_75t_L g1735 ( 
.A1(n_1669),
.A2(n_1672),
.B1(n_1660),
.B2(n_1657),
.C(n_1604),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1666),
.A2(n_1635),
.B1(n_1674),
.B2(n_1676),
.Y(n_1736)
);

A2O1A1Ixp33_ASAP7_75t_L g1737 ( 
.A1(n_1669),
.A2(n_1672),
.B(n_1664),
.C(n_1657),
.Y(n_1737)
);

HB1xp67_ASAP7_75t_L g1738 ( 
.A(n_1658),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1649),
.B(n_1670),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1664),
.A2(n_1660),
.B(n_1676),
.C(n_1674),
.Y(n_1740)
);

BUFx4f_ASAP7_75t_L g1741 ( 
.A(n_1610),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1690),
.B(n_1629),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1613),
.B(n_1614),
.Y(n_1743)
);

AOI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1635),
.A2(n_1659),
.B(n_1664),
.C(n_1609),
.Y(n_1744)
);

OAI22xp5_ASAP7_75t_L g1745 ( 
.A1(n_1666),
.A2(n_1642),
.B1(n_1615),
.B2(n_1616),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1636),
.B(n_1629),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1690),
.B(n_1693),
.Y(n_1747)
);

OA21x2_ASAP7_75t_L g1748 ( 
.A1(n_1638),
.A2(n_1659),
.B(n_1686),
.Y(n_1748)
);

AND2x4_ASAP7_75t_L g1749 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1698),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1615),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1616),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1666),
.A2(n_1601),
.B1(n_1682),
.B2(n_1681),
.Y(n_1753)
);

A2O1A1Ixp33_ASAP7_75t_L g1754 ( 
.A1(n_1647),
.A2(n_1652),
.B(n_1595),
.C(n_1605),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1618),
.A2(n_1619),
.B1(n_1621),
.B2(n_1633),
.Y(n_1755)
);

AO32x1_ASAP7_75t_L g1756 ( 
.A1(n_1708),
.A2(n_1624),
.A3(n_1630),
.B1(n_1598),
.B2(n_1599),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1636),
.B(n_1612),
.Y(n_1757)
);

BUFx3_ASAP7_75t_L g1758 ( 
.A(n_1692),
.Y(n_1758)
);

AO32x2_ASAP7_75t_L g1759 ( 
.A1(n_1663),
.A2(n_1699),
.A3(n_1640),
.B1(n_1645),
.B2(n_1597),
.Y(n_1759)
);

HB1xp67_ASAP7_75t_L g1760 ( 
.A(n_1621),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1594),
.B(n_1640),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1627),
.B(n_1612),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1634),
.B(n_1642),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1634),
.B(n_1643),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1643),
.Y(n_1765)
);

INVx1_ASAP7_75t_SL g1766 ( 
.A(n_1707),
.Y(n_1766)
);

O2A1O1Ixp33_ASAP7_75t_L g1767 ( 
.A1(n_1707),
.A2(n_1682),
.B(n_1706),
.C(n_1697),
.Y(n_1767)
);

BUFx3_ASAP7_75t_L g1768 ( 
.A(n_1692),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1600),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1651),
.A2(n_1691),
.B(n_1650),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1712),
.B(n_1651),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1738),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1751),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1752),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1651),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1760),
.B(n_1765),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1745),
.B(n_1626),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1755),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1755),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1724),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1732),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1748),
.B(n_1651),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1771),
.B(n_1654),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1732),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1722),
.A2(n_1644),
.B1(n_1689),
.B2(n_1682),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1723),
.B(n_1610),
.Y(n_1787)
);

INVxp67_ASAP7_75t_SL g1788 ( 
.A(n_1761),
.Y(n_1788)
);

OAI221xp5_ASAP7_75t_SL g1789 ( 
.A1(n_1728),
.A2(n_1625),
.B1(n_1703),
.B2(n_1626),
.C(n_1605),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1745),
.B(n_1626),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1771),
.B(n_1654),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1746),
.Y(n_1792)
);

BUFx3_ASAP7_75t_L g1793 ( 
.A(n_1758),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1747),
.B(n_1654),
.Y(n_1794)
);

NOR2xp33_ASAP7_75t_L g1795 ( 
.A(n_1768),
.B(n_1609),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1742),
.B(n_1654),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1717),
.A2(n_1650),
.B1(n_1706),
.B2(n_1702),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1730),
.B(n_1650),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1770),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1761),
.B(n_1603),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1764),
.B(n_1630),
.Y(n_1801)
);

NOR2x1_ASAP7_75t_SL g1802 ( 
.A(n_1762),
.B(n_1701),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1715),
.Y(n_1803)
);

BUFx2_ASAP7_75t_L g1804 ( 
.A(n_1746),
.Y(n_1804)
);

OAI22xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1710),
.A2(n_1617),
.B1(n_1702),
.B2(n_1706),
.Y(n_1805)
);

AND2x4_ASAP7_75t_L g1806 ( 
.A(n_1749),
.B(n_1593),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1713),
.A2(n_1689),
.B1(n_1625),
.B2(n_1702),
.Y(n_1807)
);

NAND3xp33_ASAP7_75t_L g1808 ( 
.A(n_1726),
.B(n_1711),
.C(n_1767),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1741),
.Y(n_1809)
);

BUFx3_ASAP7_75t_L g1810 ( 
.A(n_1741),
.Y(n_1810)
);

INVx1_ASAP7_75t_SL g1811 ( 
.A(n_1714),
.Y(n_1811)
);

NAND4xp25_ASAP7_75t_L g1812 ( 
.A(n_1808),
.B(n_1787),
.C(n_1726),
.D(n_1711),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1808),
.B(n_1718),
.C(n_1744),
.Y(n_1813)
);

OR2x2_ASAP7_75t_L g1814 ( 
.A(n_1777),
.B(n_1766),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1799),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1778),
.A2(n_1756),
.B(n_1744),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1794),
.B(n_1753),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1794),
.B(n_1753),
.Y(n_1818)
);

BUFx3_ASAP7_75t_L g1819 ( 
.A(n_1809),
.Y(n_1819)
);

INVx4_ASAP7_75t_L g1820 ( 
.A(n_1809),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1786),
.A2(n_1718),
.B1(n_1725),
.B2(n_1736),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1794),
.B(n_1720),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_L g1823 ( 
.A(n_1779),
.B(n_1719),
.C(n_1733),
.Y(n_1823)
);

NAND2x1_ASAP7_75t_L g1824 ( 
.A(n_1792),
.B(n_1804),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1800),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1775),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1782),
.B(n_1743),
.Y(n_1827)
);

OAI211xp5_ASAP7_75t_L g1828 ( 
.A1(n_1778),
.A2(n_1710),
.B(n_1709),
.C(n_1719),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1782),
.B(n_1763),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1789),
.B(n_1725),
.C(n_1735),
.Y(n_1830)
);

AND2x4_ASAP7_75t_L g1831 ( 
.A(n_1802),
.B(n_1757),
.Y(n_1831)
);

INVx3_ASAP7_75t_L g1832 ( 
.A(n_1781),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1772),
.B(n_1721),
.Y(n_1833)
);

OR2x6_ASAP7_75t_L g1834 ( 
.A(n_1784),
.B(n_1762),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1772),
.B(n_1729),
.Y(n_1835)
);

INVx5_ASAP7_75t_L g1836 ( 
.A(n_1781),
.Y(n_1836)
);

AND2x4_ASAP7_75t_SL g1837 ( 
.A(n_1806),
.B(n_1769),
.Y(n_1837)
);

INVx3_ASAP7_75t_L g1838 ( 
.A(n_1781),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1785),
.B(n_1736),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1796),
.B(n_1716),
.Y(n_1840)
);

OAI21xp33_ASAP7_75t_L g1841 ( 
.A1(n_1779),
.A2(n_1731),
.B(n_1734),
.Y(n_1841)
);

INVxp67_ASAP7_75t_SL g1842 ( 
.A(n_1790),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1796),
.B(n_1716),
.Y(n_1843)
);

NAND3xp33_ASAP7_75t_L g1844 ( 
.A(n_1780),
.B(n_1727),
.C(n_1754),
.Y(n_1844)
);

OAI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1790),
.A2(n_1727),
.B(n_1740),
.C(n_1737),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1776),
.Y(n_1846)
);

HB1xp67_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1776),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1776),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1798),
.B(n_1759),
.Y(n_1850)
);

NAND2x1p5_ASAP7_75t_L g1851 ( 
.A(n_1807),
.B(n_1607),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1792),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1850),
.B(n_1784),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1846),
.Y(n_1854)
);

BUFx2_ASAP7_75t_L g1855 ( 
.A(n_1842),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1850),
.B(n_1804),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1839),
.B(n_1780),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1850),
.B(n_1803),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1815),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1833),
.B(n_1803),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1826),
.Y(n_1861)
);

INVx3_ASAP7_75t_L g1862 ( 
.A(n_1851),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1842),
.B(n_1785),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1833),
.B(n_1784),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1833),
.B(n_1791),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1839),
.B(n_1774),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1835),
.B(n_1791),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1846),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1851),
.Y(n_1869)
);

HB1xp67_ASAP7_75t_L g1870 ( 
.A(n_1826),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1825),
.B(n_1777),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1827),
.B(n_1774),
.Y(n_1872)
);

OR2x2_ASAP7_75t_L g1873 ( 
.A(n_1825),
.B(n_1801),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1835),
.B(n_1822),
.Y(n_1874)
);

AND2x4_ASAP7_75t_L g1875 ( 
.A(n_1834),
.B(n_1783),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1848),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1848),
.Y(n_1877)
);

NOR2xp33_ASAP7_75t_L g1878 ( 
.A(n_1812),
.B(n_1793),
.Y(n_1878)
);

INVx3_ASAP7_75t_L g1879 ( 
.A(n_1851),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1835),
.B(n_1791),
.Y(n_1880)
);

BUFx3_ASAP7_75t_L g1881 ( 
.A(n_1851),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1827),
.B(n_1788),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1822),
.B(n_1852),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1836),
.Y(n_1884)
);

INVxp67_ASAP7_75t_L g1885 ( 
.A(n_1812),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1852),
.B(n_1811),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1836),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1832),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1847),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1848),
.B(n_1849),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1881),
.B(n_1831),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1874),
.B(n_1840),
.Y(n_1892)
);

OR2x2_ASAP7_75t_L g1893 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1885),
.B(n_1844),
.Y(n_1894)
);

BUFx2_ASAP7_75t_SL g1895 ( 
.A(n_1887),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1874),
.B(n_1840),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1874),
.B(n_1840),
.Y(n_1897)
);

AO221x1_ASAP7_75t_L g1898 ( 
.A1(n_1885),
.A2(n_1805),
.B1(n_1797),
.B2(n_1832),
.C(n_1838),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1857),
.B(n_1844),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1883),
.B(n_1864),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1854),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1878),
.B(n_1795),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1857),
.B(n_1829),
.Y(n_1903)
);

INVx2_ASAP7_75t_SL g1904 ( 
.A(n_1886),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1878),
.B(n_1793),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1861),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1881),
.B(n_1793),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1855),
.B(n_1773),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1855),
.B(n_1773),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1889),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1861),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1870),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1890),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1855),
.B(n_1813),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1890),
.Y(n_1915)
);

AOI211xp5_ASAP7_75t_L g1916 ( 
.A1(n_1881),
.A2(n_1828),
.B(n_1813),
.C(n_1816),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1883),
.B(n_1843),
.Y(n_1917)
);

OR2x2_ASAP7_75t_SL g1918 ( 
.A(n_1863),
.B(n_1823),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1881),
.B(n_1831),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1870),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1866),
.B(n_1816),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1859),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1862),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1866),
.B(n_1828),
.Y(n_1924)
);

INVx2_ASAP7_75t_L g1925 ( 
.A(n_1854),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1872),
.B(n_1814),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1883),
.B(n_1843),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1864),
.B(n_1843),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1859),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1859),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1862),
.B(n_1819),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1864),
.B(n_1837),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1889),
.B(n_1830),
.Y(n_1933)
);

AND2x4_ASAP7_75t_L g1934 ( 
.A(n_1862),
.B(n_1831),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1890),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1890),
.Y(n_1936)
);

OR2x2_ASAP7_75t_L g1937 ( 
.A(n_1872),
.B(n_1814),
.Y(n_1937)
);

INVx1_ASAP7_75t_SL g1938 ( 
.A(n_1918),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1924),
.B(n_1860),
.Y(n_1939)
);

INVx3_ASAP7_75t_L g1940 ( 
.A(n_1891),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1894),
.B(n_1820),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1900),
.B(n_1865),
.Y(n_1942)
);

INVx1_ASAP7_75t_SL g1943 ( 
.A(n_1918),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1899),
.B(n_1860),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1916),
.B(n_1860),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1916),
.B(n_1853),
.Y(n_1946)
);

AOI21xp33_ASAP7_75t_SL g1947 ( 
.A1(n_1914),
.A2(n_1705),
.B(n_1887),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1933),
.B(n_1921),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1900),
.B(n_1865),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1910),
.B(n_1853),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1904),
.B(n_1893),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1904),
.B(n_1853),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1893),
.B(n_1853),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1903),
.B(n_1865),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1892),
.B(n_1867),
.Y(n_1955)
);

AOI22xp33_ASAP7_75t_SL g1956 ( 
.A1(n_1898),
.A2(n_1845),
.B1(n_1823),
.B2(n_1879),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1922),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1902),
.B(n_1905),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1892),
.B(n_1867),
.Y(n_1959)
);

AND2x2_ASAP7_75t_L g1960 ( 
.A(n_1896),
.B(n_1867),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1913),
.Y(n_1961)
);

OR2x6_ASAP7_75t_L g1962 ( 
.A(n_1895),
.B(n_1809),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1913),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1926),
.B(n_1871),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1906),
.B(n_1880),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1907),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1926),
.B(n_1871),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1932),
.B(n_1862),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1913),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1922),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1906),
.B(n_1880),
.Y(n_1972)
);

NOR2x1_ASAP7_75t_L g1973 ( 
.A(n_1895),
.B(n_1810),
.Y(n_1973)
);

NAND3xp33_ASAP7_75t_L g1974 ( 
.A(n_1911),
.B(n_1830),
.C(n_1845),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1896),
.B(n_1880),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1911),
.B(n_1858),
.Y(n_1976)
);

NAND3xp33_ASAP7_75t_L g1977 ( 
.A(n_1956),
.B(n_1920),
.C(n_1912),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1938),
.B(n_1891),
.Y(n_1978)
);

INVxp67_ASAP7_75t_L g1979 ( 
.A(n_1958),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1957),
.Y(n_1980)
);

OR2x6_ASAP7_75t_L g1981 ( 
.A(n_1974),
.B(n_1705),
.Y(n_1981)
);

AOI32xp33_ASAP7_75t_L g1982 ( 
.A1(n_1943),
.A2(n_1946),
.A3(n_1945),
.B1(n_1948),
.B2(n_1939),
.Y(n_1982)
);

OA21x2_ASAP7_75t_L g1983 ( 
.A1(n_1974),
.A2(n_1898),
.B(n_1912),
.Y(n_1983)
);

OAI31xp33_ASAP7_75t_L g1984 ( 
.A1(n_1944),
.A2(n_1841),
.A3(n_1869),
.B(n_1862),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1951),
.B(n_1917),
.Y(n_1985)
);

OAI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1947),
.A2(n_1841),
.B1(n_1821),
.B2(n_1862),
.C(n_1869),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1947),
.B(n_1891),
.Y(n_1987)
);

A2O1A1Ixp33_ASAP7_75t_L g1988 ( 
.A1(n_1941),
.A2(n_1879),
.B(n_1869),
.C(n_1875),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1965),
.B(n_1937),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1973),
.Y(n_1990)
);

AOI22xp5_ASAP7_75t_L g1991 ( 
.A1(n_1967),
.A2(n_1807),
.B1(n_1818),
.B2(n_1817),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1957),
.Y(n_1992)
);

OAI22xp33_ASAP7_75t_L g1993 ( 
.A1(n_1953),
.A2(n_1869),
.B1(n_1879),
.B2(n_1834),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1971),
.Y(n_1994)
);

OAI221xp5_ASAP7_75t_L g1995 ( 
.A1(n_1965),
.A2(n_1879),
.B1(n_1869),
.B2(n_1935),
.C(n_1915),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1971),
.Y(n_1996)
);

INVxp67_ASAP7_75t_L g1997 ( 
.A(n_1973),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1950),
.A2(n_1817),
.B1(n_1818),
.B2(n_1783),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1942),
.B(n_1917),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1942),
.B(n_1927),
.Y(n_2000)
);

INVxp67_ASAP7_75t_L g2001 ( 
.A(n_1962),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_SL g2002 ( 
.A1(n_1962),
.A2(n_1810),
.B(n_1887),
.Y(n_2002)
);

NAND4xp25_ASAP7_75t_SL g2003 ( 
.A(n_1952),
.B(n_1927),
.C(n_1932),
.D(n_1928),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1949),
.B(n_1897),
.Y(n_2004)
);

INVx1_ASAP7_75t_SL g2005 ( 
.A(n_1962),
.Y(n_2005)
);

AOI22xp5_ASAP7_75t_L g2006 ( 
.A1(n_1968),
.A2(n_1817),
.B1(n_1818),
.B2(n_1783),
.Y(n_2006)
);

AOI22xp33_ASAP7_75t_L g2007 ( 
.A1(n_1983),
.A2(n_1875),
.B1(n_1879),
.B2(n_1869),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1999),
.B(n_1940),
.Y(n_2008)
);

OAI21xp5_ASAP7_75t_SL g2009 ( 
.A1(n_1977),
.A2(n_1940),
.B(n_1969),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1983),
.Y(n_2010)
);

OAI221xp5_ASAP7_75t_L g2011 ( 
.A1(n_1984),
.A2(n_1968),
.B1(n_1940),
.B2(n_1879),
.C(n_1962),
.Y(n_2011)
);

OAI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1991),
.A2(n_1954),
.B1(n_1976),
.B2(n_1834),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_2004),
.B(n_1949),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_SL g2014 ( 
.A(n_1982),
.B(n_1920),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1989),
.Y(n_2015)
);

AOI211x1_ASAP7_75t_L g2016 ( 
.A1(n_1986),
.A2(n_1972),
.B(n_1966),
.C(n_1909),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1981),
.B(n_1955),
.Y(n_2017)
);

AOI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1981),
.A2(n_1963),
.B1(n_1970),
.B2(n_1961),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1980),
.Y(n_2019)
);

INVx1_ASAP7_75t_SL g2020 ( 
.A(n_1981),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1992),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1994),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1996),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1979),
.B(n_1955),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1985),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2000),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1978),
.Y(n_2027)
);

OAI21xp33_ASAP7_75t_L g2028 ( 
.A1(n_2003),
.A2(n_1964),
.B(n_1960),
.Y(n_2028)
);

OAI22xp5_ASAP7_75t_L g2029 ( 
.A1(n_1998),
.A2(n_2006),
.B1(n_1990),
.B2(n_1997),
.Y(n_2029)
);

OAI221xp5_ASAP7_75t_L g2030 ( 
.A1(n_2010),
.A2(n_2005),
.B1(n_2001),
.B2(n_1995),
.C(n_1987),
.Y(n_2030)
);

AOI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_2010),
.A2(n_2005),
.B1(n_1993),
.B2(n_1961),
.Y(n_2031)
);

OAI211xp5_ASAP7_75t_L g2032 ( 
.A1(n_2016),
.A2(n_2002),
.B(n_1988),
.C(n_1964),
.Y(n_2032)
);

HB1xp67_ASAP7_75t_L g2033 ( 
.A(n_2015),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2013),
.B(n_1959),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_2015),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2013),
.B(n_1963),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_2024),
.Y(n_2037)
);

NAND2xp33_ASAP7_75t_SL g2038 ( 
.A(n_2017),
.B(n_1908),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2019),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_2008),
.Y(n_2040)
);

NAND4xp75_ASAP7_75t_L g2041 ( 
.A(n_2014),
.B(n_2018),
.C(n_2027),
.D(n_2017),
.Y(n_2041)
);

XOR2x2_ASAP7_75t_L g2042 ( 
.A(n_2014),
.B(n_1810),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_2008),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2025),
.B(n_1970),
.Y(n_2044)
);

NOR2x1_ASAP7_75t_L g2045 ( 
.A(n_2009),
.B(n_1884),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2033),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_2034),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_2043),
.B(n_2020),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_2036),
.B(n_2025),
.Y(n_2049)
);

XNOR2xp5_ASAP7_75t_L g2050 ( 
.A(n_2042),
.B(n_2027),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_2036),
.B(n_2028),
.Y(n_2051)
);

NAND3xp33_ASAP7_75t_L g2052 ( 
.A(n_2035),
.B(n_2007),
.C(n_2029),
.Y(n_2052)
);

NAND4xp25_ASAP7_75t_L g2053 ( 
.A(n_2037),
.B(n_2026),
.C(n_2023),
.D(n_2022),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_2040),
.B(n_2021),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_2030),
.A2(n_2011),
.B(n_1887),
.C(n_1884),
.Y(n_2055)
);

NOR3x1_ASAP7_75t_L g2056 ( 
.A(n_2041),
.B(n_1888),
.C(n_1824),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2044),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_2039),
.B(n_1959),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2047),
.B(n_2044),
.Y(n_2059)
);

NOR3xp33_ASAP7_75t_SL g2060 ( 
.A(n_2053),
.B(n_2051),
.C(n_2030),
.Y(n_2060)
);

NOR2xp33_ASAP7_75t_L g2061 ( 
.A(n_2049),
.B(n_2032),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_R g2062 ( 
.A(n_2046),
.B(n_1750),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_SL g2063 ( 
.A1(n_2052),
.A2(n_2031),
.B1(n_1884),
.B2(n_1923),
.Y(n_2063)
);

AOI211xp5_ASAP7_75t_L g2064 ( 
.A1(n_2055),
.A2(n_2050),
.B(n_2053),
.C(n_2048),
.Y(n_2064)
);

AO22x2_ASAP7_75t_L g2065 ( 
.A1(n_2057),
.A2(n_2038),
.B1(n_1969),
.B2(n_1923),
.Y(n_2065)
);

AOI221xp5_ASAP7_75t_L g2066 ( 
.A1(n_2054),
.A2(n_2012),
.B1(n_1901),
.B2(n_1925),
.C(n_1930),
.Y(n_2066)
);

AO21x1_ASAP7_75t_L g2067 ( 
.A1(n_2061),
.A2(n_2058),
.B(n_2056),
.Y(n_2067)
);

AOI211xp5_ASAP7_75t_L g2068 ( 
.A1(n_2064),
.A2(n_1931),
.B(n_2045),
.C(n_1960),
.Y(n_2068)
);

OAI22xp33_ASAP7_75t_L g2069 ( 
.A1(n_2059),
.A2(n_1884),
.B1(n_1925),
.B2(n_1901),
.Y(n_2069)
);

AOI21xp5_ASAP7_75t_L g2070 ( 
.A1(n_2065),
.A2(n_2063),
.B(n_2066),
.Y(n_2070)
);

NAND4xp25_ASAP7_75t_L g2071 ( 
.A(n_2060),
.B(n_1969),
.C(n_1819),
.D(n_1820),
.Y(n_2071)
);

AOI221xp5_ASAP7_75t_L g2072 ( 
.A1(n_2062),
.A2(n_1930),
.B1(n_1929),
.B2(n_1975),
.C(n_1935),
.Y(n_2072)
);

OAI221xp5_ASAP7_75t_L g2073 ( 
.A1(n_2060),
.A2(n_1923),
.B1(n_1884),
.B2(n_1936),
.C(n_1935),
.Y(n_2073)
);

OAI211xp5_ASAP7_75t_L g2074 ( 
.A1(n_2060),
.A2(n_1923),
.B(n_1884),
.C(n_1820),
.Y(n_2074)
);

NOR2xp67_ASAP7_75t_L g2075 ( 
.A(n_2071),
.B(n_1891),
.Y(n_2075)
);

AO22x1_ASAP7_75t_L g2076 ( 
.A1(n_2067),
.A2(n_1919),
.B1(n_1739),
.B2(n_1934),
.Y(n_2076)
);

NOR2x1p5_ASAP7_75t_L g2077 ( 
.A(n_2074),
.B(n_1819),
.Y(n_2077)
);

OAI211xp5_ASAP7_75t_SL g2078 ( 
.A1(n_2068),
.A2(n_1915),
.B(n_1936),
.C(n_1929),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_2070),
.B(n_1975),
.Y(n_2079)
);

NOR3xp33_ASAP7_75t_L g2080 ( 
.A(n_2073),
.B(n_1820),
.C(n_1915),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2076),
.B(n_2072),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_2075),
.B(n_1897),
.Y(n_2082)
);

NAND3xp33_ASAP7_75t_L g2083 ( 
.A(n_2079),
.B(n_2069),
.C(n_1936),
.Y(n_2083)
);

NAND4xp25_ASAP7_75t_SL g2084 ( 
.A(n_2080),
.B(n_1886),
.C(n_1928),
.D(n_1856),
.Y(n_2084)
);

OAI21xp5_ASAP7_75t_SL g2085 ( 
.A1(n_2081),
.A2(n_2078),
.B(n_2077),
.Y(n_2085)
);

OAI22xp5_ASAP7_75t_L g2086 ( 
.A1(n_2085),
.A2(n_2083),
.B1(n_2082),
.B2(n_2084),
.Y(n_2086)
);

NAND2xp33_ASAP7_75t_R g2087 ( 
.A(n_2086),
.B(n_1919),
.Y(n_2087)
);

OAI22xp5_ASAP7_75t_SL g2088 ( 
.A1(n_2086),
.A2(n_1919),
.B1(n_1934),
.B2(n_1805),
.Y(n_2088)
);

XOR2xp5_ASAP7_75t_L g2089 ( 
.A(n_2088),
.B(n_1919),
.Y(n_2089)
);

AOI22xp5_ASAP7_75t_SL g2090 ( 
.A1(n_2087),
.A2(n_1934),
.B1(n_1858),
.B2(n_1856),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2090),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2089),
.Y(n_2092)
);

AOI21xp5_ASAP7_75t_L g2093 ( 
.A1(n_2091),
.A2(n_1937),
.B(n_1882),
.Y(n_2093)
);

AO21x2_ASAP7_75t_L g2094 ( 
.A1(n_2093),
.A2(n_2092),
.B(n_1882),
.Y(n_2094)
);

OR3x2_ASAP7_75t_L g2095 ( 
.A(n_2094),
.B(n_1871),
.C(n_1873),
.Y(n_2095)
);

OAI221xp5_ASAP7_75t_L g2096 ( 
.A1(n_2095),
.A2(n_1888),
.B1(n_1876),
.B2(n_1868),
.C(n_1877),
.Y(n_2096)
);

AOI211xp5_ASAP7_75t_L g2097 ( 
.A1(n_2096),
.A2(n_1934),
.B(n_1888),
.C(n_1789),
.Y(n_2097)
);


endmodule