module fake_ariane_2509_n_1776 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1776);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1776;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_81),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_28),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_86),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_124),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_106),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g175 ( 
.A(n_93),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_31),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_8),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_125),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_60),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_100),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_60),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_6),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_42),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_104),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_49),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_41),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_168),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_22),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_3),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_49),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_108),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_52),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_90),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_19),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_38),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_35),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_68),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_31),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_37),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_51),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_27),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_24),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_120),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_115),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_57),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_25),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_72),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_55),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_50),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_6),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_9),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_20),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_80),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_61),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_143),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_119),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_63),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_58),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_26),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_30),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_23),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_127),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_45),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_151),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_117),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_51),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_85),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_32),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_65),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_44),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_39),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_70),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_91),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_136),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_7),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_79),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_123),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g256 ( 
.A(n_111),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_164),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_128),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_113),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_163),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_140),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_61),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_154),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_13),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_157),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_18),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_144),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_14),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_102),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_96),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_78),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_107),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_7),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_161),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_40),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_58),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_121),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_56),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_147),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_20),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_2),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_28),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_139),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_97),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_39),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_152),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_137),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_98),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_9),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_29),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_133),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_167),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_69),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_15),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_21),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_153),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_99),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_40),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_130),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_62),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_116),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_26),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_47),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_22),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_73),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_24),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_64),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_25),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_4),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_0),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_32),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_5),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_2),
.Y(n_319)
);

BUFx10_ASAP7_75t_L g320 ( 
.A(n_38),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_33),
.Y(n_321)
);

BUFx10_ASAP7_75t_L g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_36),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_11),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_95),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_103),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_5),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_46),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_57),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_56),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_17),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_82),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_146),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_150),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_12),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_177),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_184),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_195),
.Y(n_339)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_203),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_331),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_170),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_186),
.B(n_1),
.Y(n_343)
);

NOR2xp67_ASAP7_75t_L g344 ( 
.A(n_234),
.B(n_1),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_254),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_268),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_197),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_200),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_234),
.B(n_3),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_266),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_242),
.B(n_4),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_266),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_319),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_266),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_205),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_174),
.B(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_205),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_197),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_197),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_213),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_171),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_213),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_179),
.B(n_10),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_255),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g369 ( 
.A(n_171),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_201),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_225),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_217),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_227),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_262),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_237),
.Y(n_375)
);

INVxp33_ASAP7_75t_SL g376 ( 
.A(n_180),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_223),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_216),
.Y(n_378)
);

BUFx2_ASAP7_75t_SL g379 ( 
.A(n_225),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_225),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_181),
.B(n_10),
.Y(n_381)
);

INVxp33_ASAP7_75t_SL g382 ( 
.A(n_180),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_223),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_283),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_192),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_288),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_216),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_239),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_291),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_247),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_257),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_267),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_288),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_176),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_271),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_280),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_183),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_288),
.Y(n_398)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_284),
.B(n_11),
.Y(n_399)
);

OR2x2_ASAP7_75t_L g400 ( 
.A(n_290),
.B(n_12),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_209),
.B(n_13),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_169),
.Y(n_402)
);

NOR2xp67_ASAP7_75t_L g403 ( 
.A(n_185),
.B(n_15),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_223),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_169),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_295),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_294),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_172),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_320),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_172),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_196),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_296),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_304),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_277),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_194),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_185),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_226),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_315),
.B(n_16),
.Y(n_418)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_365),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_350),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_249),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_394),
.A2(n_306),
.B1(n_243),
.B2(n_308),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_407),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_407),
.B(n_294),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_351),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_411),
.B(n_316),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_385),
.B(n_204),
.Y(n_435)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_365),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_343),
.B(n_178),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_354),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_317),
.Y(n_439)
);

AND2x2_ASAP7_75t_SL g440 ( 
.A(n_367),
.B(n_277),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_212),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_356),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_342),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_342),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_366),
.Y(n_448)
);

OA21x2_ASAP7_75t_L g449 ( 
.A1(n_378),
.A2(n_221),
.B(n_218),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_387),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_353),
.A2(n_276),
.B1(n_248),
.B2(n_228),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_387),
.B(n_229),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_238),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_414),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_357),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_379),
.B(n_324),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_357),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_359),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_379),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_361),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_347),
.B(n_298),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_361),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_363),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_337),
.B(n_244),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_363),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_397),
.A2(n_329),
.B1(n_328),
.B2(n_327),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_346),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_345),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_338),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_339),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_348),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_370),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_372),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_373),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_375),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_388),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_402),
.B(n_214),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_347),
.B(n_298),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_395),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

BUFx8_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_402),
.B(n_256),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_344),
.B(n_253),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_413),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_450),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_440),
.A2(n_349),
.B1(n_358),
.B2(n_401),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_488),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_433),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_444),
.B(n_405),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_485),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_472),
.B(n_360),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_433),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_360),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_437),
.B(n_422),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_420),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_450),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_457),
.B(n_340),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_433),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_433),
.Y(n_509)
);

INVx5_ASAP7_75t_L g510 ( 
.A(n_426),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_SL g511 ( 
.A1(n_468),
.A2(n_355),
.B1(n_404),
.B2(n_409),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_471),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_440),
.A2(n_301),
.B1(n_403),
.B2(n_300),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g515 ( 
.A(n_419),
.B(n_436),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_346),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_433),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_461),
.B(n_405),
.Y(n_518)
);

OR2x2_ASAP7_75t_L g519 ( 
.A(n_419),
.B(n_341),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_485),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_440),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_440),
.A2(n_382),
.B1(n_369),
.B2(n_376),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_457),
.B(n_377),
.Y(n_523)
);

NOR2x1p5_ASAP7_75t_L g524 ( 
.A(n_457),
.B(n_362),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_442),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_436),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_437),
.B(n_362),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_481),
.B(n_408),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_421),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_442),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_481),
.B(n_408),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_423),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_444),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

CKINVDCx8_ASAP7_75t_R g535 ( 
.A(n_444),
.Y(n_535)
);

BUFx8_ASAP7_75t_SL g536 ( 
.A(n_446),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_463),
.B(n_410),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

OAI22xp33_ASAP7_75t_L g539 ( 
.A1(n_452),
.A2(n_383),
.B1(n_399),
.B2(n_400),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_371),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_469),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_452),
.A2(n_418),
.B1(n_399),
.B2(n_400),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_422),
.B(n_371),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_469),
.A2(n_410),
.B1(n_418),
.B2(n_329),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_429),
.Y(n_547)
);

NOR3xp33_ASAP7_75t_L g548 ( 
.A(n_468),
.B(n_190),
.C(n_189),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_450),
.Y(n_549)
);

AND3x1_ASAP7_75t_L g550 ( 
.A(n_473),
.B(n_322),
.C(n_320),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_473),
.B(n_380),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_429),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_485),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_432),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_463),
.B(n_380),
.Y(n_556)
);

NOR3xp33_ASAP7_75t_L g557 ( 
.A(n_446),
.B(n_190),
.C(n_189),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_462),
.Y(n_558)
);

AND3x2_ASAP7_75t_L g559 ( 
.A(n_446),
.B(n_175),
.C(n_260),
.Y(n_559)
);

INVx4_ASAP7_75t_L g560 ( 
.A(n_473),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_434),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_450),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_482),
.B(n_386),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_491),
.A2(n_398),
.B1(n_393),
.B2(n_386),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_470),
.A2(n_208),
.B1(n_207),
.B2(n_202),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_482),
.B(n_393),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_488),
.Y(n_567)
);

AND3x2_ASAP7_75t_L g568 ( 
.A(n_470),
.B(n_274),
.C(n_265),
.Y(n_568)
);

INVx6_ASAP7_75t_L g569 ( 
.A(n_474),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_451),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

NAND3xp33_ASAP7_75t_L g572 ( 
.A(n_489),
.B(n_198),
.C(n_193),
.Y(n_572)
);

BUFx4f_ASAP7_75t_L g573 ( 
.A(n_449),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_473),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_491),
.B(n_191),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_491),
.B(n_246),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_451),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_438),
.Y(n_578)
);

AND2x4_ASAP7_75t_L g579 ( 
.A(n_491),
.B(n_193),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_470),
.B(n_173),
.Y(n_580)
);

INVxp33_ASAP7_75t_L g581 ( 
.A(n_424),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_491),
.B(n_264),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_451),
.Y(n_583)
);

AND2x2_ASAP7_75t_SL g584 ( 
.A(n_489),
.B(n_449),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_476),
.B(n_281),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_488),
.B(n_173),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_430),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_462),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_462),
.Y(n_589)
);

INVx5_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_438),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_430),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_474),
.Y(n_593)
);

AOI22xp33_ASAP7_75t_L g594 ( 
.A1(n_488),
.A2(n_320),
.B1(n_322),
.B2(n_302),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_476),
.B(n_368),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_488),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_475),
.B(n_322),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_451),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_451),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_198),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_449),
.A2(n_230),
.B1(n_252),
.B2(n_245),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_430),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_424),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_451),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_439),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_474),
.B(n_182),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_474),
.B(n_182),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_475),
.B(n_202),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_443),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_474),
.B(n_187),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_443),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_456),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_456),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_456),
.Y(n_615)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_439),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_439),
.B(n_207),
.Y(n_617)
);

CKINVDCx11_ASAP7_75t_R g618 ( 
.A(n_430),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_456),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_462),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_443),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_456),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_462),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_474),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_443),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_462),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_462),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_478),
.B(n_480),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_459),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_480),
.B(n_374),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_430),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_443),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_483),
.Y(n_633)
);

INVx2_ASAP7_75t_SL g634 ( 
.A(n_484),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_443),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_486),
.B(n_187),
.Y(n_636)
);

AND3x2_ASAP7_75t_L g637 ( 
.A(n_486),
.B(n_303),
.C(n_275),
.Y(n_637)
);

BUFx3_ASAP7_75t_L g638 ( 
.A(n_474),
.Y(n_638)
);

NOR3xp33_ASAP7_75t_L g639 ( 
.A(n_487),
.B(n_208),
.C(n_300),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_459),
.Y(n_640)
);

AOI21x1_ASAP7_75t_L g641 ( 
.A1(n_449),
.A2(n_299),
.B(n_313),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_633),
.B(n_477),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_493),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_634),
.B(n_477),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_525),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_525),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_634),
.B(n_477),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_493),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_633),
.B(n_477),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_507),
.B(n_475),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_527),
.B(n_556),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_528),
.B(n_384),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g653 ( 
.A(n_533),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_504),
.B(n_477),
.Y(n_654)
);

A2O1A1Ixp33_ASAP7_75t_L g655 ( 
.A1(n_521),
.A2(n_466),
.B(n_487),
.C(n_492),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_505),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_530),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_505),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_514),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_514),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_633),
.B(n_477),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_521),
.A2(n_321),
.B1(n_308),
.B2(n_309),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_530),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_531),
.B(n_389),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_507),
.B(n_479),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_598),
.B(n_490),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_598),
.B(n_490),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_551),
.B(n_490),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_551),
.B(n_490),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_496),
.B(n_492),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_501),
.B(n_415),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_518),
.B(n_490),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_529),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_R g674 ( 
.A(n_512),
.B(n_417),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_609),
.B(n_490),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_521),
.A2(n_449),
.B1(n_490),
.B2(n_479),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_587),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_529),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_560),
.A2(n_466),
.B(n_453),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_609),
.B(n_523),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_523),
.B(n_479),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_602),
.A2(n_435),
.B1(n_447),
.B2(n_445),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_532),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_532),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_500),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_534),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_503),
.B(n_459),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_587),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_523),
.B(n_459),
.Y(n_690)
);

AND2x2_ASAP7_75t_SL g691 ( 
.A(n_594),
.B(n_292),
.Y(n_691)
);

NAND2x1_ASAP7_75t_L g692 ( 
.A(n_560),
.B(n_426),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_497),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_537),
.B(n_541),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_516),
.B(n_188),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_495),
.B(n_459),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_496),
.B(n_464),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_544),
.B(n_435),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_563),
.B(n_445),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_579),
.B(n_188),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_542),
.B(n_312),
.C(n_309),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_538),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_495),
.B(n_447),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_538),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_566),
.B(n_448),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_580),
.B(n_448),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_579),
.B(n_522),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_533),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_560),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_606),
.B(n_455),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_585),
.B(n_455),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_513),
.A2(n_467),
.B1(n_464),
.B2(n_465),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_500),
.B(n_458),
.Y(n_713)
);

INVx1_ASAP7_75t_SL g714 ( 
.A(n_526),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_497),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_520),
.B(n_458),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_520),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_502),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_595),
.B(n_441),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_553),
.B(n_458),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_441),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_502),
.Y(n_722)
);

CKINVDCx16_ASAP7_75t_R g723 ( 
.A(n_616),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_499),
.B(n_310),
.C(n_312),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_SL g725 ( 
.A(n_535),
.B(n_310),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_547),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_508),
.Y(n_727)
);

BUFx6f_ASAP7_75t_SL g728 ( 
.A(n_579),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_508),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_553),
.B(n_460),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_512),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_547),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_552),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_552),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_564),
.B(n_199),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_509),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_513),
.B(n_460),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_631),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_617),
.B(n_460),
.Y(n_739)
);

NOR2xp67_ASAP7_75t_L g740 ( 
.A(n_515),
.B(n_453),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_575),
.B(n_465),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_465),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_509),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_517),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_515),
.B(n_454),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_558),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_572),
.B(n_454),
.Y(n_747)
);

INVx4_ASAP7_75t_SL g748 ( 
.A(n_631),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_582),
.B(n_467),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_554),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_574),
.B(n_628),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_574),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_617),
.B(n_467),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_517),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_543),
.A2(n_467),
.B1(n_328),
.B2(n_327),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_554),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_613),
.B(n_294),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_555),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_617),
.B(n_467),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_567),
.B(n_467),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_587),
.B(n_199),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_592),
.B(n_206),
.Y(n_763)
);

NOR2xp67_ASAP7_75t_SL g764 ( 
.A(n_574),
.B(n_314),
.Y(n_764)
);

OAI22xp33_ASAP7_75t_L g765 ( 
.A1(n_535),
.A2(n_321),
.B1(n_314),
.B2(n_318),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_613),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_614),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_592),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_592),
.B(n_206),
.Y(n_769)
);

INVxp33_ASAP7_75t_L g770 ( 
.A(n_526),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_614),
.B(n_289),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_615),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_615),
.B(n_619),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_524),
.B(n_318),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_603),
.B(n_289),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_619),
.B(n_293),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_603),
.B(n_293),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_603),
.B(n_297),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_638),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_519),
.B(n_323),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_561),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_557),
.B(n_297),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_622),
.B(n_305),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_622),
.B(n_305),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_519),
.B(n_539),
.Y(n_785)
);

INVx2_ASAP7_75t_SL g786 ( 
.A(n_524),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_629),
.A2(n_325),
.B(n_326),
.C(n_323),
.Y(n_787)
);

INVxp67_ASAP7_75t_L g788 ( 
.A(n_536),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_601),
.B(n_210),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_561),
.Y(n_790)
);

INVx4_ASAP7_75t_L g791 ( 
.A(n_631),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_629),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_596),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_571),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_640),
.Y(n_795)
);

HB1xp67_ASAP7_75t_L g796 ( 
.A(n_565),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_550),
.B(n_307),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_571),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_601),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_640),
.B(n_307),
.Y(n_800)
);

NAND3xp33_ASAP7_75t_SL g801 ( 
.A(n_548),
.B(n_279),
.C(n_236),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_596),
.B(n_311),
.Y(n_802)
);

BUFx8_ASAP7_75t_L g803 ( 
.A(n_558),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_546),
.B(n_211),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_573),
.A2(n_269),
.B1(n_219),
.B2(n_222),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_581),
.B(n_224),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_578),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_578),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_636),
.B(n_311),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_639),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_679),
.A2(n_573),
.B(n_655),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_651),
.A2(n_719),
.B(n_721),
.C(n_785),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_698),
.B(n_584),
.Y(n_813)
);

INVxp67_ASAP7_75t_SL g814 ( 
.A(n_803),
.Y(n_814)
);

BUFx2_ASAP7_75t_L g815 ( 
.A(n_674),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_745),
.A2(n_643),
.B(n_656),
.C(n_648),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_807),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_751),
.A2(n_584),
.B(n_607),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_672),
.A2(n_654),
.B(n_773),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_740),
.B(n_586),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_650),
.B(n_591),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_668),
.A2(n_605),
.B(n_597),
.Y(n_822)
);

INVxp67_ASAP7_75t_L g823 ( 
.A(n_714),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_688),
.A2(n_611),
.B(n_608),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_643),
.A2(n_591),
.B(n_511),
.C(n_600),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_803),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_709),
.B(n_558),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_669),
.A2(n_624),
.B(n_593),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_810),
.B(n_618),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_SL g830 ( 
.A(n_731),
.B(n_604),
.Y(n_830)
);

INVx4_ASAP7_75t_L g831 ( 
.A(n_738),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_650),
.B(n_559),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_648),
.A2(n_506),
.B1(n_599),
.B2(n_494),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_644),
.A2(n_593),
.B(n_624),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_696),
.A2(n_593),
.B(n_624),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_645),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_694),
.B(n_494),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_665),
.B(n_568),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_656),
.A2(n_605),
.B(n_597),
.C(n_600),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_665),
.B(n_494),
.Y(n_840)
);

O2A1O1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_804),
.A2(n_626),
.B(n_627),
.C(n_599),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_645),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_647),
.A2(n_498),
.B(n_599),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_709),
.B(n_558),
.Y(n_844)
);

INVx5_ASAP7_75t_L g845 ( 
.A(n_738),
.Y(n_845)
);

AO21x1_ASAP7_75t_L g846 ( 
.A1(n_703),
.A2(n_570),
.B(n_540),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_739),
.B(n_498),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_680),
.B(n_604),
.Y(n_848)
);

NAND2x1p5_ASAP7_75t_L g849 ( 
.A(n_791),
.B(n_638),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_723),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_709),
.A2(n_506),
.B(n_626),
.Y(n_851)
);

O2A1O1Ixp33_ASAP7_75t_L g852 ( 
.A1(n_662),
.A2(n_796),
.B(n_780),
.C(n_765),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_658),
.A2(n_583),
.B(n_570),
.C(n_562),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_766),
.A2(n_540),
.B(n_549),
.Y(n_854)
);

AOI21x1_ASAP7_75t_L g855 ( 
.A1(n_764),
.A2(n_641),
.B(n_577),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_766),
.A2(n_577),
.B(n_549),
.Y(n_856)
);

INVx1_ASAP7_75t_SL g857 ( 
.A(n_731),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_788),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_653),
.Y(n_859)
);

NOR2x1_ASAP7_75t_L g860 ( 
.A(n_791),
.B(n_626),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_770),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_646),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_658),
.A2(n_627),
.B(n_583),
.C(n_562),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_680),
.B(n_637),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_752),
.B(n_558),
.Y(n_865)
);

O2A1O1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_659),
.A2(n_627),
.B(n_545),
.C(n_610),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_752),
.A2(n_545),
.B(n_635),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_708),
.B(n_235),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_659),
.Y(n_869)
);

BUFx12f_ASAP7_75t_L g870 ( 
.A(n_791),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_660),
.A2(n_610),
.B(n_635),
.C(n_632),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_707),
.B(n_569),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_752),
.A2(n_621),
.B(n_632),
.Y(n_873)
);

OAI21xp5_ASAP7_75t_L g874 ( 
.A1(n_767),
.A2(n_625),
.B(n_621),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_693),
.A2(n_625),
.B(n_612),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_693),
.A2(n_718),
.B(n_715),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_673),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_772),
.A2(n_612),
.B(n_641),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_739),
.B(n_588),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_803),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_801),
.B(n_336),
.C(n_263),
.Y(n_881)
);

BUFx3_ASAP7_75t_L g882 ( 
.A(n_738),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_677),
.B(n_588),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_761),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_673),
.A2(n_427),
.B(n_428),
.C(n_431),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_764),
.A2(n_431),
.B(n_428),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_678),
.A2(n_427),
.B(n_428),
.C(n_431),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_746),
.Y(n_888)
);

OAI21xp5_ASAP7_75t_L g889 ( 
.A1(n_772),
.A2(n_427),
.B(n_335),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_718),
.A2(n_623),
.B(n_620),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_678),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_690),
.B(n_588),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_738),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_690),
.B(n_588),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_711),
.B(n_589),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_710),
.B(n_589),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_671),
.B(n_282),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_677),
.B(n_589),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_761),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_725),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_746),
.Y(n_901)
);

CKINVDCx6p67_ASAP7_75t_R g902 ( 
.A(n_728),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_689),
.B(n_589),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_670),
.B(n_589),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_683),
.A2(n_285),
.B(n_286),
.C(n_287),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_670),
.B(n_706),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_646),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_722),
.A2(n_623),
.B(n_620),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_670),
.B(n_620),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_753),
.B(n_620),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_657),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_770),
.B(n_569),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_792),
.Y(n_913)
);

NOR2xp33_ASAP7_75t_L g914 ( 
.A(n_806),
.B(n_569),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_795),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_761),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_683),
.A2(n_623),
.B1(n_332),
.B2(n_333),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_748),
.B(n_590),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_722),
.A2(n_332),
.B(n_333),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_685),
.A2(n_334),
.B1(n_335),
.B2(n_443),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_768),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_768),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_746),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_727),
.A2(n_334),
.B(n_215),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_795),
.A2(n_426),
.B(n_510),
.Y(n_925)
);

NOR2xp67_ASAP7_75t_L g926 ( 
.A(n_652),
.B(n_590),
.Y(n_926)
);

CKINVDCx6p67_ASAP7_75t_R g927 ( 
.A(n_728),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_753),
.B(n_220),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_806),
.B(n_16),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_760),
.B(n_231),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_727),
.A2(n_261),
.B(n_233),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_685),
.A2(n_759),
.B(n_808),
.C(n_733),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_702),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_747),
.A2(n_675),
.B(n_729),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_760),
.B(n_666),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_686),
.Y(n_936)
);

AOI22x1_ASAP7_75t_L g937 ( 
.A1(n_702),
.A2(n_425),
.B1(n_294),
.B2(n_241),
.Y(n_937)
);

OAI22xp5_ASAP7_75t_L g938 ( 
.A1(n_726),
.A2(n_270),
.B1(n_240),
.B2(n_250),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_664),
.B(n_17),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_689),
.B(n_256),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_697),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_667),
.B(n_699),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_726),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_782),
.B(n_232),
.C(n_251),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_732),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_697),
.Y(n_946)
);

AO21x1_ASAP7_75t_L g947 ( 
.A1(n_732),
.A2(n_256),
.B(n_294),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_733),
.A2(n_273),
.B(n_259),
.C(n_272),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_705),
.B(n_704),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_729),
.A2(n_278),
.B(n_258),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_691),
.B(n_19),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_734),
.B(n_256),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_781),
.B(n_21),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_736),
.A2(n_590),
.B(n_510),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_736),
.A2(n_590),
.B(n_510),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_734),
.B(n_23),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_743),
.A2(n_590),
.B(n_510),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_743),
.A2(n_510),
.B(n_425),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_750),
.B(n_27),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_692),
.A2(n_425),
.B(n_426),
.Y(n_960)
);

AO21x1_ASAP7_75t_L g961 ( 
.A1(n_750),
.A2(n_759),
.B(n_808),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_744),
.A2(n_510),
.B(n_425),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_756),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_756),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_728),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_758),
.B(n_790),
.Y(n_966)
);

OAI21xp33_ASAP7_75t_L g967 ( 
.A1(n_805),
.A2(n_809),
.B(n_784),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_657),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_758),
.B(n_34),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_790),
.A2(n_425),
.B(n_37),
.C(n_43),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_663),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_794),
.B(n_256),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_744),
.A2(n_425),
.B(n_256),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_754),
.A2(n_425),
.B(n_256),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_663),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_748),
.B(n_36),
.Y(n_976)
);

AND3x1_ASAP7_75t_SL g977 ( 
.A(n_794),
.B(n_798),
.C(n_701),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_691),
.B(n_43),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_798),
.B(n_44),
.Y(n_979)
);

AO21x1_ASAP7_75t_L g980 ( 
.A1(n_737),
.A2(n_256),
.B(n_87),
.Y(n_980)
);

AOI21x1_ASAP7_75t_L g981 ( 
.A1(n_692),
.A2(n_426),
.B(n_84),
.Y(n_981)
);

INVx2_ASAP7_75t_SL g982 ( 
.A(n_786),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_787),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_697),
.B(n_48),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_799),
.B(n_48),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_754),
.A2(n_426),
.B(n_92),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_676),
.A2(n_426),
.B(n_89),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_748),
.B(n_50),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_746),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_741),
.B(n_742),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_713),
.A2(n_426),
.B(n_101),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_684),
.Y(n_992)
);

O2A1O1Ixp33_ASAP7_75t_SL g993 ( 
.A1(n_695),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_799),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_681),
.B(n_53),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_642),
.A2(n_426),
.B(n_114),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_812),
.B(n_700),
.Y(n_997)
);

OR2x6_ASAP7_75t_SL g998 ( 
.A(n_858),
.B(n_783),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_848),
.B(n_830),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_812),
.B(n_717),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_823),
.B(n_786),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_813),
.B(n_684),
.Y(n_1002)
);

OR2x6_ASAP7_75t_L g1003 ( 
.A(n_880),
.B(n_686),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_R g1004 ( 
.A(n_815),
.B(n_717),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_819),
.A2(n_649),
.B(n_661),
.Y(n_1005)
);

O2A1O1Ixp5_ASAP7_75t_SL g1006 ( 
.A1(n_952),
.A2(n_797),
.B(n_735),
.C(n_802),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_965),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_951),
.A2(n_755),
.B1(n_682),
.B2(n_712),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_900),
.B(n_774),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_869),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_877),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_990),
.B(n_687),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_951),
.A2(n_774),
.B1(n_789),
.B2(n_724),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_SL g1014 ( 
.A(n_852),
.B(n_789),
.C(n_769),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_891),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_870),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_850),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_933),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_942),
.A2(n_746),
.B(n_730),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_859),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_882),
.Y(n_1021)
);

NOR2xp67_ASAP7_75t_SL g1022 ( 
.A(n_880),
.B(n_762),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_897),
.B(n_763),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_978),
.A2(n_800),
.B1(n_771),
.B2(n_776),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_882),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_913),
.Y(n_1026)
);

INVx6_ASAP7_75t_L g1027 ( 
.A(n_845),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_861),
.B(n_775),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_845),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_949),
.A2(n_716),
.B(n_720),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_966),
.B(n_687),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_978),
.A2(n_778),
.B1(n_777),
.B2(n_793),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_929),
.A2(n_749),
.B(n_779),
.C(n_757),
.Y(n_1033)
);

O2A1O1Ixp33_ASAP7_75t_L g1034 ( 
.A1(n_929),
.A2(n_779),
.B(n_59),
.C(n_62),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_943),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_868),
.B(n_779),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_941),
.B(n_757),
.Y(n_1037)
);

OR2x6_ASAP7_75t_L g1038 ( 
.A(n_826),
.B(n_757),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_845),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_946),
.B(n_757),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_915),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_845),
.Y(n_1042)
);

CKINVDCx11_ASAP7_75t_R g1043 ( 
.A(n_857),
.Y(n_1043)
);

BUFx6f_ASAP7_75t_L g1044 ( 
.A(n_936),
.Y(n_1044)
);

CKINVDCx14_ASAP7_75t_R g1045 ( 
.A(n_902),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_825),
.A2(n_54),
.B(n_59),
.C(n_757),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_945),
.B(n_757),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_835),
.A2(n_940),
.B(n_961),
.C(n_811),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_946),
.B(n_66),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_964),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_836),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_927),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_826),
.B(n_67),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_831),
.B(n_71),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_831),
.Y(n_1055)
);

AND2x2_ASAP7_75t_SL g1056 ( 
.A(n_976),
.B(n_74),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_864),
.B(n_165),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_906),
.B(n_76),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_816),
.A2(n_83),
.B(n_88),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_821),
.B(n_110),
.Y(n_1060)
);

O2A1O1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_825),
.A2(n_122),
.B(n_129),
.C(n_141),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_816),
.B(n_932),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_SL g1063 ( 
.A1(n_932),
.A2(n_142),
.B(n_148),
.C(n_149),
.Y(n_1063)
);

NAND2xp33_ASAP7_75t_R g1064 ( 
.A(n_994),
.B(n_156),
.Y(n_1064)
);

NAND2x1p5_ASAP7_75t_L g1065 ( 
.A(n_918),
.B(n_162),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_893),
.B(n_814),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_895),
.A2(n_837),
.B(n_818),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_837),
.A2(n_873),
.B(n_867),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_936),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_829),
.B(n_832),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_918),
.Y(n_1071)
);

OAI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_967),
.A2(n_939),
.B(n_953),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_884),
.B(n_899),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_827),
.A2(n_865),
.B(n_844),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_935),
.B(n_817),
.Y(n_1075)
);

O2A1O1Ixp5_ASAP7_75t_L g1076 ( 
.A1(n_940),
.A2(n_952),
.B(n_972),
.C(n_846),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_985),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_884),
.B(n_899),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_982),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_984),
.A2(n_959),
.B1(n_969),
.B2(n_956),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_914),
.A2(n_987),
.B(n_872),
.C(n_820),
.Y(n_1081)
);

OAI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_979),
.A2(n_840),
.B1(n_892),
.B2(n_894),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_829),
.B(n_921),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_916),
.B(n_985),
.Y(n_1084)
);

BUFx12f_ASAP7_75t_L g1085 ( 
.A(n_976),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_993),
.A2(n_970),
.B(n_983),
.C(n_963),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_844),
.A2(n_865),
.B(n_828),
.Y(n_1087)
);

A2O1A1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_944),
.A2(n_881),
.B(n_841),
.C(n_824),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_916),
.B(n_914),
.Y(n_1089)
);

BUFx2_ASAP7_75t_L g1090 ( 
.A(n_988),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_912),
.A2(n_838),
.B1(n_977),
.B2(n_872),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_912),
.A2(n_977),
.B1(n_938),
.B2(n_921),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_922),
.B(n_905),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_922),
.B(n_995),
.Y(n_1094)
);

BUFx12f_ASAP7_75t_L g1095 ( 
.A(n_988),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_842),
.B(n_862),
.Y(n_1096)
);

AOI33xp33_ASAP7_75t_L g1097 ( 
.A1(n_993),
.A2(n_970),
.A3(n_887),
.B1(n_885),
.B2(n_866),
.B3(n_863),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_822),
.A2(n_834),
.B(n_851),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_904),
.A2(n_909),
.B1(n_928),
.B2(n_930),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_975),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_888),
.Y(n_1101)
);

O2A1O1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_948),
.A2(n_972),
.B(n_839),
.C(n_917),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_907),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_843),
.A2(n_890),
.B(n_908),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_888),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_883),
.A2(n_898),
.B(n_903),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_911),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_849),
.Y(n_1108)
);

HB1xp67_ASAP7_75t_L g1109 ( 
.A(n_879),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_911),
.Y(n_1110)
);

O2A1O1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_948),
.A2(n_839),
.B(n_847),
.C(n_871),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_888),
.B(n_923),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_910),
.B(n_896),
.Y(n_1113)
);

AO32x1_ASAP7_75t_L g1114 ( 
.A1(n_833),
.A2(n_920),
.A3(n_971),
.B1(n_968),
.B2(n_992),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_968),
.B(n_992),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_853),
.A2(n_878),
.B(n_875),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_854),
.A2(n_874),
.B(n_856),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_876),
.A2(n_934),
.B(n_889),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_919),
.A2(n_924),
.B(n_950),
.C(n_931),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_901),
.B(n_923),
.Y(n_1120)
);

CKINVDCx8_ASAP7_75t_R g1121 ( 
.A(n_901),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_971),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_901),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_980),
.A2(n_991),
.B(n_974),
.C(n_973),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_926),
.A2(n_860),
.B1(n_947),
.B2(n_923),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_SL g1126 ( 
.A1(n_849),
.A2(n_989),
.B1(n_923),
.B2(n_925),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_989),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_989),
.Y(n_1128)
);

OAI22x1_ASAP7_75t_L g1129 ( 
.A1(n_937),
.A2(n_855),
.B1(n_960),
.B2(n_981),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_989),
.B(n_954),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_886),
.Y(n_1131)
);

BUFx2_ASAP7_75t_L g1132 ( 
.A(n_996),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_958),
.B(n_962),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_SL g1134 ( 
.A(n_986),
.B(n_955),
.C(n_957),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_815),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_812),
.A2(n_651),
.B(n_852),
.C(n_951),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_812),
.A2(n_819),
.B(n_813),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_812),
.A2(n_819),
.B(n_813),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_812),
.B(n_535),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_812),
.A2(n_819),
.B(n_813),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_882),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_812),
.A2(n_819),
.B(n_813),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1077),
.B(n_1139),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_L g1144 ( 
.A1(n_1008),
.A2(n_997),
.B1(n_1056),
.B2(n_999),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1136),
.A2(n_1008),
.B(n_1054),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_1080),
.A2(n_1118),
.A3(n_1116),
.B(n_1142),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1137),
.A2(n_1140),
.B(n_1138),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_1020),
.Y(n_1148)
);

AO21x1_ASAP7_75t_L g1149 ( 
.A1(n_1080),
.A2(n_1024),
.B(n_1061),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1067),
.A2(n_1068),
.B(n_1098),
.Y(n_1150)
);

NAND2xp33_ASAP7_75t_SL g1151 ( 
.A(n_1083),
.B(n_1004),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1046),
.A2(n_1072),
.B(n_1086),
.C(n_1024),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1104),
.A2(n_1062),
.B(n_1082),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1010),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1062),
.A2(n_1082),
.B(n_1060),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1070),
.B(n_1009),
.Y(n_1156)
);

BUFx4_ASAP7_75t_SL g1157 ( 
.A(n_1135),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1075),
.B(n_1036),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1090),
.B(n_1023),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1011),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1013),
.A2(n_1032),
.B1(n_1018),
.B2(n_1035),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1081),
.A2(n_1019),
.B(n_1087),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1088),
.A2(n_1000),
.B(n_1049),
.C(n_1093),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1121),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1030),
.A2(n_1117),
.B(n_1005),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1075),
.B(n_1073),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1117),
.A2(n_1133),
.B(n_1012),
.Y(n_1167)
);

OR2x2_ASAP7_75t_L g1168 ( 
.A(n_1069),
.B(n_1015),
.Y(n_1168)
);

AO31x2_ASAP7_75t_L g1169 ( 
.A1(n_1129),
.A2(n_1033),
.A3(n_1002),
.B(n_1113),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1012),
.A2(n_1031),
.B(n_1124),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1028),
.A2(n_1014),
.B1(n_1001),
.B2(n_1084),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1031),
.A2(n_1002),
.B(n_1132),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1073),
.B(n_1071),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_1074),
.A2(n_1096),
.A3(n_1106),
.B(n_1110),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1096),
.A2(n_1122),
.A3(n_1115),
.B(n_1051),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1043),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1134),
.A2(n_1059),
.B(n_1048),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1034),
.A2(n_1102),
.B(n_1091),
.C(n_1094),
.Y(n_1178)
);

AOI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1112),
.A2(n_1037),
.B(n_1040),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1111),
.A2(n_1126),
.B(n_1119),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1050),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_1092),
.B(n_1089),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1076),
.A2(n_1099),
.B(n_1006),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1058),
.A2(n_1089),
.B(n_1047),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1063),
.A2(n_1078),
.B(n_1079),
.C(n_1017),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1125),
.A2(n_1047),
.B(n_1108),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1097),
.A2(n_1130),
.B(n_1120),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1029),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1100),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_1052),
.Y(n_1190)
);

O2A1O1Ixp5_ASAP7_75t_L g1191 ( 
.A1(n_1022),
.A2(n_1130),
.B(n_1128),
.C(n_1127),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1078),
.A2(n_1109),
.B(n_1054),
.Y(n_1192)
);

INVx1_ASAP7_75t_SL g1193 ( 
.A(n_1123),
.Y(n_1193)
);

AOI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1085),
.A2(n_1095),
.B1(n_1057),
.B2(n_1007),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1065),
.A2(n_1103),
.B(n_1107),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1026),
.A2(n_1041),
.B(n_1065),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1044),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_1003),
.B(n_1053),
.Y(n_1198)
);

CKINVDCx11_ASAP7_75t_R g1199 ( 
.A(n_998),
.Y(n_1199)
);

INVx1_ASAP7_75t_SL g1200 ( 
.A(n_1044),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1066),
.B(n_1044),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1066),
.A2(n_1055),
.B(n_1141),
.C(n_1021),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1101),
.B(n_1105),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1114),
.A2(n_1131),
.A3(n_1038),
.B(n_1105),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1038),
.A2(n_1053),
.B(n_1003),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1038),
.A2(n_1053),
.B(n_1114),
.Y(n_1206)
);

BUFx12f_ASAP7_75t_L g1207 ( 
.A(n_1016),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1101),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1045),
.B(n_1141),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1021),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_SL g1211 ( 
.A(n_1025),
.B(n_1029),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1025),
.A2(n_1101),
.B1(n_1027),
.B2(n_1039),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1064),
.A2(n_1027),
.A3(n_1029),
.B(n_1039),
.Y(n_1213)
);

NAND3xp33_ASAP7_75t_L g1214 ( 
.A(n_1042),
.B(n_812),
.C(n_1136),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1042),
.A2(n_1139),
.B1(n_951),
.B2(n_978),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1136),
.A2(n_812),
.B(n_1137),
.Y(n_1216)
);

NAND2xp33_ASAP7_75t_L g1217 ( 
.A(n_1136),
.B(n_812),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1136),
.A2(n_812),
.B(n_1137),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1077),
.B(n_812),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1139),
.B(n_812),
.Y(n_1221)
);

OAI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1136),
.A2(n_812),
.B(n_1137),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1080),
.A2(n_846),
.A3(n_835),
.B(n_980),
.Y(n_1224)
);

OAI21xp33_ASAP7_75t_L g1225 ( 
.A1(n_1136),
.A2(n_812),
.B(n_651),
.Y(n_1225)
);

AO31x2_ASAP7_75t_L g1226 ( 
.A1(n_1080),
.A2(n_846),
.A3(n_835),
.B(n_980),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1139),
.A2(n_725),
.B1(n_785),
.B2(n_951),
.Y(n_1227)
);

AOI22x1_ASAP7_75t_L g1228 ( 
.A1(n_1137),
.A2(n_1140),
.B1(n_1142),
.B2(n_1138),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1010),
.Y(n_1229)
);

AOI221x1_ASAP7_75t_L g1230 ( 
.A1(n_1136),
.A2(n_812),
.B1(n_978),
.B2(n_951),
.C(n_825),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1077),
.B(n_812),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1010),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1010),
.Y(n_1234)
);

AOI221x1_ASAP7_75t_L g1235 ( 
.A1(n_1136),
.A2(n_812),
.B1(n_978),
.B2(n_951),
.C(n_825),
.Y(n_1235)
);

AOI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1129),
.A2(n_1138),
.B(n_1137),
.Y(n_1236)
);

NAND2xp33_ASAP7_75t_L g1237 ( 
.A(n_1136),
.B(n_812),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1139),
.B(n_812),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_SL g1240 ( 
.A1(n_1102),
.A2(n_961),
.B(n_1111),
.Y(n_1240)
);

NOR2xp33_ASAP7_75t_L g1241 ( 
.A(n_1139),
.B(n_812),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1139),
.A2(n_725),
.B1(n_785),
.B2(n_951),
.Y(n_1242)
);

AOI221x1_ASAP7_75t_L g1243 ( 
.A1(n_1136),
.A2(n_812),
.B1(n_978),
.B2(n_951),
.C(n_825),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1139),
.A2(n_812),
.B(n_651),
.C(n_997),
.Y(n_1244)
);

NAND3xp33_ASAP7_75t_L g1245 ( 
.A(n_1136),
.B(n_812),
.C(n_1139),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1043),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1139),
.B(n_812),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1104),
.A2(n_1116),
.B(n_1098),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1080),
.A2(n_846),
.A3(n_835),
.B(n_980),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1136),
.A2(n_812),
.B(n_816),
.C(n_1088),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1136),
.A2(n_812),
.B1(n_1139),
.B2(n_978),
.Y(n_1251)
);

AND2x4_ASAP7_75t_L g1252 ( 
.A(n_1073),
.B(n_882),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_999),
.B(n_848),
.Y(n_1253)
);

AOI31xp67_ASAP7_75t_L g1254 ( 
.A1(n_1133),
.A2(n_1000),
.A3(n_1062),
.B(n_972),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1256)
);

NOR2xp67_ASAP7_75t_L g1257 ( 
.A(n_1135),
.B(n_823),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1136),
.B(n_812),
.Y(n_1258)
);

OAI22x1_ASAP7_75t_L g1259 ( 
.A1(n_1139),
.A2(n_951),
.B1(n_978),
.B2(n_1077),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1077),
.B(n_812),
.Y(n_1260)
);

O2A1O1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1136),
.A2(n_812),
.B(n_651),
.C(n_1139),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1262)
);

NAND2x2_ASAP7_75t_L g1263 ( 
.A(n_1017),
.B(n_601),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1136),
.A2(n_812),
.B(n_1137),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1104),
.A2(n_1116),
.B(n_1098),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_SL g1266 ( 
.A1(n_1136),
.A2(n_812),
.B(n_816),
.C(n_1088),
.Y(n_1266)
);

AOI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1129),
.A2(n_1138),
.B(n_1137),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1043),
.Y(n_1268)
);

INVx3_ASAP7_75t_SL g1269 ( 
.A(n_1135),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_1043),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1139),
.A2(n_725),
.B1(n_785),
.B2(n_951),
.Y(n_1271)
);

CKINVDCx6p67_ASAP7_75t_R g1272 ( 
.A(n_1043),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1139),
.B(n_812),
.Y(n_1273)
);

AND3x2_ASAP7_75t_L g1274 ( 
.A(n_1070),
.B(n_815),
.C(n_725),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1077),
.B(n_812),
.Y(n_1275)
);

BUFx8_ASAP7_75t_L g1276 ( 
.A(n_1020),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1139),
.A2(n_812),
.B(n_651),
.C(n_997),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1043),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1078),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1136),
.A2(n_812),
.B(n_813),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1227),
.A2(n_1271),
.B1(n_1242),
.B2(n_1247),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1159),
.B(n_1253),
.Y(n_1282)
);

CKINVDCx20_ASAP7_75t_R g1283 ( 
.A(n_1246),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1154),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1198),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1160),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1181),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1221),
.A2(n_1238),
.B1(n_1241),
.B2(n_1273),
.Y(n_1288)
);

INVx2_ASAP7_75t_SL g1289 ( 
.A(n_1157),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1229),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1232),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1244),
.B(n_1277),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1234),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1272),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1144),
.A2(n_1251),
.B1(n_1259),
.B2(n_1215),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1258),
.B(n_1251),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1245),
.A2(n_1258),
.B1(n_1225),
.B2(n_1275),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1245),
.A2(n_1261),
.B(n_1235),
.Y(n_1298)
);

BUFx2_ASAP7_75t_L g1299 ( 
.A(n_1276),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1156),
.A2(n_1143),
.B1(n_1278),
.B2(n_1270),
.Y(n_1300)
);

INVx8_ASAP7_75t_L g1301 ( 
.A(n_1198),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1164),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1217),
.A2(n_1237),
.B1(n_1149),
.B2(n_1182),
.Y(n_1303)
);

AOI22xp5_ASAP7_75t_L g1304 ( 
.A1(n_1171),
.A2(n_1161),
.B1(n_1198),
.B2(n_1151),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_1176),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1161),
.A2(n_1206),
.B1(n_1214),
.B2(n_1260),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1230),
.A2(n_1243),
.B1(n_1231),
.B2(n_1194),
.Y(n_1307)
);

OAI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1145),
.A2(n_1280),
.B(n_1223),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1152),
.A2(n_1219),
.B1(n_1255),
.B2(n_1239),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_L g1310 ( 
.A(n_1207),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1279),
.B(n_1220),
.Y(n_1311)
);

OAI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1214),
.A2(n_1166),
.B1(n_1263),
.B2(n_1158),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1276),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1199),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1233),
.B(n_1256),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1178),
.B1(n_1222),
.B2(n_1218),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1268),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1192),
.A2(n_1274),
.B1(n_1205),
.B2(n_1189),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1190),
.Y(n_1319)
);

OAI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1168),
.A2(n_1264),
.B1(n_1222),
.B2(n_1218),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1205),
.A2(n_1206),
.B1(n_1264),
.B2(n_1216),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1148),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1216),
.A2(n_1155),
.B1(n_1153),
.B2(n_1180),
.Y(n_1323)
);

INVx4_ASAP7_75t_R g1324 ( 
.A(n_1209),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1240),
.A2(n_1183),
.B1(n_1196),
.B2(n_1184),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1187),
.A2(n_1177),
.B1(n_1228),
.B2(n_1170),
.Y(n_1326)
);

INVx6_ASAP7_75t_L g1327 ( 
.A(n_1252),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1193),
.B(n_1173),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1183),
.A2(n_1196),
.B1(n_1187),
.B2(n_1257),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1201),
.A2(n_1212),
.B1(n_1173),
.B2(n_1193),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1210),
.A2(n_1172),
.B1(n_1186),
.B2(n_1200),
.Y(n_1331)
);

BUFx4f_ASAP7_75t_SL g1332 ( 
.A(n_1197),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1197),
.B(n_1200),
.Y(n_1333)
);

BUFx8_ASAP7_75t_L g1334 ( 
.A(n_1208),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_1211),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_SL g1336 ( 
.A1(n_1212),
.A2(n_1195),
.B1(n_1266),
.B2(n_1250),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1213),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1167),
.B(n_1175),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1163),
.A2(n_1202),
.B1(n_1188),
.B2(n_1203),
.Y(n_1339)
);

BUFx8_ASAP7_75t_SL g1340 ( 
.A(n_1179),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1175),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1146),
.B(n_1169),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1191),
.Y(n_1343)
);

OAI22xp5_ASAP7_75t_L g1344 ( 
.A1(n_1147),
.A2(n_1165),
.B1(n_1185),
.B2(n_1162),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1174),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1254),
.Y(n_1346)
);

INVx4_ASAP7_75t_L g1347 ( 
.A(n_1146),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1169),
.B(n_1249),
.Y(n_1348)
);

OAI22xp5_ASAP7_75t_L g1349 ( 
.A1(n_1150),
.A2(n_1236),
.B1(n_1267),
.B2(n_1249),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1204),
.B(n_1224),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1224),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1265),
.A2(n_1248),
.B1(n_1204),
.B2(n_1226),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1204),
.A2(n_581),
.B1(n_1242),
.B2(n_1227),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1154),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1157),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1227),
.A2(n_1242),
.B1(n_1271),
.B2(n_1139),
.Y(n_1356)
);

HB1xp67_ASAP7_75t_L g1357 ( 
.A(n_1148),
.Y(n_1357)
);

BUFx2_ASAP7_75t_L g1358 ( 
.A(n_1276),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1221),
.A2(n_812),
.B(n_1238),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1221),
.B(n_1238),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1221),
.A2(n_812),
.B1(n_1241),
.B2(n_1238),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1143),
.B(n_1148),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1154),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1154),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1154),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1367)
);

BUFx8_ASAP7_75t_SL g1368 ( 
.A(n_1246),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1221),
.A2(n_1139),
.B1(n_424),
.B2(n_978),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1154),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1221),
.B(n_1238),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_SL g1372 ( 
.A1(n_1221),
.A2(n_1139),
.B1(n_1241),
.B2(n_1238),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1157),
.Y(n_1373)
);

INVx6_ASAP7_75t_L g1374 ( 
.A(n_1164),
.Y(n_1374)
);

BUFx12f_ASAP7_75t_L g1375 ( 
.A(n_1176),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1221),
.A2(n_812),
.B1(n_1241),
.B2(n_1238),
.Y(n_1376)
);

BUFx10_ASAP7_75t_L g1377 ( 
.A(n_1176),
.Y(n_1377)
);

INVx11_ASAP7_75t_L g1378 ( 
.A(n_1276),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_1157),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1269),
.Y(n_1381)
);

CKINVDCx16_ASAP7_75t_R g1382 ( 
.A(n_1246),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1276),
.Y(n_1383)
);

BUFx2_ASAP7_75t_R g1384 ( 
.A(n_1176),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1154),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1154),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1190),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_L g1390 ( 
.A(n_1221),
.B(n_1238),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1221),
.A2(n_812),
.B1(n_1241),
.B2(n_1238),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1269),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1227),
.A2(n_581),
.B1(n_1271),
.B2(n_1242),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1227),
.A2(n_1242),
.B1(n_1271),
.B2(n_725),
.Y(n_1396)
);

NAND2xp33_ASAP7_75t_L g1397 ( 
.A(n_1303),
.B(n_1362),
.Y(n_1397)
);

INVx3_ASAP7_75t_L g1398 ( 
.A(n_1347),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1311),
.Y(n_1399)
);

OR2x6_ASAP7_75t_L g1400 ( 
.A(n_1301),
.B(n_1308),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1369),
.A2(n_1389),
.B1(n_1395),
.B2(n_1393),
.Y(n_1401)
);

AND2x6_ASAP7_75t_L g1402 ( 
.A(n_1304),
.B(n_1356),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1372),
.A2(n_1288),
.B1(n_1359),
.B2(n_1281),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1372),
.B(n_1360),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1311),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1341),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1326),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1360),
.B(n_1371),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1371),
.B(n_1390),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1390),
.B(n_1321),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1362),
.B(n_1376),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1338),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1338),
.Y(n_1413)
);

OR2x2_ASAP7_75t_L g1414 ( 
.A(n_1296),
.B(n_1376),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1351),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1392),
.B(n_1296),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1348),
.A2(n_1342),
.B(n_1352),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1392),
.B(n_1284),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1315),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1315),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1344),
.A2(n_1349),
.B(n_1326),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1345),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1346),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1337),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1286),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1287),
.B(n_1290),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1291),
.B(n_1293),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1323),
.A2(n_1342),
.B(n_1348),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1361),
.A2(n_1391),
.B1(n_1388),
.B2(n_1380),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1322),
.B(n_1297),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1323),
.A2(n_1309),
.B(n_1316),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1357),
.Y(n_1432)
);

BUFx4f_ASAP7_75t_SL g1433 ( 
.A(n_1283),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1396),
.A2(n_1307),
.B(n_1320),
.Y(n_1434)
);

NAND2x1_ASAP7_75t_L g1435 ( 
.A(n_1316),
.B(n_1343),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1367),
.A2(n_1306),
.B1(n_1295),
.B2(n_1353),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1309),
.A2(n_1325),
.B(n_1331),
.Y(n_1437)
);

OR2x2_ASAP7_75t_L g1438 ( 
.A(n_1363),
.B(n_1350),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1354),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1364),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1365),
.Y(n_1441)
);

O2A1O1Ixp33_ASAP7_75t_SL g1442 ( 
.A1(n_1292),
.A2(n_1394),
.B(n_1312),
.C(n_1355),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1366),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1370),
.B(n_1385),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1350),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1386),
.B(n_1282),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1297),
.B(n_1292),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1343),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1298),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1343),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1336),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1339),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1285),
.B2(n_1340),
.Y(n_1453)
);

OAI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1335),
.A2(n_1313),
.B1(n_1310),
.B2(n_1332),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1328),
.B(n_1333),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1330),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1313),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1300),
.A2(n_1334),
.B1(n_1314),
.B2(n_1319),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1327),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1387),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1313),
.B(n_1302),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1368),
.Y(n_1462)
);

INVx2_ASAP7_75t_SL g1463 ( 
.A(n_1302),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1302),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1381),
.B(n_1358),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_1418),
.Y(n_1466)
);

NAND4xp25_ASAP7_75t_L g1467 ( 
.A(n_1403),
.B(n_1381),
.C(n_1383),
.D(n_1299),
.Y(n_1467)
);

NOR2xp33_ASAP7_75t_L g1468 ( 
.A(n_1408),
.B(n_1382),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1433),
.B(n_1384),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1406),
.Y(n_1470)
);

OA21x2_ASAP7_75t_L g1471 ( 
.A1(n_1407),
.A2(n_1374),
.B(n_1294),
.Y(n_1471)
);

AOI22xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1411),
.A2(n_1317),
.B1(n_1324),
.B2(n_1289),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1416),
.B(n_1411),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1418),
.B(n_1373),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1404),
.B(n_1416),
.Y(n_1475)
);

BUFx2_ASAP7_75t_L g1476 ( 
.A(n_1399),
.Y(n_1476)
);

AOI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1449),
.A2(n_1310),
.B1(n_1305),
.B2(n_1379),
.C(n_1384),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1414),
.B(n_1377),
.Y(n_1478)
);

OR2x2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1378),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1397),
.A2(n_1377),
.B(n_1375),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1414),
.B(n_1447),
.Y(n_1481)
);

O2A1O1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1442),
.A2(n_1401),
.B(n_1434),
.C(n_1430),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1447),
.B(n_1446),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_SL g1484 ( 
.A1(n_1431),
.A2(n_1436),
.B(n_1452),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1446),
.B(n_1426),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1427),
.B(n_1444),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1444),
.B(n_1455),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1438),
.B(n_1412),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1455),
.B(n_1425),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1415),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1436),
.A2(n_1435),
.B(n_1429),
.C(n_1410),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1439),
.B(n_1440),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1440),
.B(n_1443),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1399),
.Y(n_1494)
);

A2O1A1Ixp33_ASAP7_75t_L g1495 ( 
.A1(n_1435),
.A2(n_1410),
.B(n_1437),
.C(n_1451),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1443),
.B(n_1413),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1419),
.B(n_1420),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1402),
.A2(n_1437),
.B(n_1407),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1409),
.B(n_1460),
.Y(n_1499)
);

INVxp67_ASAP7_75t_SL g1500 ( 
.A(n_1405),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1415),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1405),
.B(n_1428),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1453),
.A2(n_1432),
.B1(n_1458),
.B2(n_1456),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1428),
.B(n_1445),
.Y(n_1504)
);

OAI21xp5_ASAP7_75t_L g1505 ( 
.A1(n_1402),
.A2(n_1421),
.B(n_1448),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1434),
.A2(n_1402),
.B1(n_1456),
.B2(n_1454),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_SL g1507 ( 
.A1(n_1462),
.A2(n_1457),
.B(n_1463),
.C(n_1464),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1421),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1417),
.B(n_1423),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1400),
.B(n_1424),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1470),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1466),
.B(n_1417),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1470),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1508),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1481),
.B(n_1417),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1476),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1476),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1502),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1501),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1481),
.B(n_1422),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1473),
.B(n_1417),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.B(n_1398),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1494),
.B(n_1497),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1483),
.B(n_1398),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1471),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1506),
.A2(n_1402),
.B1(n_1450),
.B2(n_1400),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1494),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1502),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1486),
.B(n_1485),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1509),
.Y(n_1531)
);

NAND2x1_ASAP7_75t_L g1532 ( 
.A(n_1471),
.B(n_1450),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1509),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1491),
.A2(n_1461),
.B1(n_1457),
.B2(n_1459),
.Y(n_1534)
);

NAND2xp33_ASAP7_75t_R g1535 ( 
.A(n_1512),
.B(n_1471),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1516),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1514),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1522),
.B(n_1475),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1518),
.Y(n_1540)
);

AOI221xp5_ASAP7_75t_L g1541 ( 
.A1(n_1512),
.A2(n_1482),
.B1(n_1503),
.B2(n_1484),
.C(n_1495),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1515),
.B(n_1487),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1517),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

INVx1_ASAP7_75t_SL g1545 ( 
.A(n_1517),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1522),
.B(n_1500),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1528),
.Y(n_1547)
);

AOI22xp33_ASAP7_75t_L g1548 ( 
.A1(n_1527),
.A2(n_1506),
.B1(n_1498),
.B2(n_1467),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1518),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1515),
.B(n_1489),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1512),
.B(n_1489),
.Y(n_1551)
);

NAND3xp33_ASAP7_75t_L g1552 ( 
.A(n_1519),
.B(n_1467),
.C(n_1472),
.Y(n_1552)
);

INVxp67_ASAP7_75t_L g1553 ( 
.A(n_1528),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1529),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1520),
.Y(n_1555)
);

OAI222xp33_ASAP7_75t_L g1556 ( 
.A1(n_1534),
.A2(n_1472),
.B1(n_1504),
.B2(n_1510),
.C1(n_1474),
.C2(n_1478),
.Y(n_1556)
);

BUFx3_ASAP7_75t_L g1557 ( 
.A(n_1526),
.Y(n_1557)
);

NAND4xp25_ASAP7_75t_SL g1558 ( 
.A(n_1527),
.B(n_1477),
.C(n_1480),
.D(n_1478),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1531),
.B(n_1488),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1530),
.B(n_1471),
.Y(n_1560)
);

NAND4xp25_ASAP7_75t_L g1561 ( 
.A(n_1524),
.B(n_1468),
.C(n_1469),
.D(n_1499),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1531),
.A2(n_1505),
.B1(n_1496),
.B2(n_1493),
.C(n_1492),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1563)
);

OR2x6_ASAP7_75t_L g1564 ( 
.A(n_1532),
.B(n_1510),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1530),
.B(n_1474),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1540),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1545),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1544),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1544),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1560),
.B(n_1533),
.Y(n_1572)
);

OR2x2_ASAP7_75t_L g1573 ( 
.A(n_1539),
.B(n_1521),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1537),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1537),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1539),
.B(n_1524),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1539),
.B(n_1521),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1560),
.B(n_1523),
.Y(n_1579)
);

AND2x4_ASAP7_75t_SL g1580 ( 
.A(n_1563),
.B(n_1474),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1549),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1549),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1546),
.B(n_1553),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1557),
.Y(n_1584)
);

AND2x6_ASAP7_75t_SL g1585 ( 
.A(n_1563),
.B(n_1465),
.Y(n_1585)
);

OR2x6_ASAP7_75t_L g1586 ( 
.A(n_1564),
.B(n_1532),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1538),
.B(n_1542),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1555),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1511),
.Y(n_1589)
);

INVxp67_ASAP7_75t_L g1590 ( 
.A(n_1552),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1557),
.Y(n_1591)
);

AND2x4_ASAP7_75t_SL g1592 ( 
.A(n_1563),
.B(n_1525),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1511),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1590),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1574),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1574),
.Y(n_1598)
);

NAND2x2_ASAP7_75t_L g1599 ( 
.A(n_1591),
.B(n_1479),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1567),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1574),
.Y(n_1601)
);

NAND2x1_ASAP7_75t_L g1602 ( 
.A(n_1594),
.B(n_1543),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1567),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1590),
.B(n_1551),
.Y(n_1605)
);

INVx6_ASAP7_75t_L g1606 ( 
.A(n_1585),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1565),
.Y(n_1607)
);

NAND2x1p5_ASAP7_75t_L g1608 ( 
.A(n_1584),
.B(n_1532),
.Y(n_1608)
);

INVx4_ASAP7_75t_L g1609 ( 
.A(n_1585),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1568),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1587),
.B(n_1565),
.Y(n_1611)
);

NOR2xp33_ASAP7_75t_L g1612 ( 
.A(n_1580),
.B(n_1561),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1569),
.B(n_1551),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1568),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1587),
.B(n_1565),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1570),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1592),
.B(n_1550),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1569),
.B(n_1551),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1570),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1571),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1571),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1575),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1581),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1577),
.B(n_1554),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_L g1626 ( 
.A(n_1584),
.B(n_1558),
.C(n_1552),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1550),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1592),
.B(n_1550),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1581),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1582),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1582),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1588),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1580),
.B(n_1547),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1588),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1573),
.B(n_1559),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1575),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1596),
.B(n_1583),
.Y(n_1639)
);

OAI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1635),
.A2(n_1548),
.B1(n_1534),
.B2(n_1586),
.C1(n_1526),
.C2(n_1594),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1605),
.B(n_1578),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1598),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1609),
.B(n_1594),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_SL g1644 ( 
.A1(n_1626),
.A2(n_1625),
.B(n_1603),
.C(n_1610),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1604),
.B(n_1578),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1600),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1598),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1598),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1606),
.Y(n_1649)
);

INVxp67_ASAP7_75t_L g1650 ( 
.A(n_1612),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1600),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1603),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1604),
.B(n_1589),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1610),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_SL g1656 ( 
.A(n_1609),
.B(n_1594),
.Y(n_1656)
);

NOR3xp33_ASAP7_75t_L g1657 ( 
.A(n_1609),
.B(n_1558),
.C(n_1541),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1618),
.B(n_1594),
.Y(n_1658)
);

CKINVDCx16_ASAP7_75t_R g1659 ( 
.A(n_1630),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1637),
.B(n_1589),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1591),
.Y(n_1662)
);

HB1xp67_ASAP7_75t_L g1663 ( 
.A(n_1614),
.Y(n_1663)
);

INVx1_ASAP7_75t_SL g1664 ( 
.A(n_1606),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1637),
.B(n_1593),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1616),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1606),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1628),
.B(n_1591),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1628),
.B(n_1579),
.Y(n_1669)
);

INVx3_ASAP7_75t_L g1670 ( 
.A(n_1606),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1602),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1617),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1616),
.B(n_1593),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1627),
.B(n_1576),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1651),
.Y(n_1675)
);

AOI31xp33_ASAP7_75t_L g1676 ( 
.A1(n_1650),
.A2(n_1608),
.A3(n_1630),
.B(n_1634),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1644),
.B(n_1561),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1653),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1613),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1657),
.B(n_1607),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1657),
.A2(n_1644),
.B1(n_1541),
.B2(n_1649),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1649),
.Y(n_1682)
);

XNOR2x1_ASAP7_75t_L g1683 ( 
.A(n_1664),
.B(n_1608),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1639),
.B(n_1607),
.Y(n_1684)
);

OAI32xp33_ASAP7_75t_L g1685 ( 
.A1(n_1659),
.A2(n_1599),
.A3(n_1667),
.B1(n_1664),
.B2(n_1639),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1663),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1640),
.A2(n_1619),
.B(n_1602),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1666),
.Y(n_1688)
);

CKINVDCx14_ASAP7_75t_R g1689 ( 
.A(n_1651),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1646),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1646),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1645),
.B(n_1611),
.Y(n_1692)
);

INVx2_ASAP7_75t_SL g1693 ( 
.A(n_1643),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1652),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1652),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1640),
.A2(n_1656),
.B(n_1667),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1655),
.Y(n_1697)
);

AOI211x1_ASAP7_75t_L g1698 ( 
.A1(n_1662),
.A2(n_1556),
.B(n_1634),
.C(n_1611),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1659),
.B(n_1615),
.Y(n_1699)
);

OAI321xp33_ASAP7_75t_L g1700 ( 
.A1(n_1650),
.A2(n_1608),
.A3(n_1548),
.B1(n_1586),
.B2(n_1638),
.C(n_1617),
.Y(n_1700)
);

AOI22xp5_ASAP7_75t_L g1701 ( 
.A1(n_1677),
.A2(n_1535),
.B1(n_1670),
.B2(n_1599),
.Y(n_1701)
);

INVx1_ASAP7_75t_SL g1702 ( 
.A(n_1682),
.Y(n_1702)
);

XNOR2x1_ASAP7_75t_SL g1703 ( 
.A(n_1693),
.B(n_1670),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1699),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1677),
.A2(n_1535),
.B1(n_1670),
.B2(n_1599),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1693),
.Y(n_1706)
);

AOI22xp33_ASAP7_75t_L g1707 ( 
.A1(n_1681),
.A2(n_1526),
.B1(n_1670),
.B2(n_1672),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1680),
.B(n_1641),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1690),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1681),
.B(n_1662),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1689),
.B(n_1662),
.Y(n_1711)
);

NOR2xp33_ASAP7_75t_L g1712 ( 
.A(n_1689),
.B(n_1643),
.Y(n_1712)
);

NOR2xp33_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1643),
.Y(n_1713)
);

INVxp67_ASAP7_75t_SL g1714 ( 
.A(n_1683),
.Y(n_1714)
);

OAI21xp5_ASAP7_75t_SL g1715 ( 
.A1(n_1676),
.A2(n_1643),
.B(n_1668),
.Y(n_1715)
);

HB1xp67_ASAP7_75t_L g1716 ( 
.A(n_1699),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1678),
.B(n_1668),
.Y(n_1717)
);

AOI211xp5_ASAP7_75t_L g1718 ( 
.A1(n_1685),
.A2(n_1643),
.B(n_1655),
.C(n_1660),
.Y(n_1718)
);

OAI21xp33_ASAP7_75t_L g1719 ( 
.A1(n_1687),
.A2(n_1668),
.B(n_1641),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1716),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1704),
.B(n_1686),
.Y(n_1722)
);

NAND2xp33_ASAP7_75t_SL g1723 ( 
.A(n_1710),
.B(n_1688),
.Y(n_1723)
);

HB1xp67_ASAP7_75t_L g1724 ( 
.A(n_1703),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1702),
.B(n_1692),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1706),
.Y(n_1726)
);

XOR2xp5_ASAP7_75t_L g1727 ( 
.A(n_1708),
.B(n_1683),
.Y(n_1727)
);

OAI22xp5_ASAP7_75t_L g1728 ( 
.A1(n_1718),
.A2(n_1698),
.B1(n_1705),
.B2(n_1701),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1706),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1658),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1717),
.Y(n_1731)
);

XNOR2xp5_ASAP7_75t_L g1732 ( 
.A(n_1714),
.B(n_1696),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1732),
.A2(n_1719),
.B1(n_1707),
.B2(n_1712),
.Y(n_1733)
);

NOR2xp33_ASAP7_75t_L g1734 ( 
.A(n_1724),
.B(n_1711),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1725),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1730),
.B(n_1700),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1724),
.B(n_1715),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1723),
.B(n_1671),
.Y(n_1738)
);

NAND3x1_ASAP7_75t_L g1739 ( 
.A(n_1722),
.B(n_1713),
.C(n_1709),
.Y(n_1739)
);

NOR3xp33_ASAP7_75t_L g1740 ( 
.A(n_1723),
.B(n_1729),
.C(n_1726),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1721),
.Y(n_1741)
);

NOR2x1p5_ASAP7_75t_L g1742 ( 
.A(n_1731),
.B(n_1720),
.Y(n_1742)
);

AOI211xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1728),
.A2(n_1684),
.B(n_1695),
.C(n_1694),
.Y(n_1743)
);

NAND2xp33_ASAP7_75t_SL g1744 ( 
.A(n_1735),
.B(n_1671),
.Y(n_1744)
);

AOI221xp5_ASAP7_75t_L g1745 ( 
.A1(n_1736),
.A2(n_1727),
.B1(n_1697),
.B2(n_1672),
.C(n_1642),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1740),
.A2(n_1642),
.B1(n_1672),
.B2(n_1647),
.C(n_1648),
.Y(n_1746)
);

OAI222xp33_ASAP7_75t_L g1747 ( 
.A1(n_1733),
.A2(n_1679),
.B1(n_1642),
.B2(n_1647),
.C1(n_1648),
.C2(n_1671),
.Y(n_1747)
);

AOI221xp5_ASAP7_75t_L g1748 ( 
.A1(n_1734),
.A2(n_1647),
.B1(n_1648),
.B2(n_1660),
.C(n_1673),
.Y(n_1748)
);

NAND4xp75_ASAP7_75t_L g1749 ( 
.A(n_1737),
.B(n_1658),
.C(n_1665),
.D(n_1669),
.Y(n_1749)
);

AOI222xp33_ASAP7_75t_L g1750 ( 
.A1(n_1745),
.A2(n_1738),
.B1(n_1741),
.B2(n_1742),
.C1(n_1743),
.C2(n_1739),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1747),
.A2(n_1665),
.B(n_1658),
.C(n_1661),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1746),
.A2(n_1673),
.B1(n_1661),
.B2(n_1654),
.C(n_1617),
.Y(n_1752)
);

OAI211xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1748),
.A2(n_1654),
.B(n_1674),
.C(n_1631),
.Y(n_1753)
);

OAI211xp5_ASAP7_75t_SL g1754 ( 
.A1(n_1749),
.A2(n_1674),
.B(n_1631),
.C(n_1629),
.Y(n_1754)
);

OAI321xp33_ASAP7_75t_L g1755 ( 
.A1(n_1744),
.A2(n_1586),
.A3(n_1669),
.B1(n_1638),
.B2(n_1597),
.C(n_1601),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1750),
.A2(n_1669),
.B(n_1636),
.C(n_1633),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1751),
.B(n_1620),
.Y(n_1757)
);

NOR2x1_ASAP7_75t_L g1758 ( 
.A(n_1754),
.B(n_1620),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1753),
.B(n_1621),
.Y(n_1759)
);

NOR2x1_ASAP7_75t_L g1760 ( 
.A(n_1755),
.B(n_1621),
.Y(n_1760)
);

AOI221xp5_ASAP7_75t_L g1761 ( 
.A1(n_1756),
.A2(n_1752),
.B1(n_1638),
.B2(n_1597),
.C(n_1601),
.Y(n_1761)
);

OAI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1760),
.A2(n_1623),
.B1(n_1633),
.B2(n_1632),
.C(n_1629),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1757),
.B(n_1622),
.Y(n_1763)
);

OAI22x1_ASAP7_75t_L g1764 ( 
.A1(n_1763),
.A2(n_1758),
.B1(n_1759),
.B2(n_1465),
.Y(n_1764)
);

AOI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1764),
.A2(n_1762),
.B1(n_1761),
.B2(n_1623),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1765),
.Y(n_1766)
);

INVx4_ASAP7_75t_L g1767 ( 
.A(n_1765),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1767),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1767),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1769),
.A2(n_1766),
.B1(n_1636),
.B2(n_1632),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_L g1771 ( 
.A1(n_1768),
.A2(n_1624),
.B(n_1622),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1771),
.B(n_1624),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1772),
.A2(n_1770),
.B1(n_1566),
.B2(n_1572),
.Y(n_1773)
);

NAND2xp33_ASAP7_75t_L g1774 ( 
.A(n_1773),
.B(n_1615),
.Y(n_1774)
);

OAI221xp5_ASAP7_75t_R g1775 ( 
.A1(n_1774),
.A2(n_1545),
.B1(n_1580),
.B2(n_1595),
.C(n_1536),
.Y(n_1775)
);

AOI211xp5_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1457),
.B(n_1479),
.C(n_1507),
.Y(n_1776)
);


endmodule