module fake_netlist_6_2358_n_925 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_925);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_925;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_832;
wire n_280;
wire n_287;
wire n_685;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_758;
wire n_720;
wire n_842;
wire n_525;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_850;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_7),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_39),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_97),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_55),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_18),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_43),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_127),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_77),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_117),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_82),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_37),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_11),
.Y(n_201)
);

BUFx8_ASAP7_75t_SL g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_94),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_169),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_108),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_71),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_1),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_112),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_45),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_46),
.Y(n_215)
);

BUFx8_ASAP7_75t_SL g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_22),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_44),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_7),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_19),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_17),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_73),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_96),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_123),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_1),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_90),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_163),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_9),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_158),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_22),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_143),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_48),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_165),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_56),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_162),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_101),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_83),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_0),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_28),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_157),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_104),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_87),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_161),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_144),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_67),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_125),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_17),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_168),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_202),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_199),
.B(n_0),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_202),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_251),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_230),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_191),
.B(n_185),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_201),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_188),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_195),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_187),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_215),
.B(n_2),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_216),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_189),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_190),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_189),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_250),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_193),
.Y(n_278)
);

BUFx6f_ASAP7_75t_SL g279 ( 
.A(n_250),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_184),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_217),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_218),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_194),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_221),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_199),
.B(n_3),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_196),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_210),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_226),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_229),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_208),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_197),
.Y(n_298)
);

INVxp33_ASAP7_75t_SL g299 ( 
.A(n_231),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_236),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_256),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_3),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_254),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_192),
.B(n_4),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_198),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_214),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_273),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_306),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_276),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_259),
.B(n_243),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_280),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_270),
.B(n_192),
.Y(n_319)
);

BUFx8_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_277),
.B(n_204),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_264),
.Y(n_322)
);

NAND2x1_ASAP7_75t_L g323 ( 
.A(n_271),
.B(n_214),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_271),
.B(n_214),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_274),
.B(n_200),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_200),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_263),
.B(n_248),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g330 ( 
.A1(n_261),
.A2(n_222),
.B(n_205),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_281),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_299),
.B(n_203),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_269),
.B(n_205),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_299),
.B(n_206),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_268),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_300),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_234),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_260),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_286),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_290),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_281),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_267),
.B(n_245),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_245),
.Y(n_354)
);

BUFx8_ASAP7_75t_L g355 ( 
.A(n_279),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_275),
.Y(n_356)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_289),
.Y(n_357)
);

OAI21x1_ASAP7_75t_L g358 ( 
.A1(n_279),
.A2(n_247),
.B(n_244),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_289),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_307),
.Y(n_360)
);

OR2x6_ASAP7_75t_L g361 ( 
.A(n_359),
.B(n_357),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_335),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_337),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_265),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_252),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_329),
.B(n_293),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_339),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_323),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_329),
.B(n_257),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_309),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_329),
.B(n_294),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_312),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_354),
.B(n_294),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_344),
.Y(n_377)
);

AND2x4_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_207),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_347),
.B(n_209),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_325),
.B(n_301),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_340),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_301),
.B1(n_238),
.B2(n_237),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_326),
.B(n_211),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_262),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_354),
.B(n_212),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVx4_ASAP7_75t_L g391 ( 
.A(n_336),
.Y(n_391)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_336),
.Y(n_392)
);

AND2x6_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_27),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

AND2x4_ASAP7_75t_L g395 ( 
.A(n_344),
.B(n_213),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_311),
.B(n_262),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_340),
.Y(n_397)
);

OR2x2_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_258),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_223),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_342),
.B(n_224),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_333),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_345),
.B(n_225),
.Y(n_405)
);

AND2x4_ASAP7_75t_SL g406 ( 
.A(n_357),
.B(n_272),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_343),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_324),
.B(n_227),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_357),
.B(n_228),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_341),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_356),
.B(n_282),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_232),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_352),
.B(n_235),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_320),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_341),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_313),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_315),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_314),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_314),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_346),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_322),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_327),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_327),
.B(n_239),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_331),
.B(n_241),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_317),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_317),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_338),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_331),
.B(n_242),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_394),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_417),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_417),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_358),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_420),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_420),
.Y(n_439)
);

NAND2x1p5_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_349),
.Y(n_440)
);

AO22x2_ASAP7_75t_L g441 ( 
.A1(n_375),
.A2(n_321),
.B1(n_328),
.B2(n_332),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_419),
.Y(n_442)
);

NAND2x1p5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_349),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_422),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

NAND2x1p5_ASAP7_75t_L g446 ( 
.A(n_403),
.B(n_350),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_368),
.Y(n_448)
);

OAI221xp5_ASAP7_75t_L g449 ( 
.A1(n_385),
.A2(n_318),
.B1(n_334),
.B2(n_249),
.C(n_255),
.Y(n_449)
);

AO22x2_ASAP7_75t_L g450 ( 
.A1(n_375),
.A2(n_316),
.B1(n_243),
.B2(n_6),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_381),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_383),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_397),
.B(n_358),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_416),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_330),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_425),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_318),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_384),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_367),
.A2(n_351),
.B1(n_246),
.B2(n_330),
.Y(n_459)
);

NAND2x1p5_ASAP7_75t_L g460 ( 
.A(n_369),
.B(n_320),
.Y(n_460)
);

NAND2x1p5_ASAP7_75t_L g461 ( 
.A(n_369),
.B(n_320),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_367),
.A2(n_373),
.B1(n_382),
.B2(n_380),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_362),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_364),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_401),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_401),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_399),
.B(n_316),
.Y(n_468)
);

AO22x2_ASAP7_75t_L g469 ( 
.A1(n_418),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_401),
.B(n_355),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_421),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_421),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_428),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_384),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_390),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_429),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_429),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_399),
.B(n_355),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_373),
.B(n_365),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_396),
.Y(n_482)
);

NAND2x1_ASAP7_75t_L g483 ( 
.A(n_393),
.B(n_29),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_418),
.A2(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_361),
.A2(n_369),
.B1(n_400),
.B2(n_386),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_411),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_411),
.Y(n_489)
);

AO22x2_ASAP7_75t_L g490 ( 
.A1(n_388),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_388),
.B(n_355),
.Y(n_491)
);

OAI221xp5_ASAP7_75t_L g492 ( 
.A1(n_389),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_492)
);

OAI221xp5_ASAP7_75t_L g493 ( 
.A1(n_389),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.C(n_15),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_387),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_378),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_387),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_378),
.B(n_30),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_372),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_360),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_415),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_360),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_363),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_415),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_409),
.A2(n_98),
.B1(n_182),
.B2(n_181),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_363),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_370),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_370),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_374),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_374),
.Y(n_510)
);

AO22x2_ASAP7_75t_L g511 ( 
.A1(n_427),
.A2(n_432),
.B1(n_398),
.B2(n_412),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_372),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_423),
.B(n_16),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_372),
.Y(n_514)
);

NAND2xp33_ASAP7_75t_SL g515 ( 
.A(n_480),
.B(n_409),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_463),
.B(n_369),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_SL g517 ( 
.A(n_470),
.B(n_395),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_505),
.B(n_366),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_495),
.B(n_391),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_444),
.B(n_361),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_481),
.B(n_391),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_442),
.B(n_414),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_497),
.B(n_426),
.Y(n_523)
);

NAND2xp33_ASAP7_75t_SL g524 ( 
.A(n_491),
.B(n_395),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_497),
.B(n_405),
.Y(n_525)
);

NAND2xp33_ASAP7_75t_SL g526 ( 
.A(n_513),
.B(n_395),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_447),
.B(n_459),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_484),
.B(n_405),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_482),
.B(n_378),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_445),
.B(n_379),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_464),
.B(n_379),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_501),
.B(n_379),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_448),
.B(n_407),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_468),
.B(n_361),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_465),
.B(n_443),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_504),
.B(n_483),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_451),
.B(n_407),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_446),
.B(n_407),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_486),
.B(n_407),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_452),
.B(n_408),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_457),
.B(n_454),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_456),
.B(n_413),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_462),
.B(n_361),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_457),
.B(n_406),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_479),
.B(n_487),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_489),
.B(n_406),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_440),
.B(n_437),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_437),
.B(n_392),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_433),
.B(n_392),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_433),
.B(n_392),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_434),
.B(n_371),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_434),
.B(n_392),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_435),
.B(n_392),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_466),
.B(n_393),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_435),
.B(n_410),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_436),
.B(n_410),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_436),
.B(n_410),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_511),
.B(n_366),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_438),
.B(n_410),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_438),
.B(n_410),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_467),
.B(n_393),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_494),
.B(n_393),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_439),
.B(n_371),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_439),
.B(n_376),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_471),
.B(n_376),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_472),
.B(n_376),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_473),
.B(n_476),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_477),
.B(n_478),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_460),
.B(n_393),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_461),
.B(n_393),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_453),
.B(n_371),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_453),
.B(n_371),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_509),
.B(n_371),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_496),
.B(n_371),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_SL g575 ( 
.A(n_538),
.B(n_492),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_534),
.A2(n_441),
.B1(n_511),
.B2(n_449),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_516),
.A2(n_455),
.B(n_518),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_533),
.Y(n_578)
);

OAI21x1_ASAP7_75t_L g579 ( 
.A1(n_551),
.A2(n_512),
.B(n_510),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_537),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_561),
.A2(n_498),
.B(n_512),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_522),
.B(n_509),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_564),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_530),
.B(n_441),
.Y(n_584)
);

AO31x2_ASAP7_75t_L g585 ( 
.A1(n_563),
.A2(n_510),
.A3(n_502),
.B(n_508),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_523),
.B(n_518),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_525),
.A2(n_490),
.B1(n_534),
.B2(n_493),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_558),
.Y(n_589)
);

A2O1A1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_526),
.A2(n_488),
.B(n_474),
.C(n_458),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_567),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_543),
.B(n_500),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_R g593 ( 
.A(n_520),
.B(n_554),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_573),
.A2(n_475),
.B(n_499),
.Y(n_594)
);

OAI21xp33_ASAP7_75t_SL g595 ( 
.A1(n_531),
.A2(n_507),
.B(n_506),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_554),
.A2(n_490),
.B1(n_450),
.B2(n_485),
.Y(n_597)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_562),
.A2(n_514),
.B(n_503),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_515),
.Y(n_599)
);

AOI211x1_ASAP7_75t_L g600 ( 
.A1(n_541),
.A2(n_450),
.B(n_485),
.C(n_469),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_571),
.A2(n_95),
.B(n_183),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_520),
.B(n_469),
.Y(n_602)
);

A2O1A1Ixp33_ASAP7_75t_L g603 ( 
.A1(n_540),
.A2(n_542),
.B(n_524),
.C(n_527),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_565),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_521),
.B(n_31),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_528),
.B(n_16),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_SL g607 ( 
.A1(n_539),
.A2(n_18),
.B(n_19),
.Y(n_607)
);

AO22x2_ASAP7_75t_L g608 ( 
.A1(n_535),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_566),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_532),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_544),
.B(n_20),
.Y(n_611)
);

OAI21x1_ASAP7_75t_L g612 ( 
.A1(n_572),
.A2(n_100),
.B(n_179),
.Y(n_612)
);

A2O1A1Ixp33_ASAP7_75t_L g613 ( 
.A1(n_517),
.A2(n_21),
.B(n_23),
.C(n_24),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_555),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_547),
.B(n_25),
.Y(n_615)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_546),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

O2A1O1Ixp5_ASAP7_75t_L g618 ( 
.A1(n_569),
.A2(n_106),
.B(n_177),
.C(n_32),
.Y(n_618)
);

NOR2xp67_ASAP7_75t_SL g619 ( 
.A(n_570),
.B(n_25),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_548),
.B(n_26),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_519),
.B(n_26),
.Y(n_621)
);

BUFx12f_ASAP7_75t_L g622 ( 
.A(n_536),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_545),
.Y(n_623)
);

OAI21x1_ASAP7_75t_L g624 ( 
.A1(n_574),
.A2(n_33),
.B(n_34),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_549),
.B(n_35),
.Y(n_625)
);

AO21x2_ASAP7_75t_L g626 ( 
.A1(n_577),
.A2(n_560),
.B(n_559),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_591),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_589),
.B(n_550),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_584),
.A2(n_553),
.B(n_552),
.C(n_557),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_577),
.A2(n_36),
.B(n_38),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_599),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_633)
);

NAND2x1p5_ASAP7_75t_L g634 ( 
.A(n_623),
.B(n_47),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_589),
.B(n_49),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

OAI21x1_ASAP7_75t_L g637 ( 
.A1(n_594),
.A2(n_50),
.B(n_51),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_609),
.Y(n_638)
);

NAND2x1p5_ASAP7_75t_L g639 ( 
.A(n_623),
.B(n_52),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_592),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_576),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_604),
.Y(n_642)
);

AO221x2_ASAP7_75t_L g643 ( 
.A1(n_597),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.C(n_61),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_585),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_579),
.A2(n_62),
.B(n_63),
.Y(n_645)
);

OR2x6_ASAP7_75t_L g646 ( 
.A(n_622),
.B(n_65),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_583),
.Y(n_647)
);

AND2x4_ASAP7_75t_L g648 ( 
.A(n_616),
.B(n_66),
.Y(n_648)
);

AO21x2_ASAP7_75t_L g649 ( 
.A1(n_603),
.A2(n_68),
.B(n_69),
.Y(n_649)
);

OAI22xp5_ASAP7_75t_L g650 ( 
.A1(n_582),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_620),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_582),
.B(n_78),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_578),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_580),
.B(n_80),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_610),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_617),
.Y(n_656)
);

OA21x2_ASAP7_75t_L g657 ( 
.A1(n_587),
.A2(n_81),
.B(n_84),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_615),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_614),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_593),
.Y(n_660)
);

AOI21x1_ASAP7_75t_L g661 ( 
.A1(n_605),
.A2(n_85),
.B(n_86),
.Y(n_661)
);

BUFx8_ASAP7_75t_L g662 ( 
.A(n_608),
.Y(n_662)
);

BUFx12f_ASAP7_75t_L g663 ( 
.A(n_608),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_611),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_606),
.B(n_92),
.Y(n_665)
);

A2O1A1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_588),
.A2(n_99),
.B(n_103),
.C(n_109),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

OR2x6_ASAP7_75t_L g668 ( 
.A(n_600),
.B(n_110),
.Y(n_668)
);

BUFx12f_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_581),
.A2(n_111),
.B(n_114),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_597),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_602),
.A2(n_115),
.B1(n_116),
.B2(n_118),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_653),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_627),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_653),
.Y(n_676)
);

HB1xp67_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_640),
.B(n_613),
.Y(n_678)
);

INVxp67_ASAP7_75t_L g679 ( 
.A(n_651),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_670),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_644),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_668),
.B(n_575),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_659),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_658),
.B(n_621),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g685 ( 
.A1(n_660),
.A2(n_625),
.B1(n_590),
.B2(n_598),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_659),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_648),
.B(n_612),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_655),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_668),
.B(n_607),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_629),
.B(n_619),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_668),
.B(n_643),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_648),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_651),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_636),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_638),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_656),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_637),
.A2(n_624),
.B(n_618),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_642),
.B(n_119),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_630),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_667),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_663),
.A2(n_595),
.B1(n_121),
.B2(n_124),
.Y(n_703)
);

CKINVDCx11_ASAP7_75t_R g704 ( 
.A(n_646),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_649),
.Y(n_705)
);

OA21x2_ASAP7_75t_L g706 ( 
.A1(n_666),
.A2(n_120),
.B(n_126),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_635),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_657),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_657),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_626),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_657),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_645),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_634),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_635),
.Y(n_714)
);

HB1xp67_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

BUFx2_ASAP7_75t_SL g716 ( 
.A(n_671),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_634),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_654),
.Y(n_718)
);

AOI21x1_ASAP7_75t_L g719 ( 
.A1(n_661),
.A2(n_128),
.B(n_131),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_652),
.A2(n_132),
.B(n_133),
.Y(n_720)
);

BUFx6f_ASAP7_75t_L g721 ( 
.A(n_639),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_626),
.Y(n_722)
);

OR2x6_ASAP7_75t_L g723 ( 
.A(n_663),
.B(n_669),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_669),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_643),
.B(n_135),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_707),
.B(n_662),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_677),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_R g728 ( 
.A(n_704),
.B(n_692),
.Y(n_728)
);

CKINVDCx6p67_ASAP7_75t_R g729 ( 
.A(n_688),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_700),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_R g731 ( 
.A(n_692),
.B(n_671),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_674),
.Y(n_732)
);

XNOR2xp5_ASAP7_75t_L g733 ( 
.A(n_716),
.B(n_646),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_R g734 ( 
.A(n_682),
.B(n_646),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_R g735 ( 
.A(n_692),
.B(n_721),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_714),
.B(n_643),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_R g737 ( 
.A(n_692),
.B(n_662),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_692),
.B(n_672),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_R g739 ( 
.A(n_682),
.B(n_632),
.Y(n_739)
);

INVxp67_ASAP7_75t_L g740 ( 
.A(n_716),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_SL g741 ( 
.A(n_725),
.B(n_641),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_674),
.B(n_666),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_R g743 ( 
.A(n_721),
.B(n_136),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_698),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_718),
.B(n_672),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_721),
.B(n_137),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_725),
.B(n_650),
.Y(n_747)
);

OR2x2_ASAP7_75t_L g748 ( 
.A(n_715),
.B(n_696),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_683),
.Y(n_749)
);

BUFx10_ASAP7_75t_L g750 ( 
.A(n_698),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_679),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_693),
.B(n_639),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_R g753 ( 
.A(n_706),
.B(n_138),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_717),
.B(n_633),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_R g755 ( 
.A(n_721),
.B(n_140),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_683),
.Y(n_756)
);

INVx8_ASAP7_75t_L g757 ( 
.A(n_698),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_694),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_R g759 ( 
.A(n_721),
.B(n_142),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_R g760 ( 
.A(n_706),
.B(n_145),
.Y(n_760)
);

XOR2xp5_ASAP7_75t_L g761 ( 
.A(n_687),
.B(n_664),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_696),
.B(n_146),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_678),
.B(n_631),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_686),
.Y(n_764)
);

CKINVDCx12_ASAP7_75t_R g765 ( 
.A(n_723),
.Y(n_765)
);

XNOR2xp5_ASAP7_75t_L g766 ( 
.A(n_724),
.B(n_147),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_678),
.B(n_631),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_676),
.B(n_149),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_732),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_749),
.Y(n_770)
);

NOR2x1_ASAP7_75t_L g771 ( 
.A(n_745),
.B(n_726),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_756),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_758),
.B(n_713),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_748),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_767),
.B(n_722),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_764),
.Y(n_776)
);

NOR2x1_ASAP7_75t_L g777 ( 
.A(n_726),
.B(n_713),
.Y(n_777)
);

NOR2xp67_ASAP7_75t_SL g778 ( 
.A(n_738),
.B(n_706),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_736),
.B(n_722),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_SL g780 ( 
.A1(n_766),
.A2(n_691),
.B(n_703),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_727),
.B(n_695),
.Y(n_781)
);

HB1xp67_ASAP7_75t_L g782 ( 
.A(n_730),
.Y(n_782)
);

BUFx2_ASAP7_75t_L g783 ( 
.A(n_735),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_763),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_741),
.A2(n_691),
.B1(n_723),
.B2(n_689),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_763),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_751),
.B(n_699),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_740),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_742),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_742),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_752),
.B(n_710),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_731),
.B(n_710),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_737),
.B(n_673),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_762),
.B(n_673),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_747),
.B(n_708),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_765),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_768),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_761),
.B(n_684),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_744),
.B(n_675),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_769),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_770),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_780),
.A2(n_723),
.B1(n_739),
.B2(n_760),
.Y(n_802)
);

BUFx2_ASAP7_75t_L g803 ( 
.A(n_795),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_SL g804 ( 
.A(n_798),
.B(n_759),
.C(n_755),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_779),
.B(n_709),
.Y(n_805)
);

AND2x2_ASAP7_75t_L g806 ( 
.A(n_779),
.B(n_709),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_783),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_770),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_769),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_772),
.Y(n_810)
);

OAI211xp5_ASAP7_75t_L g811 ( 
.A1(n_771),
.A2(n_746),
.B(n_743),
.C(n_724),
.Y(n_811)
);

AND2x4_ASAP7_75t_L g812 ( 
.A(n_791),
.B(n_711),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_784),
.B(n_708),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_775),
.B(n_711),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_775),
.B(n_705),
.Y(n_815)
);

OA21x2_ASAP7_75t_L g816 ( 
.A1(n_795),
.A2(n_705),
.B(n_701),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_784),
.B(n_701),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_772),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_818),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_818),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_802),
.B(n_786),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_800),
.B(n_774),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_808),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_809),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_807),
.B(n_791),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_809),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_803),
.B(n_790),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_810),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_810),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_801),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_808),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_803),
.B(n_782),
.Y(n_832)
);

OAI221xp5_ASAP7_75t_L g833 ( 
.A1(n_821),
.A2(n_811),
.B1(n_796),
.B2(n_785),
.C(n_734),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_832),
.B(n_800),
.Y(n_834)
);

OAI221xp5_ASAP7_75t_L g835 ( 
.A1(n_821),
.A2(n_811),
.B1(n_796),
.B2(n_733),
.C(n_804),
.Y(n_835)
);

NOR2x1_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_807),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_825),
.A2(n_802),
.B1(n_804),
.B2(n_723),
.Y(n_837)
);

OAI22xp33_ASAP7_75t_L g838 ( 
.A1(n_827),
.A2(n_753),
.B1(n_807),
.B2(n_783),
.Y(n_838)
);

AO221x2_ASAP7_75t_L g839 ( 
.A1(n_824),
.A2(n_787),
.B1(n_781),
.B2(n_789),
.C(n_797),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_834),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_839),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_836),
.B(n_837),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_833),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_835),
.B(n_729),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_839),
.B(n_826),
.Y(n_846)
);

NOR2x1_ASAP7_75t_L g847 ( 
.A(n_836),
.B(n_819),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_847),
.B(n_820),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_843),
.B(n_822),
.Y(n_849)
);

XNOR2xp5_ASAP7_75t_L g850 ( 
.A(n_844),
.B(n_777),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_840),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_848),
.Y(n_853)
);

NOR2xp33_ASAP7_75t_L g854 ( 
.A(n_849),
.B(n_845),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_850),
.B(n_842),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_852),
.B(n_841),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_853),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_856),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_855),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_854),
.Y(n_860)
);

NOR3x1_ASAP7_75t_L g861 ( 
.A(n_859),
.B(n_851),
.C(n_846),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_860),
.A2(n_848),
.B(n_720),
.Y(n_862)
);

AOI211xp5_ASAP7_75t_L g863 ( 
.A1(n_858),
.A2(n_728),
.B(n_778),
.C(n_788),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_857),
.Y(n_864)
);

AOI221xp5_ASAP7_75t_L g865 ( 
.A1(n_857),
.A2(n_778),
.B1(n_829),
.B2(n_828),
.C(n_789),
.Y(n_865)
);

NOR3xp33_ASAP7_75t_L g866 ( 
.A(n_859),
.B(n_690),
.C(n_685),
.Y(n_866)
);

NAND4xp25_ASAP7_75t_SL g867 ( 
.A(n_860),
.B(n_793),
.C(n_792),
.D(n_823),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_864),
.A2(n_830),
.B1(n_689),
.B2(n_823),
.C(n_831),
.Y(n_868)
);

AOI211xp5_ASAP7_75t_L g869 ( 
.A1(n_862),
.A2(n_773),
.B(n_793),
.C(n_754),
.Y(n_869)
);

AOI221x1_ASAP7_75t_L g870 ( 
.A1(n_866),
.A2(n_831),
.B1(n_808),
.B2(n_801),
.C(n_776),
.Y(n_870)
);

OAI221xp5_ASAP7_75t_L g871 ( 
.A1(n_863),
.A2(n_706),
.B1(n_797),
.B2(n_713),
.C(n_717),
.Y(n_871)
);

AOI211xp5_ASAP7_75t_L g872 ( 
.A1(n_867),
.A2(n_754),
.B(n_687),
.C(n_792),
.Y(n_872)
);

AOI221x1_ASAP7_75t_L g873 ( 
.A1(n_861),
.A2(n_808),
.B1(n_801),
.B2(n_776),
.C(n_712),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_865),
.A2(n_757),
.B1(n_812),
.B2(n_815),
.Y(n_874)
);

NOR2x1_ASAP7_75t_L g875 ( 
.A(n_871),
.B(n_816),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_874),
.A2(n_790),
.B1(n_812),
.B2(n_813),
.Y(n_876)
);

NOR2xp67_ASAP7_75t_L g877 ( 
.A(n_873),
.B(n_869),
.Y(n_877)
);

NOR3x2_ASAP7_75t_L g878 ( 
.A(n_870),
.B(n_813),
.C(n_152),
.Y(n_878)
);

NOR2x1_ASAP7_75t_L g879 ( 
.A(n_872),
.B(n_816),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_868),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_871),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_872),
.B(n_814),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_873),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_R g884 ( 
.A(n_881),
.B(n_150),
.Y(n_884)
);

NAND2xp33_ASAP7_75t_SL g885 ( 
.A(n_883),
.B(n_799),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_877),
.B(n_812),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_879),
.B(n_812),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_880),
.B(n_814),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_875),
.B(n_817),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_SL g890 ( 
.A(n_882),
.B(n_799),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_876),
.B(n_878),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_877),
.B(n_817),
.Y(n_892)
);

NAND2x1_ASAP7_75t_SL g893 ( 
.A(n_883),
.B(n_816),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_SL g894 ( 
.A(n_883),
.B(n_806),
.Y(n_894)
);

AOI211xp5_ASAP7_75t_L g895 ( 
.A1(n_891),
.A2(n_687),
.B(n_794),
.C(n_815),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_890),
.A2(n_757),
.B1(n_806),
.B2(n_805),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_885),
.Y(n_897)
);

OR2x2_ASAP7_75t_L g898 ( 
.A(n_888),
.B(n_805),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_893),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_884),
.B(n_816),
.Y(n_900)
);

AOI221xp5_ASAP7_75t_L g901 ( 
.A1(n_894),
.A2(n_757),
.B1(n_794),
.B2(n_712),
.C(n_686),
.Y(n_901)
);

XNOR2x1_ASAP7_75t_L g902 ( 
.A(n_886),
.B(n_153),
.Y(n_902)
);

NAND4xp25_ASAP7_75t_L g903 ( 
.A(n_897),
.B(n_892),
.C(n_889),
.D(n_887),
.Y(n_903)
);

XNOR2xp5_ASAP7_75t_L g904 ( 
.A(n_902),
.B(n_154),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_899),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_898),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_900),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_901),
.A2(n_697),
.B(n_680),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_905),
.A2(n_896),
.B1(n_895),
.B2(n_816),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_903),
.A2(n_697),
.B(n_680),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_906),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_904),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_911),
.A2(n_907),
.B1(n_908),
.B2(n_750),
.Y(n_913)
);

AOI31xp33_ASAP7_75t_L g914 ( 
.A1(n_909),
.A2(n_155),
.A3(n_156),
.B(n_159),
.Y(n_914)
);

AOI211xp5_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_912),
.B(n_910),
.C(n_913),
.Y(n_915)
);

XOR2xp5_ASAP7_75t_L g916 ( 
.A(n_913),
.B(n_160),
.Y(n_916)
);

NAND4xp25_ASAP7_75t_L g917 ( 
.A(n_913),
.B(n_164),
.C(n_166),
.D(n_170),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_916),
.A2(n_171),
.B(n_172),
.Y(n_918)
);

OAI222xp33_ASAP7_75t_L g919 ( 
.A1(n_915),
.A2(n_719),
.B1(n_680),
.B2(n_681),
.C1(n_675),
.C2(n_702),
.Y(n_919)
);

NOR3xp33_ASAP7_75t_SL g920 ( 
.A(n_917),
.B(n_173),
.C(n_174),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_920),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_918),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_919),
.Y(n_923)
);

AOI221xp5_ASAP7_75t_L g924 ( 
.A1(n_921),
.A2(n_175),
.B1(n_176),
.B2(n_180),
.C(n_702),
.Y(n_924)
);

AOI211xp5_ASAP7_75t_L g925 ( 
.A1(n_924),
.A2(n_923),
.B(n_922),
.C(n_719),
.Y(n_925)
);


endmodule