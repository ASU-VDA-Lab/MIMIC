module real_aes_17166_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_874, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_874;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_617;
wire n_139;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g863 ( .A(n_0), .B(n_864), .Y(n_863) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_1), .A2(n_4), .B1(n_239), .B2(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g133 ( .A1(n_2), .A2(n_43), .B1(n_134), .B2(n_136), .Y(n_133) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_3), .A2(n_26), .B1(n_136), .B2(n_179), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_5), .A2(n_17), .B1(n_161), .B2(n_230), .Y(n_229) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_6), .A2(n_60), .B1(n_181), .B2(n_206), .Y(n_562) );
AOI22xp5_ASAP7_75t_L g615 ( .A1(n_7), .A2(n_18), .B1(n_134), .B2(n_165), .Y(n_615) );
INVx1_ASAP7_75t_L g864 ( .A(n_8), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g598 ( .A(n_9), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_10), .A2(n_102), .B1(n_856), .B2(n_870), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_11), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_12), .A2(n_19), .B1(n_163), .B2(n_205), .Y(n_204) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_13), .A2(n_86), .B1(n_117), .B2(n_118), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
OR2x2_ASAP7_75t_L g112 ( .A(n_14), .B(n_38), .Y(n_112) );
BUFx2_ASAP7_75t_L g869 ( .A(n_14), .Y(n_869) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_15), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_16), .Y(n_233) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_20), .A2(n_99), .B1(n_161), .B2(n_239), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_21), .A2(n_39), .B1(n_197), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_22), .B(n_162), .Y(n_194) );
OAI21x1_ASAP7_75t_L g150 ( .A1(n_23), .A2(n_57), .B(n_151), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g516 ( .A(n_24), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_25), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_27), .B(n_140), .Y(n_523) );
INVx4_ASAP7_75t_R g578 ( .A(n_28), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_29), .A2(n_47), .B1(n_142), .B2(n_144), .Y(n_141) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_30), .A2(n_53), .B1(n_144), .B2(n_161), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_31), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_32), .B(n_197), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_33), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_34), .B(n_136), .Y(n_530) );
INVx1_ASAP7_75t_L g539 ( .A(n_35), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_SL g596 ( .A1(n_36), .A2(n_134), .B(n_146), .C(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_37), .A2(n_54), .B1(n_134), .B2(n_144), .Y(n_512) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_38), .Y(n_867) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_40), .A2(n_85), .B1(n_134), .B2(n_178), .Y(n_177) );
AOI22x1_ASAP7_75t_SL g845 ( .A1(n_41), .A2(n_55), .B1(n_846), .B2(n_847), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_41), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_42), .A2(n_46), .B1(n_134), .B2(n_165), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_44), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g241 ( .A1(n_45), .A2(n_59), .B1(n_161), .B2(n_216), .Y(n_241) );
INVx1_ASAP7_75t_L g527 ( .A(n_48), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_49), .B(n_134), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_50), .Y(n_548) );
INVx2_ASAP7_75t_L g482 ( .A(n_51), .Y(n_482) );
INVx1_ASAP7_75t_L g110 ( .A(n_52), .Y(n_110) );
BUFx3_ASAP7_75t_L g490 ( .A(n_52), .Y(n_490) );
INVx1_ASAP7_75t_L g847 ( .A(n_55), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_56), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g616 ( .A1(n_58), .A2(n_87), .B1(n_134), .B2(n_144), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_61), .A2(n_73), .B1(n_142), .B2(n_216), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_62), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_63), .A2(n_75), .B1(n_134), .B2(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g160 ( .A1(n_64), .A2(n_97), .B1(n_161), .B2(n_163), .Y(n_160) );
AND2x4_ASAP7_75t_L g130 ( .A(n_65), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g151 ( .A(n_66), .Y(n_151) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_67), .A2(n_89), .B1(n_142), .B2(n_144), .Y(n_535) );
AO22x1_ASAP7_75t_L g565 ( .A1(n_68), .A2(n_74), .B1(n_227), .B2(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g131 ( .A(n_69), .Y(n_131) );
AND2x2_ASAP7_75t_L g599 ( .A(n_70), .B(n_148), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_71), .B(n_181), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g592 ( .A(n_72), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_76), .B(n_136), .Y(n_549) );
INVx2_ASAP7_75t_L g140 ( .A(n_77), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_78), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_79), .B(n_148), .Y(n_520) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_80), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g180 ( .A1(n_81), .A2(n_98), .B1(n_144), .B2(n_181), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_82), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_83), .B(n_158), .Y(n_563) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_84), .Y(n_153) );
INVx1_ASAP7_75t_L g118 ( .A(n_86), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_88), .B(n_148), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_90), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_91), .B(n_148), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g498 ( .A(n_92), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g849 ( .A(n_93), .Y(n_849) );
NAND2xp33_ASAP7_75t_L g198 ( .A(n_94), .B(n_162), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_95), .A2(n_167), .B(n_181), .C(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g580 ( .A(n_96), .B(n_581), .Y(n_580) );
NAND2xp33_ASAP7_75t_L g553 ( .A(n_100), .B(n_143), .Y(n_553) );
INVx4_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_483), .Y(n_103) );
A2O1A1O1Ixp25_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_113), .B(n_475), .C(n_478), .D(n_874), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
CKINVDCx8_ASAP7_75t_R g477 ( .A(n_107), .Y(n_477) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_110), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_111), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1_ASAP7_75t_L g855 ( .A(n_112), .B(n_490), .Y(n_855) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
XNOR2x1_ASAP7_75t_L g114 ( .A(n_115), .B(n_119), .Y(n_114) );
INVx2_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
OA22x2_ASAP7_75t_L g493 ( .A1(n_119), .A2(n_494), .B1(n_499), .B2(n_501), .Y(n_493) );
AND2x4_ASAP7_75t_L g119 ( .A(n_120), .B(n_371), .Y(n_119) );
NOR2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_323), .Y(n_120) );
NAND3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_270), .C(n_308), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_201), .B1(n_221), .B2(n_249), .C(n_255), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_123), .A2(n_448), .B1(n_451), .B2(n_452), .Y(n_447) );
INVx2_ASAP7_75t_SL g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_172), .Y(n_124) );
INVx1_ASAP7_75t_L g362 ( .A(n_125), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_154), .Y(n_125) );
INVx1_ASAP7_75t_L g314 ( .A(n_126), .Y(n_314) );
AND2x4_ASAP7_75t_L g357 ( .A(n_126), .B(n_278), .Y(n_357) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g285 ( .A(n_127), .B(n_188), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_127), .B(n_254), .Y(n_345) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g253 ( .A(n_128), .B(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g269 ( .A(n_128), .B(n_174), .Y(n_269) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_128), .Y(n_276) );
INVx1_ASAP7_75t_L g332 ( .A(n_128), .Y(n_332) );
AO31x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .A3(n_147), .B(n_152), .Y(n_128) );
INVx2_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
AO31x2_ASAP7_75t_L g202 ( .A1(n_129), .A2(n_156), .A3(n_203), .B(n_209), .Y(n_202) );
AO31x2_ASAP7_75t_L g224 ( .A1(n_129), .A2(n_175), .A3(n_225), .B(n_232), .Y(n_224) );
AO31x2_ASAP7_75t_L g613 ( .A1(n_129), .A2(n_220), .A3(n_614), .B(n_617), .Y(n_613) );
BUFx10_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g184 ( .A(n_130), .Y(n_184) );
BUFx10_ASAP7_75t_L g514 ( .A(n_130), .Y(n_514) );
INVx1_ASAP7_75t_L g569 ( .A(n_130), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B1(n_141), .B2(n_145), .Y(n_132) );
INVx1_ASAP7_75t_L g163 ( .A(n_134), .Y(n_163) );
INVx4_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
INVx1_ASAP7_75t_L g216 ( .A(n_134), .Y(n_216) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_135), .Y(n_136) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_135), .Y(n_144) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
INVx2_ASAP7_75t_L g179 ( .A(n_135), .Y(n_179) );
INVx1_ASAP7_75t_L g181 ( .A(n_135), .Y(n_181) );
INVx1_ASAP7_75t_L g207 ( .A(n_135), .Y(n_207) );
INVx1_ASAP7_75t_L g228 ( .A(n_135), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_135), .Y(n_231) );
INVx1_ASAP7_75t_L g240 ( .A(n_135), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_136), .B(n_592), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_137), .A2(n_145), .B1(n_215), .B2(n_217), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g225 ( .A1(n_137), .A2(n_145), .B1(n_226), .B2(n_229), .Y(n_225) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_137), .A2(n_145), .B1(n_238), .B2(n_241), .Y(n_237) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g513 ( .A(n_138), .Y(n_513) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g551 ( .A(n_139), .Y(n_551) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx8_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx1_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
INVx1_ASAP7_75t_L g526 ( .A(n_140), .Y(n_526) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_143), .A2(n_231), .B1(n_578), .B2(n_579), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_144), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g537 ( .A(n_144), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_145), .A2(n_160), .B1(n_164), .B2(n_166), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g176 ( .A1(n_145), .A2(n_177), .B1(n_180), .B2(n_182), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_145), .A2(n_196), .B(n_198), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_145), .A2(n_166), .B1(n_204), .B2(n_208), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_145), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_145), .A2(n_182), .B1(n_535), .B2(n_536), .Y(n_534) );
OAI22x1_ASAP7_75t_L g614 ( .A1(n_145), .A2(n_182), .B1(n_615), .B2(n_616), .Y(n_614) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
O2A1O1Ixp5_ASAP7_75t_L g192 ( .A1(n_146), .A2(n_165), .B(n_193), .C(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_146), .A2(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_146), .B(n_565), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g627 ( .A1(n_146), .A2(n_561), .B(n_565), .C(n_568), .Y(n_627) );
AO31x2_ASAP7_75t_L g509 ( .A1(n_147), .A2(n_510), .A3(n_514), .B(n_515), .Y(n_509) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
NOR2x1_ASAP7_75t_L g555 ( .A(n_148), .B(n_556), .Y(n_555) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_149), .B(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_149), .B(n_171), .Y(n_170) );
BUFx3_ASAP7_75t_L g175 ( .A(n_149), .Y(n_175) );
INVx2_ASAP7_75t_SL g190 ( .A(n_149), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_149), .B(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g531 ( .A(n_149), .B(n_514), .Y(n_531) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
INVx3_ASAP7_75t_L g252 ( .A(n_154), .Y(n_252) );
AND2x2_ASAP7_75t_L g267 ( .A(n_154), .B(n_188), .Y(n_267) );
INVx2_ASAP7_75t_L g273 ( .A(n_154), .Y(n_273) );
AND2x4_ASAP7_75t_L g335 ( .A(n_154), .B(n_174), .Y(n_335) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_154), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_154), .B(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
AND2x2_ASAP7_75t_L g284 ( .A(n_155), .B(n_174), .Y(n_284) );
AND2x2_ASAP7_75t_L g312 ( .A(n_155), .B(n_313), .Y(n_312) );
BUFx2_ASAP7_75t_L g391 ( .A(n_155), .Y(n_391) );
AO31x2_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_159), .A3(n_168), .B(n_170), .Y(n_155) );
AO31x2_ASAP7_75t_L g533 ( .A1(n_156), .A2(n_183), .A3(n_534), .B(n_538), .Y(n_533) );
AOI21x1_ASAP7_75t_L g588 ( .A1(n_156), .A2(n_589), .B(n_599), .Y(n_588) );
BUFx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_157), .B(n_516), .Y(n_515) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_157), .B(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g581 ( .A(n_157), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_157), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
INVx2_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
OAI21xp33_ASAP7_75t_L g568 ( .A1(n_158), .A2(n_563), .B(n_569), .Y(n_568) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_162), .Y(n_566) );
O2A1O1Ixp33_ASAP7_75t_L g547 ( .A1(n_165), .A2(n_548), .B(n_549), .C(n_550), .Y(n_547) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
INVx1_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
AO31x2_ASAP7_75t_L g236 ( .A1(n_168), .A2(n_212), .A3(n_237), .B(n_242), .Y(n_236) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g572 ( .A1(n_169), .A2(n_573), .B(n_576), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_188), .Y(n_172) );
INVx1_ASAP7_75t_L g347 ( .A(n_173), .Y(n_347) );
NAND2x1_ASAP7_75t_L g375 ( .A(n_173), .B(n_267), .Y(n_375) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OR2x2_ASAP7_75t_L g277 ( .A(n_174), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g313 ( .A(n_174), .Y(n_313) );
INVx1_ASAP7_75t_L g389 ( .A(n_174), .Y(n_389) );
AO31x2_ASAP7_75t_L g174 ( .A1(n_175), .A2(n_176), .A3(n_183), .B(n_185), .Y(n_174) );
INVx2_ASAP7_75t_SL g178 ( .A(n_179), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_179), .B(n_598), .Y(n_597) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_182), .B(n_577), .Y(n_576) );
AO31x2_ASAP7_75t_L g211 ( .A1(n_183), .A2(n_212), .A3(n_214), .B(n_218), .Y(n_211) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_SL g199 ( .A(n_184), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_SL g209 ( .A(n_186), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g213 ( .A(n_186), .Y(n_213) );
AND2x4_ASAP7_75t_L g328 ( .A(n_188), .B(n_313), .Y(n_328) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
BUFx2_ASAP7_75t_L g350 ( .A(n_189), .Y(n_350) );
OAI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B(n_200), .Y(n_189) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_190), .A2(n_191), .B(n_200), .Y(n_254) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_195), .B(n_199), .Y(n_191) );
AND2x4_ASAP7_75t_L g222 ( .A(n_201), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
INVx4_ASAP7_75t_SL g246 ( .A(n_202), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_202), .B(n_248), .Y(n_258) );
BUFx2_ASAP7_75t_L g322 ( .A(n_202), .Y(n_322) );
AND2x2_ASAP7_75t_L g366 ( .A(n_202), .B(n_224), .Y(n_366) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_207), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g244 ( .A(n_211), .Y(n_244) );
OR2x2_ASAP7_75t_L g282 ( .A(n_211), .B(n_224), .Y(n_282) );
INVx2_ASAP7_75t_L g293 ( .A(n_211), .Y(n_293) );
AND2x4_ASAP7_75t_L g296 ( .A(n_211), .B(n_297), .Y(n_296) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_211), .Y(n_337) );
INVx1_ASAP7_75t_L g378 ( .A(n_211), .Y(n_378) );
AO21x2_ASAP7_75t_L g571 ( .A1(n_212), .A2(n_572), .B(n_580), .Y(n_571) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_220), .B(n_243), .Y(n_242) );
OR2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_234), .Y(n_221) );
INVx2_ASAP7_75t_L g471 ( .A(n_222), .Y(n_471) );
AND2x4_ASAP7_75t_L g432 ( .A(n_223), .B(n_235), .Y(n_432) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
INVx2_ASAP7_75t_L g297 ( .A(n_224), .Y(n_297) );
INVx1_ASAP7_75t_L g353 ( .A(n_224), .Y(n_353) );
AND2x2_ASAP7_75t_L g379 ( .A(n_224), .B(n_304), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_224), .B(n_292), .Y(n_383) );
OAI21xp33_ASAP7_75t_SL g522 ( .A1(n_227), .A2(n_523), .B(n_524), .Y(n_522) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_245), .Y(n_234) );
INVx3_ASAP7_75t_L g360 ( .A(n_235), .Y(n_360) );
AND2x4_ASAP7_75t_L g235 ( .A(n_236), .B(n_244), .Y(n_235) );
INVx2_ASAP7_75t_L g264 ( .A(n_236), .Y(n_264) );
INVx2_ASAP7_75t_L g304 ( .A(n_236), .Y(n_304) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_240), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_244), .B(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g333 ( .A(n_244), .B(n_304), .Y(n_333) );
INVx1_ASAP7_75t_L g259 ( .A(n_245), .Y(n_259) );
NAND2x1_ASAP7_75t_L g395 ( .A(n_245), .B(n_369), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_245), .B(n_333), .Y(n_444) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx2_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_246), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g352 ( .A(n_246), .B(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_246), .Y(n_429) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_249), .A2(n_442), .B1(n_443), .B2(n_445), .Y(n_441) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_251), .B(n_285), .Y(n_320) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x4_ASAP7_75t_L g343 ( .A(n_252), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g442 ( .A(n_252), .B(n_253), .Y(n_442) );
AND2x2_ASAP7_75t_L g315 ( .A(n_253), .B(n_284), .Y(n_315) );
AND2x4_ASAP7_75t_L g334 ( .A(n_253), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g385 ( .A(n_253), .B(n_312), .Y(n_385) );
INVx1_ASAP7_75t_L g278 ( .A(n_254), .Y(n_278) );
AOI31xp33_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_259), .A3(n_260), .B(n_265), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_257), .B(n_300), .Y(n_299) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_257), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g469 ( .A1(n_257), .A2(n_259), .B(n_289), .Y(n_469) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g311 ( .A(n_258), .Y(n_311) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g446 ( .A(n_261), .B(n_282), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
INVx1_ASAP7_75t_L g301 ( .A(n_263), .Y(n_301) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_263), .Y(n_408) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g290 ( .A(n_264), .Y(n_290) );
OR2x2_ASAP7_75t_L g318 ( .A(n_264), .B(n_293), .Y(n_318) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NOR2x1p5_ASAP7_75t_L g307 ( .A(n_269), .B(n_273), .Y(n_307) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_279), .B1(n_283), .B2(n_286), .C(n_298), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g387 ( .A(n_276), .B(n_290), .Y(n_387) );
AND2x2_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
OR2x2_ASAP7_75t_L g317 ( .A(n_280), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g404 ( .A(n_280), .B(n_296), .Y(n_404) );
AND2x4_ASAP7_75t_L g321 ( .A(n_281), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g340 ( .A(n_282), .B(n_303), .Y(n_340) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_SL g356 ( .A(n_284), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_SL g397 ( .A(n_284), .Y(n_397) );
INVx2_ASAP7_75t_L g406 ( .A(n_284), .Y(n_406) );
AND2x2_ASAP7_75t_L g420 ( .A(n_284), .B(n_350), .Y(n_420) );
INVx1_ASAP7_75t_L g398 ( .A(n_285), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_287), .B(n_294), .Y(n_286) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_288), .B(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2x1p5_ASAP7_75t_L g330 ( .A(n_289), .B(n_296), .Y(n_330) );
AND2x2_ASAP7_75t_L g351 ( .A(n_289), .B(n_352), .Y(n_351) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_289), .B(n_321), .Y(n_459) );
INVx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B(n_306), .Y(n_298) );
NAND2x1_ASAP7_75t_L g460 ( .A(n_300), .B(n_404), .Y(n_460) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_301), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx4_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
AND2x2_ASAP7_75t_L g439 ( .A(n_303), .B(n_344), .Y(n_439) );
INVx3_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g336 ( .A(n_304), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g349 ( .A(n_307), .B(n_350), .Y(n_349) );
NOR2x1_ASAP7_75t_L g419 ( .A(n_307), .B(n_420), .Y(n_419) );
AOI322xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_312), .A3(n_314), .B1(n_315), .B2(n_316), .C1(n_319), .C2(n_321), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g402 ( .A(n_312), .B(n_350), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_312), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g426 ( .A(n_312), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g431 ( .A(n_312), .B(n_416), .Y(n_431) );
INVx1_ASAP7_75t_L g440 ( .A(n_312), .Y(n_440) );
OR2x2_ASAP7_75t_L g326 ( .A(n_314), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g453 ( .A(n_314), .Y(n_453) );
AND2x2_ASAP7_75t_L g456 ( .A(n_315), .B(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NOR3xp33_ASAP7_75t_L g392 ( .A(n_318), .B(n_332), .C(n_393), .Y(n_392) );
INVx2_ASAP7_75t_L g434 ( .A(n_318), .Y(n_434) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND3xp33_ASAP7_75t_SL g323 ( .A(n_324), .B(n_338), .C(n_348), .Y(n_323) );
AOI222xp33_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_329), .B1(n_331), .B2(n_333), .C1(n_334), .C2(n_336), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22x1_ASAP7_75t_L g470 ( .A1(n_327), .A2(n_471), .B1(n_472), .B2(n_473), .Y(n_470) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g331 ( .A(n_328), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_328), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g424 ( .A(n_328), .B(n_390), .Y(n_424) );
AND2x4_ASAP7_75t_L g454 ( .A(n_328), .B(n_391), .Y(n_454) );
AND2x2_ASAP7_75t_L g435 ( .A(n_329), .B(n_402), .Y(n_435) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g427 ( .A(n_332), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_333), .B(n_366), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_333), .B(n_352), .Y(n_450) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
INVx2_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
INVx1_ASAP7_75t_L g364 ( .A(n_337), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_343), .B(n_346), .Y(n_342) );
AOI221xp5_ASAP7_75t_SL g430 ( .A1(n_343), .A2(n_431), .B1(n_432), .B2(n_433), .C(n_435), .Y(n_430) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVxp67_ASAP7_75t_SL g468 ( .A(n_345), .Y(n_468) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_347), .B(n_453), .Y(n_462) );
AOI221xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_354), .B2(n_365), .C(n_367), .Y(n_348) );
OR2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_406), .Y(n_405) );
AOI32xp33_ASAP7_75t_L g386 ( .A1(n_352), .A2(n_366), .A3(n_387), .B1(n_388), .B2(n_392), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_352), .B(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_361), .B2(n_363), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_357), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR2x2_ASAP7_75t_L g428 ( .A(n_360), .B(n_429), .Y(n_428) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g421 ( .A(n_364), .B(n_366), .Y(n_421) );
AND2x2_ASAP7_75t_L g474 ( .A(n_364), .B(n_379), .Y(n_474) );
AND2x2_ASAP7_75t_L g433 ( .A(n_365), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_366), .B(n_369), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
NOR2x1_ASAP7_75t_L g371 ( .A(n_372), .B(n_436), .Y(n_371) );
NAND4xp75_ASAP7_75t_L g372 ( .A(n_373), .B(n_399), .C(n_417), .D(n_430), .Y(n_372) );
AOI211x1_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B(n_380), .C(n_394), .Y(n_373) );
INVxp67_ASAP7_75t_L g472 ( .A(n_374), .Y(n_472) );
INVx2_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_384), .B(n_386), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
BUFx2_ASAP7_75t_L g393 ( .A(n_389), .Y(n_393) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g465 ( .A(n_393), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .C(n_398), .Y(n_394) );
INVx2_ASAP7_75t_L g457 ( .A(n_395), .Y(n_457) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_409), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B1(n_405), .B2(n_407), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_414), .B2(n_415), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_422), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_425), .B(n_428), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_429), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g449 ( .A(n_432), .Y(n_449) );
NAND4xp75_ASAP7_75t_SL g436 ( .A(n_437), .B(n_447), .C(n_455), .D(n_463), .Y(n_436) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
NOR2xp67_ASAP7_75t_SL g455 ( .A(n_456), .B(n_458), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_461), .Y(n_458) );
INVxp67_ASAP7_75t_SL g461 ( .A(n_462), .Y(n_461) );
AOI21x1_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_469), .B(n_470), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
NOR2xp33_ASAP7_75t_SL g475 ( .A(n_476), .B(n_477), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_479), .Y(n_478) );
INVx2_ASAP7_75t_SL g479 ( .A(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g487 ( .A(n_482), .Y(n_487) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_482), .B(n_853), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_491), .B(n_848), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx6_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x6_ASAP7_75t_SL g486 ( .A(n_487), .B(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI22xp33_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B1(n_844), .B2(n_845), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx8_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx12f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_497), .Y(n_496) );
BUFx8_ASAP7_75t_SL g500 ( .A(n_497), .Y(n_500) );
AND2x2_ASAP7_75t_L g854 ( .A(n_497), .B(n_855), .Y(n_854) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
BUFx2_ASAP7_75t_L g862 ( .A(n_498), .Y(n_862) );
INVx3_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_734), .Y(n_501) );
NOR4xp25_ASAP7_75t_L g502 ( .A(n_503), .B(n_634), .C(n_676), .D(n_708), .Y(n_502) );
OAI211xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_540), .B(n_582), .C(n_619), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_517), .Y(n_506) );
INVx2_ASAP7_75t_L g647 ( .A(n_507), .Y(n_647) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g726 ( .A(n_508), .B(n_519), .Y(n_726) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_509), .B(n_533), .Y(n_585) );
AND2x2_ASAP7_75t_L g608 ( .A(n_509), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_SL g633 ( .A(n_509), .Y(n_633) );
OR2x2_ASAP7_75t_L g696 ( .A(n_509), .B(n_533), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_513), .A2(n_529), .B(n_530), .Y(n_528) );
OAI21x1_ASAP7_75t_L g561 ( .A1(n_513), .A2(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g556 ( .A(n_514), .Y(n_556) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x2_ASAP7_75t_L g630 ( .A(n_518), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g642 ( .A(n_518), .Y(n_642) );
INVxp67_ASAP7_75t_SL g820 ( .A(n_518), .Y(n_820) );
OR2x2_ASAP7_75t_L g833 ( .A(n_518), .B(n_834), .Y(n_833) );
OR2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_532), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_519), .B(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g606 ( .A(n_519), .Y(n_606) );
AND2x2_ASAP7_75t_L g653 ( .A(n_519), .B(n_654), .Y(n_653) );
NAND2x1p5_ASAP7_75t_SL g672 ( .A(n_519), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_519), .B(n_607), .Y(n_722) );
INVx1_ASAP7_75t_L g811 ( .A(n_519), .Y(n_811) );
AND2x2_ASAP7_75t_L g840 ( .A(n_519), .B(n_533), .Y(n_840) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_528), .B(n_531), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
BUFx4f_ASAP7_75t_L g595 ( .A(n_526), .Y(n_595) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g607 ( .A(n_533), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_533), .B(n_633), .Y(n_655) );
INVx1_ASAP7_75t_L g675 ( .A(n_533), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_533), .B(n_609), .Y(n_727) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_557), .Y(n_541) );
OR2x2_ASAP7_75t_L g624 ( .A(n_542), .B(n_625), .Y(n_624) );
OR2x2_ASAP7_75t_L g731 ( .A(n_542), .B(n_680), .Y(n_731) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g640 ( .A(n_543), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_543), .B(n_660), .Y(n_659) );
NOR2x1_ASAP7_75t_L g745 ( .A(n_543), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_L g603 ( .A(n_544), .Y(n_603) );
BUFx3_ASAP7_75t_L g651 ( .A(n_544), .Y(n_651) );
AND2x2_ASAP7_75t_L g687 ( .A(n_544), .B(n_668), .Y(n_687) );
AND2x2_ASAP7_75t_L g767 ( .A(n_544), .B(n_613), .Y(n_767) );
AND2x2_ASAP7_75t_L g780 ( .A(n_544), .B(n_571), .Y(n_780) );
NAND2x1p5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_552), .B(n_555), .Y(n_546) );
INVx2_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g720 ( .A(n_557), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_557), .B(n_650), .Y(n_728) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_570), .Y(n_557) );
AND2x2_ASAP7_75t_L g639 ( .A(n_558), .B(n_571), .Y(n_639) );
INVx1_ASAP7_75t_L g747 ( .A(n_558), .Y(n_747) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x4_ASAP7_75t_L g601 ( .A(n_559), .B(n_571), .Y(n_601) );
AND2x2_ASAP7_75t_L g664 ( .A(n_559), .B(n_570), .Y(n_664) );
AOI21x1_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B(n_567), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g589 ( .A1(n_569), .A2(n_590), .B(n_596), .Y(n_589) );
AND2x2_ASAP7_75t_L g622 ( .A(n_570), .B(n_613), .Y(n_622) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g612 ( .A(n_571), .B(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g680 ( .A(n_571), .B(n_613), .Y(n_680) );
INVx1_ASAP7_75t_L g691 ( .A(n_571), .Y(n_691) );
AND2x2_ASAP7_75t_L g754 ( .A(n_571), .B(n_603), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_600), .B1(n_604), .B2(n_610), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_583), .A2(n_653), .B1(n_656), .B2(n_658), .Y(n_652) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g732 ( .A(n_585), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g838 ( .A(n_585), .Y(n_838) );
INVx1_ASAP7_75t_L g697 ( .A(n_586), .Y(n_697) );
OR2x2_ASAP7_75t_L g760 ( .A(n_586), .B(n_655), .Y(n_760) );
OR2x2_ASAP7_75t_L g631 ( .A(n_587), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_587), .B(n_606), .Y(n_707) );
AND2x2_ASAP7_75t_L g724 ( .A(n_587), .B(n_651), .Y(n_724) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_587), .Y(n_741) );
INVxp67_ASAP7_75t_L g789 ( .A(n_587), .Y(n_789) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g609 ( .A(n_588), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g590 ( .A1(n_591), .A2(n_593), .B(n_595), .Y(n_590) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_601), .Y(n_699) );
INVx3_ASAP7_75t_L g704 ( .A(n_601), .Y(n_704) );
AND2x2_ASAP7_75t_L g717 ( .A(n_601), .B(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g817 ( .A(n_601), .B(n_779), .Y(n_817) );
INVx1_ASAP7_75t_L g611 ( .A(n_602), .Y(n_611) );
OR2x2_ASAP7_75t_L g794 ( .A(n_602), .B(n_769), .Y(n_794) );
BUFx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g718 ( .A(n_603), .B(n_628), .Y(n_718) );
AND2x2_ASAP7_75t_L g739 ( .A(n_603), .B(n_664), .Y(n_739) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_605), .B(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g740 ( .A(n_605), .Y(n_740) );
AND2x2_ASAP7_75t_L g782 ( .A(n_605), .B(n_783), .Y(n_782) );
AND2x4_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx2_ASAP7_75t_L g683 ( .A(n_606), .Y(n_683) );
AND2x2_ASAP7_75t_L g714 ( .A(n_606), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_606), .B(n_673), .Y(n_733) );
AND2x2_ASAP7_75t_L g682 ( .A(n_608), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g798 ( .A(n_608), .Y(n_798) );
AND2x2_ASAP7_75t_L g821 ( .A(n_608), .B(n_811), .Y(n_821) );
INVx1_ASAP7_75t_L g834 ( .A(n_608), .Y(n_834) );
INVx2_ASAP7_75t_L g673 ( .A(n_609), .Y(n_673) );
OR2x2_ASAP7_75t_L g769 ( .A(n_609), .B(n_633), .Y(n_769) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_612), .B(n_650), .Y(n_657) );
INVx2_ASAP7_75t_L g628 ( .A(n_613), .Y(n_628) );
INVx2_ASAP7_75t_L g668 ( .A(n_613), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_613), .B(n_626), .Y(n_690) );
OAI21xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_623), .B(n_629), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_622), .B(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g763 ( .A(n_625), .B(n_764), .Y(n_763) );
OR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx2_ASAP7_75t_L g669 ( .A(n_626), .Y(n_669) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g660 ( .A(n_628), .Y(n_660) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g643 ( .A(n_631), .Y(n_643) );
INVxp67_ASAP7_75t_L g814 ( .A(n_631), .Y(n_814) );
OR2x2_ASAP7_75t_L g716 ( .A(n_632), .B(n_673), .Y(n_716) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g634 ( .A(n_635), .B(n_644), .C(n_652), .D(n_661), .Y(n_634) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_641), .C(n_643), .Y(n_635) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g830 ( .A1(n_637), .A2(n_831), .B(n_833), .C(n_835), .Y(n_830) );
OR2x6_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_639), .B(n_687), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g742 ( .A(n_639), .B(n_743), .C(n_745), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_639), .B(n_718), .Y(n_823) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_639), .A2(n_744), .B1(n_836), .B2(n_839), .C(n_841), .Y(n_835) );
INVx1_ASAP7_75t_L g826 ( .A(n_640), .Y(n_826) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_648), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g761 ( .A1(n_645), .A2(n_653), .B1(n_688), .B2(n_762), .C(n_765), .Y(n_761) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_647), .B(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g712 ( .A(n_648), .Y(n_712) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_650), .B(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g827 ( .A(n_650), .B(n_678), .Y(n_827) );
INVx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g663 ( .A(n_651), .Y(n_663) );
AND3x1_ASAP7_75t_L g836 ( .A(n_651), .B(n_837), .C(n_838), .Y(n_836) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g706 ( .A(n_655), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g776 ( .A(n_658), .Y(n_776) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OR2x2_ASAP7_75t_L g752 ( .A(n_660), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g779 ( .A(n_660), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_670), .Y(n_661) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
NAND2x1_ASAP7_75t_L g677 ( .A(n_663), .B(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g744 ( .A(n_664), .Y(n_744) );
INVxp67_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_L g700 ( .A(n_668), .Y(n_700) );
OR2x2_ASAP7_75t_L g679 ( .A(n_669), .B(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g792 ( .A(n_669), .Y(n_792) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_671), .B(n_819), .Y(n_818) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_674), .Y(n_671) );
OR2x2_ASAP7_75t_L g748 ( .A(n_672), .B(n_696), .Y(n_748) );
INVx2_ASAP7_75t_L g837 ( .A(n_672), .Y(n_837) );
INVx1_ASAP7_75t_L g711 ( .A(n_673), .Y(n_711) );
NOR4xp25_ASAP7_75t_L g841 ( .A(n_673), .B(n_704), .C(n_842), .D(n_843), .Y(n_841) );
INVx1_ASAP7_75t_L g843 ( .A(n_674), .Y(n_843) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
BUFx3_ASAP7_75t_L g829 ( .A(n_675), .Y(n_829) );
OAI211xp5_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_681), .B(n_684), .C(n_692), .Y(n_676) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g816 ( .A(n_679), .Y(n_816) );
INVx2_ASAP7_75t_L g801 ( .A(n_680), .Y(n_801) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_682), .A2(n_685), .B(n_688), .Y(n_684) );
OR2x2_ASAP7_75t_L g768 ( .A(n_683), .B(n_769), .Y(n_768) );
AND2x2_ASAP7_75t_L g786 ( .A(n_683), .B(n_787), .Y(n_786) );
INVxp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g702 ( .A(n_687), .Y(n_702) );
AND2x4_ASAP7_75t_SL g791 ( .A(n_687), .B(n_792), .Y(n_791) );
INVx3_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_690), .Y(n_757) );
INVx1_ASAP7_75t_L g764 ( .A(n_691), .Y(n_764) );
AOI32xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_698), .A3(n_700), .B1(n_701), .B2(n_705), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_695), .B(n_711), .Y(n_710) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_695), .Y(n_756) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g773 ( .A(n_696), .B(n_711), .Y(n_773) );
INVx2_ASAP7_75t_L g787 ( .A(n_696), .Y(n_787) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_704), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI211xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_712), .B(n_713), .C(n_729), .Y(n_708) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_717), .B(n_719), .Y(n_713) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g770 ( .A(n_718), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_718), .B(n_805), .Y(n_804) );
OAI32xp33_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .A3(n_723), .B1(n_725), .B2(n_728), .Y(n_719) );
INVx1_ASAP7_75t_L g805 ( .A(n_720), .Y(n_805) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
OR2x2_ASAP7_75t_L g797 ( .A(n_722), .B(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
NOR2x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_806), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_736), .B(n_761), .C(n_774), .D(n_802), .Y(n_735) );
NOR2xp67_ASAP7_75t_L g736 ( .A(n_737), .B(n_749), .Y(n_736) );
OAI32xp33_ASAP7_75t_L g737 ( .A1(n_738), .A2(n_740), .A3(n_741), .B1(n_742), .B2(n_748), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g788 ( .A(n_740), .B(n_789), .Y(n_788) );
OAI32xp33_ASAP7_75t_L g793 ( .A1(n_740), .A2(n_794), .A3(n_795), .B1(n_797), .B2(n_799), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_741), .B(n_829), .Y(n_828) );
NAND2xp5_ASAP7_75t_SL g807 ( .A(n_743), .B(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g800 ( .A(n_746), .B(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g832 ( .A(n_746), .Y(n_832) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g796 ( .A(n_747), .Y(n_796) );
OAI22x1_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_755), .B1(n_757), .B2(n_758), .Y(n_749) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_759), .B(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NOR2x1_ASAP7_75t_L g825 ( .A(n_763), .B(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_770), .B2(n_771), .Y(n_765) );
NAND2x1_ASAP7_75t_L g831 ( .A(n_767), .B(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g842 ( .A(n_767), .Y(n_842) );
INVx2_ASAP7_75t_L g783 ( .A(n_769), .Y(n_783) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
NOR3xp33_ASAP7_75t_SL g774 ( .A(n_775), .B(n_784), .C(n_793), .Y(n_774) );
AOI21xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_777), .B(n_781), .Y(n_775) );
NAND2xp33_ASAP7_75t_L g803 ( .A(n_777), .B(n_804), .Y(n_803) );
INVx2_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
AND2x4_ASAP7_75t_L g839 ( .A(n_783), .B(n_840), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_788), .B(n_790), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x4_ASAP7_75t_L g810 ( .A(n_787), .B(n_811), .Y(n_810) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_789), .Y(n_809) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVxp67_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND3xp33_ASAP7_75t_SL g806 ( .A(n_807), .B(n_812), .C(n_824), .Y(n_806) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g815 ( .A(n_811), .Y(n_815) );
AOI222xp33_ASAP7_75t_L g812 ( .A1(n_813), .A2(n_816), .B1(n_817), .B2(n_818), .C1(n_821), .C2(n_822), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
O2A1O1Ixp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_827), .B(n_828), .C(n_830), .Y(n_824) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx6_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
BUFx10_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
CKINVDCx11_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
OR2x6_ASAP7_75t_L g857 ( .A(n_858), .B(n_865), .Y(n_857) );
OR2x6_ASAP7_75t_L g872 ( .A(n_858), .B(n_865), .Y(n_872) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2x1p5_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
NOR2x1p5_ASAP7_75t_L g866 ( .A(n_867), .B(n_868), .Y(n_866) );
INVx1_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
INVx3_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
CKINVDCx11_ASAP7_75t_R g871 ( .A(n_872), .Y(n_871) );
endmodule