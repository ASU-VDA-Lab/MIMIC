module fake_ariane_633_n_1468 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_332, n_294, n_197, n_176, n_34, n_404, n_172, n_347, n_183, n_373, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_416, n_283, n_50, n_187, n_367, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_57, n_387, n_406, n_117, n_139, n_85, n_130, n_349, n_391, n_346, n_214, n_348, n_2, n_32, n_410, n_379, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_405, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_401, n_267, n_335, n_350, n_291, n_344, n_381, n_398, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_365, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_390, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_388, n_333, n_413, n_392, n_376, n_221, n_321, n_86, n_361, n_89, n_149, n_383, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_362, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_371, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_414, n_287, n_302, n_380, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_409, n_171, n_384, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_407, n_13, n_27, n_254, n_219, n_55, n_231, n_366, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_415, n_78, n_63, n_99, n_216, n_5, n_223, n_403, n_25, n_83, n_389, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_378, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_358, n_105, n_30, n_131, n_263, n_360, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_364, n_258, n_118, n_121, n_411, n_353, n_22, n_241, n_29, n_357, n_412, n_191, n_382, n_80, n_211, n_97, n_408, n_322, n_251, n_116, n_397, n_351, n_39, n_393, n_359, n_155, n_127, n_1468);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_183;
input n_373;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_367;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_57;
input n_387;
input n_406;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_391;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_410;
input n_379;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_405;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_401;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_381;
input n_398;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_365;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_413;
input n_392;
input n_376;
input n_221;
input n_321;
input n_86;
input n_361;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_362;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_414;
input n_287;
input n_302;
input n_380;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_409;
input n_171;
input n_384;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_407;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_366;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_378;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_358;
input n_105;
input n_30;
input n_131;
input n_263;
input n_360;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_364;
input n_258;
input n_118;
input n_121;
input n_411;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_191;
input n_382;
input n_80;
input n_211;
input n_97;
input n_408;
input n_322;
input n_251;
input n_116;
input n_397;
input n_351;
input n_39;
input n_393;
input n_359;
input n_155;
input n_127;

output n_1468;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_1013;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_1352;
wire n_643;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_519;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_826;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_917;
wire n_1271;
wire n_631;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_946;
wire n_757;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_849;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_1451;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_227),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_192),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_247),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_315),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_49),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_13),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_305),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_112),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

BUFx5_ASAP7_75t_L g426 ( 
.A(n_299),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_385),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_337),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_125),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_207),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_67),
.Y(n_432)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_39),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_150),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_160),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_82),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_267),
.Y(n_438)
);

BUFx2_ASAP7_75t_L g439 ( 
.A(n_231),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_334),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_114),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_265),
.Y(n_442)
);

BUFx10_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_253),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_111),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_203),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_127),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_390),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_393),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_68),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_270),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_55),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_213),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_196),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_45),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_141),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_322),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_273),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_255),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_54),
.Y(n_461)
);

BUFx2_ASAP7_75t_SL g462 ( 
.A(n_193),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_271),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_29),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_122),
.B(n_90),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_278),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_110),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_48),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_183),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_54),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_304),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_38),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_399),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_409),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_200),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_113),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_47),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_182),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_232),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_256),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_94),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_204),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_11),
.Y(n_483)
);

INVx2_ASAP7_75t_SL g484 ( 
.A(n_220),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_178),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_371),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_238),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_306),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_246),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_236),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_339),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_109),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_35),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_149),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_292),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_283),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_300),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_261),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_389),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_272),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_32),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_205),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_152),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_190),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_310),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_40),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_189),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_403),
.Y(n_508)
);

BUFx10_ASAP7_75t_L g509 ( 
.A(n_266),
.Y(n_509)
);

INVx1_ASAP7_75t_SL g510 ( 
.A(n_296),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_155),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_294),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_153),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_307),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_326),
.Y(n_515)
);

BUFx3_ASAP7_75t_L g516 ( 
.A(n_115),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_187),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_128),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_75),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_228),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_291),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_214),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_169),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_41),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_199),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_248),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_15),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_70),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_309),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_78),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_38),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_416),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_244),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_344),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_327),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_70),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_191),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_188),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_108),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_368),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_99),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_404),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_6),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_280),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_351),
.Y(n_545)
);

BUFx5_ASAP7_75t_L g546 ( 
.A(n_340),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_317),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_275),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_215),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_355),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g551 ( 
.A(n_26),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_384),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_262),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_313),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_161),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_148),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_245),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_46),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_171),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_250),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_202),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_151),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_348),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_230),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_185),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_5),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_36),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_222),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_13),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_51),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_15),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_314),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_302),
.Y(n_573)
);

CKINVDCx16_ASAP7_75t_R g574 ( 
.A(n_224),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_34),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_100),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_359),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_154),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_360),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_45),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_27),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_86),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_118),
.Y(n_583)
);

NOR2xp67_ASAP7_75t_L g584 ( 
.A(n_60),
.B(n_373),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_412),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_440),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_461),
.Y(n_587)
);

OA21x2_ASAP7_75t_L g588 ( 
.A1(n_420),
.A2(n_0),
.B(n_1),
.Y(n_588)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_551),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_434),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_485),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_456),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_434),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_466),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_501),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_476),
.Y(n_596)
);

BUFx8_ASAP7_75t_SL g597 ( 
.A(n_452),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_572),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_582),
.Y(n_599)
);

BUFx8_ASAP7_75t_SL g600 ( 
.A(n_524),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_476),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_572),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g603 ( 
.A(n_433),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_516),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_516),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_578),
.B(n_2),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_421),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_485),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_444),
.Y(n_610)
);

INVx5_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_485),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_575),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_469),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_580),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_439),
.Y(n_616)
);

INVx3_ASAP7_75t_L g617 ( 
.A(n_576),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_582),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_618)
);

BUFx12f_ASAP7_75t_L g619 ( 
.A(n_443),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_578),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_468),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_509),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_521),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_425),
.B(n_7),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_427),
.B(n_8),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_492),
.B(n_9),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_430),
.B(n_10),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_487),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_487),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_487),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_499),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_481),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_431),
.B(n_10),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_11),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_438),
.B(n_12),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_506),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_569),
.Y(n_637)
);

OA21x2_ASAP7_75t_L g638 ( 
.A1(n_442),
.A2(n_447),
.B(n_446),
.Y(n_638)
);

AND2x6_ASAP7_75t_L g639 ( 
.A(n_547),
.B(n_116),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_517),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_547),
.Y(n_642)
);

HB1xp67_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_547),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_529),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_547),
.B(n_117),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_455),
.B(n_12),
.Y(n_647)
);

OAI22x1_ASAP7_75t_R g648 ( 
.A1(n_422),
.A2(n_17),
.B1(n_14),
.B2(n_16),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_532),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_571),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_457),
.B(n_14),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_458),
.B(n_471),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_473),
.Y(n_654)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_557),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_655)
);

AND2x6_ASAP7_75t_L g656 ( 
.A(n_453),
.B(n_119),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_429),
.B(n_18),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_554),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_474),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_475),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_591),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_610),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_586),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_614),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_589),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_R g666 ( 
.A(n_587),
.B(n_432),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_445),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_591),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_631),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_640),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_593),
.Y(n_671)
);

NAND2xp33_ASAP7_75t_L g672 ( 
.A(n_606),
.B(n_465),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_591),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_R g674 ( 
.A(n_645),
.B(n_574),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_R g675 ( 
.A(n_641),
.B(n_417),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_621),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_636),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g678 ( 
.A(n_597),
.Y(n_678)
);

BUFx10_ASAP7_75t_L g679 ( 
.A(n_653),
.Y(n_679)
);

CKINVDCx20_ASAP7_75t_R g680 ( 
.A(n_600),
.Y(n_680)
);

CKINVDCx20_ASAP7_75t_R g681 ( 
.A(n_619),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_603),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_649),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_616),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_608),
.Y(n_685)
);

BUFx6f_ASAP7_75t_L g686 ( 
.A(n_608),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_623),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_649),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_658),
.B(n_622),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_650),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_649),
.Y(n_691)
);

INVxp33_ASAP7_75t_SL g692 ( 
.A(n_655),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_658),
.Y(n_693)
);

CKINVDCx16_ASAP7_75t_R g694 ( 
.A(n_599),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_590),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_594),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_654),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_596),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_608),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_R g700 ( 
.A(n_638),
.B(n_598),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_601),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_604),
.Y(n_702)
);

NAND2xp33_ASAP7_75t_R g703 ( 
.A(n_638),
.B(n_437),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_R g704 ( 
.A(n_602),
.B(n_418),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_648),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_605),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_R g707 ( 
.A(n_620),
.B(n_450),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_667),
.B(n_695),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_672),
.B(n_657),
.C(n_606),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_698),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_704),
.B(n_657),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_667),
.B(n_676),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_671),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_683),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_677),
.B(n_652),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_693),
.B(n_652),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_697),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_696),
.B(n_629),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_701),
.B(n_629),
.Y(n_719)
);

NAND3xp33_ASAP7_75t_L g720 ( 
.A(n_707),
.B(n_626),
.C(n_635),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_661),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_675),
.B(n_634),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_668),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_705),
.B(n_613),
.C(n_592),
.Y(n_724)
);

AO221x1_ASAP7_75t_L g725 ( 
.A1(n_692),
.A2(n_615),
.B1(n_618),
.B2(n_459),
.C(n_654),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_679),
.B(n_659),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_673),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_682),
.Y(n_728)
);

NOR2xp67_ASAP7_75t_L g729 ( 
.A(n_684),
.B(n_660),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_679),
.B(n_624),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_702),
.B(n_624),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_706),
.B(n_625),
.Y(n_732)
);

NAND2xp33_ASAP7_75t_L g733 ( 
.A(n_689),
.B(n_627),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_687),
.B(n_643),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_690),
.B(n_627),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_699),
.B(n_633),
.Y(n_736)
);

INVxp33_ASAP7_75t_L g737 ( 
.A(n_674),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_700),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_665),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_688),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_691),
.B(n_633),
.Y(n_741)
);

INVxp33_ASAP7_75t_L g742 ( 
.A(n_694),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_685),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_662),
.B(n_643),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_685),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_664),
.B(n_647),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_685),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_685),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_686),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_686),
.B(n_651),
.Y(n_750)
);

NAND3xp33_ASAP7_75t_L g751 ( 
.A(n_666),
.B(n_651),
.C(n_470),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_686),
.B(n_656),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_686),
.B(n_656),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_670),
.B(n_607),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_681),
.B(n_595),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_703),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_703),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_663),
.B(n_472),
.Y(n_758)
);

NOR3xp33_ASAP7_75t_L g759 ( 
.A(n_669),
.B(n_483),
.C(n_477),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_678),
.B(n_609),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_680),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_665),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_693),
.B(n_632),
.Y(n_763)
);

BUFx6f_ASAP7_75t_L g764 ( 
.A(n_685),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_698),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_693),
.B(n_637),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_667),
.B(n_656),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_667),
.B(n_611),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_667),
.B(n_611),
.Y(n_769)
);

INVx8_ASAP7_75t_L g770 ( 
.A(n_682),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_698),
.Y(n_771)
);

INVx1_ASAP7_75t_SL g772 ( 
.A(n_744),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_713),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_731),
.B(n_510),
.Y(n_774)
);

INVx2_ASAP7_75t_SL g775 ( 
.A(n_734),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_717),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_746),
.B(n_519),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_720),
.A2(n_584),
.B1(n_463),
.B2(n_484),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_730),
.B(n_527),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_716),
.B(n_528),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_770),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_741),
.B(n_530),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_770),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_750),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_741),
.B(n_531),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_764),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_750),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_765),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_764),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_721),
.Y(n_790)
);

AND2x6_ASAP7_75t_SL g791 ( 
.A(n_760),
.B(n_480),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_736),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_739),
.B(n_757),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_736),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_770),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_768),
.A2(n_769),
.B(n_767),
.Y(n_796)
);

INVx2_ASAP7_75t_SL g797 ( 
.A(n_755),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_754),
.B(n_617),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_712),
.B(n_708),
.Y(n_799)
);

INVx3_ASAP7_75t_L g800 ( 
.A(n_748),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_723),
.Y(n_801)
);

BUFx8_ASAP7_75t_SL g802 ( 
.A(n_761),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_771),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_725),
.A2(n_588),
.B1(n_462),
.B2(n_577),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_729),
.B(n_536),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_764),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_711),
.A2(n_491),
.B1(n_494),
.B2(n_488),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_748),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_710),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_757),
.Y(n_810)
);

AND2x6_ASAP7_75t_SL g811 ( 
.A(n_763),
.B(n_496),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_727),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_756),
.A2(n_646),
.B1(n_639),
.B2(n_502),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_708),
.B(n_541),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_732),
.B(n_543),
.Y(n_815)
);

OAI22xp33_ASAP7_75t_L g816 ( 
.A1(n_751),
.A2(n_566),
.B1(n_567),
.B2(n_558),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_762),
.B(n_581),
.Y(n_817)
);

INVx1_ASAP7_75t_SL g818 ( 
.A(n_742),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_715),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_737),
.B(n_500),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_718),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_766),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_SL g823 ( 
.A(n_724),
.B(n_423),
.C(n_419),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_757),
.A2(n_646),
.B1(n_639),
.B2(n_505),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_735),
.B(n_424),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_715),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_714),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_745),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_749),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_726),
.Y(n_830)
);

BUFx4f_ASAP7_75t_L g831 ( 
.A(n_740),
.Y(n_831)
);

AND2x6_ASAP7_75t_L g832 ( 
.A(n_767),
.B(n_507),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_738),
.B(n_428),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_SL g834 ( 
.A(n_759),
.B(n_436),
.C(n_435),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_747),
.Y(n_835)
);

INVx3_ASAP7_75t_L g836 ( 
.A(n_747),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_743),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_733),
.B(n_719),
.Y(n_838)
);

INVx1_ASAP7_75t_SL g839 ( 
.A(n_722),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_752),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_758),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_753),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_768),
.B(n_769),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_720),
.A2(n_512),
.B1(n_513),
.B2(n_511),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_713),
.Y(n_845)
);

HB1xp67_ASAP7_75t_L g846 ( 
.A(n_734),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_746),
.B(n_441),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_R g848 ( 
.A(n_762),
.B(n_448),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_731),
.B(n_449),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_713),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_709),
.A2(n_523),
.B1(n_533),
.B2(n_522),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_746),
.B(n_451),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_720),
.A2(n_540),
.B1(n_549),
.B2(n_537),
.Y(n_853)
);

INVx5_ASAP7_75t_L g854 ( 
.A(n_770),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_720),
.A2(n_555),
.B1(n_559),
.B2(n_552),
.Y(n_855)
);

INVx2_ASAP7_75t_SL g856 ( 
.A(n_744),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_729),
.B(n_561),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_713),
.Y(n_858)
);

AND2x4_ASAP7_75t_L g859 ( 
.A(n_729),
.B(n_562),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_770),
.Y(n_860)
);

AO22x1_ASAP7_75t_L g861 ( 
.A1(n_724),
.A2(n_646),
.B1(n_639),
.B2(n_564),
.Y(n_861)
);

AND2x4_ASAP7_75t_SL g862 ( 
.A(n_728),
.B(n_563),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_770),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_731),
.B(n_454),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_750),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_746),
.B(n_565),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_750),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_731),
.B(n_460),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_770),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_SL g870 ( 
.A1(n_777),
.A2(n_482),
.B(n_539),
.C(n_467),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_819),
.B(n_478),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_866),
.A2(n_646),
.B1(n_560),
.B2(n_479),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_826),
.B(n_486),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_856),
.B(n_490),
.C(n_489),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_843),
.A2(n_497),
.B(n_495),
.Y(n_875)
);

INVx6_ASAP7_75t_L g876 ( 
.A(n_854),
.Y(n_876)
);

BUFx10_ASAP7_75t_L g877 ( 
.A(n_783),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_854),
.B(n_498),
.Y(n_878)
);

O2A1O1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_814),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_796),
.A2(n_504),
.B(n_503),
.Y(n_880)
);

CKINVDCx8_ASAP7_75t_R g881 ( 
.A(n_854),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_792),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_772),
.Y(n_883)
);

NAND2x1p5_ASAP7_75t_L g884 ( 
.A(n_795),
.B(n_611),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_SL g885 ( 
.A(n_860),
.B(n_514),
.C(n_508),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_774),
.B(n_515),
.Y(n_886)
);

O2A1O1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_794),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_838),
.A2(n_867),
.B(n_865),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_865),
.A2(n_520),
.B(n_518),
.Y(n_889)
);

AO32x1_ASAP7_75t_L g890 ( 
.A1(n_851),
.A2(n_546),
.A3(n_426),
.B1(n_27),
.B2(n_25),
.Y(n_890)
);

XNOR2xp5_ASAP7_75t_L g891 ( 
.A(n_869),
.B(n_525),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_822),
.B(n_526),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_R g893 ( 
.A(n_781),
.B(n_534),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_830),
.B(n_535),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_784),
.B(n_538),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_804),
.A2(n_542),
.B1(n_545),
.B2(n_544),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_839),
.B(n_775),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_863),
.B(n_28),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_849),
.A2(n_550),
.B1(n_553),
.B2(n_548),
.Y(n_899)
);

BUFx8_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_845),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_846),
.B(n_30),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_831),
.B(n_556),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_863),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_786),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_802),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_864),
.A2(n_573),
.B1(n_579),
.B2(n_568),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_821),
.B(n_583),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_SL g909 ( 
.A(n_834),
.B(n_585),
.C(n_30),
.Y(n_909)
);

OAI21xp5_ASAP7_75t_L g910 ( 
.A1(n_840),
.A2(n_630),
.B(n_546),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_841),
.B(n_31),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_776),
.Y(n_912)
);

AOI22x1_ASAP7_75t_L g913 ( 
.A1(n_867),
.A2(n_628),
.B1(n_642),
.B2(n_612),
.Y(n_913)
);

OAI22x1_ASAP7_75t_L g914 ( 
.A1(n_807),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_787),
.A2(n_630),
.B(n_628),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_818),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_798),
.B(n_33),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_868),
.B(n_37),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_786),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_848),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_780),
.B(n_37),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_793),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_850),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_858),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_789),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_801),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_825),
.A2(n_815),
.B1(n_852),
.B2(n_847),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_810),
.B(n_39),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_817),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_803),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_810),
.B(n_42),
.Y(n_931)
);

NOR3xp33_ASAP7_75t_SL g932 ( 
.A(n_823),
.B(n_43),
.C(n_44),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_820),
.A2(n_546),
.B1(n_426),
.B2(n_644),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_844),
.A2(n_642),
.B(n_644),
.C(n_612),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_R g935 ( 
.A(n_805),
.B(n_120),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_853),
.B(n_43),
.Y(n_936)
);

A2O1A1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_855),
.A2(n_644),
.B(n_48),
.C(n_46),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_857),
.A2(n_546),
.B1(n_426),
.B2(n_50),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_859),
.B(n_49),
.Y(n_939)
);

INVx6_ASAP7_75t_L g940 ( 
.A(n_791),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_837),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_790),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_862),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_835),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_789),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_812),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_782),
.B(n_51),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_831),
.B(n_426),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_785),
.B(n_52),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_805),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_789),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_842),
.A2(n_546),
.B(n_426),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_779),
.A2(n_778),
.B1(n_836),
.B2(n_808),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_827),
.B(n_53),
.Y(n_954)
);

OAI22xp5_ASAP7_75t_L g955 ( 
.A1(n_836),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_809),
.B(n_56),
.Y(n_956)
);

INVxp33_ASAP7_75t_SL g957 ( 
.A(n_833),
.Y(n_957)
);

BUFx12f_ASAP7_75t_L g958 ( 
.A(n_811),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_806),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_800),
.B(n_58),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_788),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_806),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_832),
.B(n_59),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_828),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_829),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_816),
.B(n_60),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_813),
.A2(n_824),
.B(n_832),
.C(n_63),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_832),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_832),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_861),
.B(n_61),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_866),
.A2(n_64),
.B(n_62),
.C(n_63),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_819),
.B(n_62),
.Y(n_972)
);

NAND3xp33_ASAP7_75t_SL g973 ( 
.A(n_777),
.B(n_64),
.C(n_65),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_R g974 ( 
.A(n_783),
.B(n_121),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_819),
.B(n_65),
.Y(n_975)
);

INVxp67_ASAP7_75t_SL g976 ( 
.A(n_786),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_799),
.A2(n_124),
.B(n_123),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_799),
.B(n_66),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_799),
.B(n_66),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_799),
.B(n_67),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_819),
.B(n_69),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_799),
.B(n_69),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_863),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_799),
.A2(n_129),
.B(n_126),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_866),
.A2(n_73),
.B(n_71),
.C(n_72),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_799),
.B(n_71),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_772),
.B(n_72),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_799),
.A2(n_131),
.B(n_130),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_799),
.A2(n_133),
.B(n_132),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_799),
.B(n_73),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_772),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_799),
.A2(n_135),
.B(n_134),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_819),
.B(n_74),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_819),
.B(n_74),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_866),
.A2(n_77),
.B(n_75),
.C(n_76),
.Y(n_995)
);

BUFx10_ASAP7_75t_L g996 ( 
.A(n_783),
.Y(n_996)
);

A2O1A1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_866),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_863),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_773),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_799),
.A2(n_137),
.B(n_136),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_799),
.B(n_79),
.Y(n_1001)
);

O2A1O1Ixp5_ASAP7_75t_L g1002 ( 
.A1(n_866),
.A2(n_81),
.B(n_79),
.C(n_80),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_773),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_819),
.B(n_81),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_799),
.A2(n_84),
.B1(n_82),
.B2(n_83),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_799),
.B(n_84),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_772),
.B(n_85),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_866),
.A2(n_89),
.B(n_87),
.C(n_88),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_R g1009 ( 
.A(n_783),
.B(n_138),
.Y(n_1009)
);

OR2x6_ASAP7_75t_L g1010 ( 
.A(n_863),
.B(n_88),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_R g1011 ( 
.A(n_783),
.B(n_139),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_772),
.B(n_90),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_L g1013 ( 
.A1(n_777),
.A2(n_91),
.B(n_92),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_819),
.B(n_91),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_866),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_772),
.B(n_95),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_952),
.A2(n_142),
.B(n_140),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_883),
.Y(n_1018)
);

OR2x6_ASAP7_75t_L g1019 ( 
.A(n_906),
.B(n_1010),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_SL g1020 ( 
.A1(n_888),
.A2(n_96),
.B(n_97),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_916),
.B(n_991),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_969),
.A2(n_144),
.B(n_143),
.Y(n_1022)
);

NAND2x1p5_ASAP7_75t_L g1023 ( 
.A(n_922),
.B(n_145),
.Y(n_1023)
);

AO21x2_ASAP7_75t_L g1024 ( 
.A1(n_910),
.A2(n_147),
.B(n_146),
.Y(n_1024)
);

BUFx5_ASAP7_75t_L g1025 ( 
.A(n_926),
.Y(n_1025)
);

BUFx12f_ASAP7_75t_L g1026 ( 
.A(n_996),
.Y(n_1026)
);

AOI22x1_ASAP7_75t_L g1027 ( 
.A1(n_977),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1027)
);

INVx1_ASAP7_75t_SL g1028 ( 
.A(n_929),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_941),
.Y(n_1029)
);

BUFx3_ASAP7_75t_L g1030 ( 
.A(n_900),
.Y(n_1030)
);

OAI21x1_ASAP7_75t_L g1031 ( 
.A1(n_984),
.A2(n_157),
.B(n_156),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_988),
.A2(n_159),
.B(n_158),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_876),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_1016),
.B(n_98),
.Y(n_1034)
);

INVx8_ASAP7_75t_L g1035 ( 
.A(n_1010),
.Y(n_1035)
);

AOI22x1_ASAP7_75t_L g1036 ( 
.A1(n_989),
.A2(n_1000),
.B1(n_992),
.B2(n_875),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_959),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_901),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_915),
.A2(n_163),
.B(n_162),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_996),
.Y(n_1040)
);

INVx6_ASAP7_75t_SL g1041 ( 
.A(n_877),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_876),
.Y(n_1042)
);

NAND2x1p5_ASAP7_75t_L g1043 ( 
.A(n_944),
.B(n_164),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_900),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_923),
.Y(n_1045)
);

BUFx2_ASAP7_75t_SL g1046 ( 
.A(n_881),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_920),
.Y(n_1047)
);

AOI22x1_ASAP7_75t_L g1048 ( 
.A1(n_880),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_930),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_SL g1050 ( 
.A1(n_978),
.A2(n_980),
.B(n_979),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_928),
.A2(n_166),
.B(n_165),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_959),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_912),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_959),
.B(n_167),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_898),
.Y(n_1055)
);

OR2x6_ASAP7_75t_L g1056 ( 
.A(n_950),
.B(n_940),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_957),
.B(n_102),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_924),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_966),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_964),
.Y(n_1060)
);

OAI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_982),
.A2(n_104),
.B(n_105),
.Y(n_1061)
);

OA21x2_ASAP7_75t_L g1062 ( 
.A1(n_918),
.A2(n_170),
.B(n_168),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_894),
.B(n_105),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_SL g1064 ( 
.A(n_968),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_942),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_931),
.A2(n_173),
.B(n_172),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_987),
.B(n_1007),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_905),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_986),
.A2(n_106),
.B(n_107),
.Y(n_1069)
);

BUFx4f_ASAP7_75t_SL g1070 ( 
.A(n_943),
.Y(n_1070)
);

OA21x2_ASAP7_75t_L g1071 ( 
.A1(n_913),
.A2(n_175),
.B(n_174),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_SL g1072 ( 
.A1(n_990),
.A2(n_106),
.B(n_107),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_999),
.Y(n_1073)
);

CKINVDCx20_ASAP7_75t_R g1074 ( 
.A(n_891),
.Y(n_1074)
);

OAI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1001),
.A2(n_176),
.B(n_177),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_967),
.A2(n_179),
.B(n_180),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_940),
.Y(n_1077)
);

NAND2x1p5_ASAP7_75t_L g1078 ( 
.A(n_904),
.B(n_181),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1003),
.Y(n_1079)
);

CKINVDCx8_ASAP7_75t_R g1080 ( 
.A(n_897),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_905),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_983),
.B(n_184),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_956),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_946),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_974),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_965),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_905),
.Y(n_1087)
);

INVx6_ASAP7_75t_L g1088 ( 
.A(n_958),
.Y(n_1088)
);

INVx5_ASAP7_75t_L g1089 ( 
.A(n_968),
.Y(n_1089)
);

INVx3_ASAP7_75t_SL g1090 ( 
.A(n_902),
.Y(n_1090)
);

NAND2x1p5_ASAP7_75t_L g1091 ( 
.A(n_998),
.B(n_186),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1012),
.B(n_415),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1006),
.Y(n_1093)
);

AOI21x1_ASAP7_75t_L g1094 ( 
.A1(n_927),
.A2(n_194),
.B(n_195),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_953),
.A2(n_197),
.B(n_198),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_954),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_908),
.B(n_201),
.Y(n_1097)
);

AO21x2_ASAP7_75t_L g1098 ( 
.A1(n_933),
.A2(n_206),
.B(n_208),
.Y(n_1098)
);

AO21x2_ASAP7_75t_L g1099 ( 
.A1(n_948),
.A2(n_209),
.B(n_210),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_884),
.Y(n_1100)
);

OAI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_873),
.A2(n_211),
.B(n_212),
.Y(n_1101)
);

CKINVDCx6p67_ASAP7_75t_R g1102 ( 
.A(n_914),
.Y(n_1102)
);

INVx6_ASAP7_75t_L g1103 ( 
.A(n_919),
.Y(n_1103)
);

BUFx12f_ASAP7_75t_L g1104 ( 
.A(n_919),
.Y(n_1104)
);

INVx2_ASAP7_75t_SL g1105 ( 
.A(n_1009),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_963),
.A2(n_216),
.B(n_217),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_961),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_962),
.B(n_218),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_925),
.Y(n_1109)
);

AO21x2_ASAP7_75t_L g1110 ( 
.A1(n_870),
.A2(n_219),
.B(n_221),
.Y(n_1110)
);

OAI21x1_ASAP7_75t_L g1111 ( 
.A1(n_960),
.A2(n_223),
.B(n_225),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_972),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_911),
.B(n_226),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_975),
.Y(n_1114)
);

BUFx4_ASAP7_75t_SL g1115 ( 
.A(n_1011),
.Y(n_1115)
);

BUFx3_ASAP7_75t_L g1116 ( 
.A(n_925),
.Y(n_1116)
);

OA21x2_ASAP7_75t_L g1117 ( 
.A1(n_934),
.A2(n_229),
.B(n_233),
.Y(n_1117)
);

INVx6_ASAP7_75t_SL g1118 ( 
.A(n_935),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_945),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_951),
.B(n_234),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_951),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_981),
.Y(n_1122)
);

NAND2x1_ASAP7_75t_L g1123 ( 
.A(n_951),
.B(n_235),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_993),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_917),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_878),
.B(n_237),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_994),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_886),
.A2(n_239),
.B(n_240),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_893),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1004),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_936),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_909),
.Y(n_1132)
);

AOI22x1_ASAP7_75t_L g1133 ( 
.A1(n_889),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_892),
.B(n_939),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_895),
.A2(n_249),
.B(n_251),
.Y(n_1135)
);

AOI22x1_ASAP7_75t_L g1136 ( 
.A1(n_1002),
.A2(n_252),
.B1(n_254),
.B2(n_257),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_976),
.B(n_258),
.Y(n_1137)
);

AOI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_896),
.A2(n_259),
.B1(n_260),
.B2(n_263),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1014),
.Y(n_1139)
);

NAND2x1p5_ASAP7_75t_L g1140 ( 
.A(n_903),
.B(n_264),
.Y(n_1140)
);

BUFx2_ASAP7_75t_SL g1141 ( 
.A(n_871),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_879),
.A2(n_938),
.B(n_970),
.Y(n_1142)
);

HB1xp67_ASAP7_75t_L g1143 ( 
.A(n_947),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_882),
.A2(n_268),
.B(n_269),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_887),
.A2(n_274),
.B(n_276),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_872),
.A2(n_277),
.B(n_279),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_937),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_1013),
.A2(n_281),
.B(n_282),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_955),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_874),
.B(n_284),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1005),
.A2(n_285),
.B(n_286),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_949),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_921),
.A2(n_287),
.B(n_288),
.Y(n_1153)
);

INVx8_ASAP7_75t_L g1154 ( 
.A(n_885),
.Y(n_1154)
);

AO21x2_ASAP7_75t_L g1155 ( 
.A1(n_899),
.A2(n_289),
.B(n_290),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_907),
.A2(n_293),
.B(n_295),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_932),
.B(n_297),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_971),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1018),
.Y(n_1159)
);

OAI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1102),
.A2(n_973),
.B1(n_1008),
.B2(n_997),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1060),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1038),
.Y(n_1162)
);

BUFx4f_ASAP7_75t_SL g1163 ( 
.A(n_1041),
.Y(n_1163)
);

AO21x2_ASAP7_75t_L g1164 ( 
.A1(n_1050),
.A2(n_1015),
.B(n_995),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1063),
.A2(n_1067),
.B1(n_1149),
.B2(n_1143),
.Y(n_1165)
);

AO21x2_ASAP7_75t_L g1166 ( 
.A1(n_1050),
.A2(n_985),
.B(n_890),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1118),
.A2(n_890),
.B1(n_301),
.B2(n_303),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1049),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1083),
.B(n_414),
.Y(n_1169)
);

NAND2x1p5_ASAP7_75t_L g1170 ( 
.A(n_1033),
.B(n_298),
.Y(n_1170)
);

BUFx4f_ASAP7_75t_SL g1171 ( 
.A(n_1041),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1028),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1080),
.B(n_413),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1057),
.B(n_308),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1118),
.A2(n_311),
.B1(n_316),
.B2(n_318),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1029),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1029),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_SL g1178 ( 
.A(n_1059),
.B(n_319),
.C(n_320),
.Y(n_1178)
);

CKINVDCx11_ASAP7_75t_R g1179 ( 
.A(n_1074),
.Y(n_1179)
);

OA21x2_ASAP7_75t_L g1180 ( 
.A1(n_1101),
.A2(n_321),
.B(n_323),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_1090),
.B(n_324),
.Y(n_1181)
);

INVxp33_ASAP7_75t_L g1182 ( 
.A(n_1021),
.Y(n_1182)
);

AOI22xp33_ASAP7_75t_SL g1183 ( 
.A1(n_1092),
.A2(n_325),
.B1(n_328),
.B2(n_329),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1070),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1053),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1149),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1113),
.A2(n_333),
.B1(n_335),
.B2(n_336),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1045),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1056),
.B(n_338),
.Y(n_1189)
);

NAND2x1p5_ASAP7_75t_L g1190 ( 
.A(n_1033),
.B(n_341),
.Y(n_1190)
);

AOI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1094),
.A2(n_342),
.B(n_343),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1058),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_1085),
.Y(n_1193)
);

AOI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1094),
.A2(n_345),
.B(n_346),
.Y(n_1194)
);

AOI222xp33_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_347),
.B1(n_349),
.B2(n_350),
.C1(n_352),
.C2(n_353),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1115),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1095),
.A2(n_354),
.B(n_357),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_SL g1198 ( 
.A1(n_1061),
.A2(n_358),
.B(n_361),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1035),
.B(n_411),
.Y(n_1199)
);

INVx4_ASAP7_75t_L g1200 ( 
.A(n_1104),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1142),
.A2(n_362),
.B(n_364),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1107),
.B(n_365),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1107),
.B(n_410),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1026),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1089),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1065),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1073),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1152),
.A2(n_366),
.B1(n_367),
.B2(n_369),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1129),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1025),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1150),
.A2(n_370),
.B1(n_372),
.B2(n_374),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_SL g1212 ( 
.A1(n_1150),
.A2(n_1125),
.B1(n_1035),
.B2(n_1069),
.Y(n_1212)
);

AOI22xp5_ASAP7_75t_L g1213 ( 
.A1(n_1132),
.A2(n_1055),
.B1(n_1105),
.B2(n_1141),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1109),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1079),
.Y(n_1215)
);

AO22x1_ASAP7_75t_L g1216 ( 
.A1(n_1157),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1036),
.A2(n_378),
.B(n_379),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1100),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1141),
.A2(n_380),
.B1(n_381),
.B2(n_386),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1147),
.A2(n_387),
.B1(n_388),
.B2(n_391),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1134),
.B(n_392),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1019),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_1222)
);

AOI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1097),
.A2(n_397),
.B(n_398),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1084),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1096),
.B(n_408),
.Y(n_1225)
);

BUFx12f_ASAP7_75t_L g1226 ( 
.A(n_1040),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1086),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1086),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1131),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1077),
.Y(n_1230)
);

CKINVDCx11_ASAP7_75t_R g1231 ( 
.A(n_1030),
.Y(n_1231)
);

INVx4_ASAP7_75t_SL g1232 ( 
.A(n_1088),
.Y(n_1232)
);

AOI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_1158),
.A2(n_407),
.B(n_405),
.Y(n_1233)
);

AO21x1_ASAP7_75t_SL g1234 ( 
.A1(n_1156),
.A2(n_406),
.B(n_1093),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1112),
.Y(n_1235)
);

AOI21xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1154),
.A2(n_1157),
.B(n_1042),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1046),
.B(n_1047),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1114),
.A2(n_1130),
.B1(n_1139),
.B2(n_1127),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1116),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1088),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1122),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1147),
.A2(n_1114),
.B1(n_1139),
.B2(n_1127),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1089),
.B(n_1119),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1025),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1025),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1044),
.Y(n_1246)
);

CKINVDCx20_ASAP7_75t_R g1247 ( 
.A(n_1047),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_1081),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1025),
.Y(n_1249)
);

BUFx2_ASAP7_75t_SL g1250 ( 
.A(n_1064),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1124),
.Y(n_1251)
);

BUFx2_ASAP7_75t_SL g1252 ( 
.A(n_1064),
.Y(n_1252)
);

INVx8_ASAP7_75t_L g1253 ( 
.A(n_1154),
.Y(n_1253)
);

CKINVDCx6p67_ASAP7_75t_R g1254 ( 
.A(n_1046),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1130),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1020),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1037),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1103),
.B(n_1037),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1103),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1017),
.A2(n_1031),
.B(n_1032),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1108),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1048),
.A2(n_1027),
.B1(n_1136),
.B2(n_1138),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1020),
.Y(n_1263)
);

BUFx10_ASAP7_75t_L g1264 ( 
.A(n_1081),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1137),
.A2(n_1148),
.B1(n_1135),
.B2(n_1072),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1120),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1022),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_1262),
.A2(n_1128),
.A3(n_1024),
.B(n_1068),
.Y(n_1268)
);

HB1xp67_ASAP7_75t_L g1269 ( 
.A(n_1172),
.Y(n_1269)
);

CKINVDCx9p33_ASAP7_75t_R g1270 ( 
.A(n_1218),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1247),
.B(n_1052),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1168),
.Y(n_1272)
);

CKINVDCx14_ASAP7_75t_R g1273 ( 
.A(n_1179),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1253),
.Y(n_1274)
);

NOR3xp33_ASAP7_75t_SL g1275 ( 
.A(n_1196),
.B(n_1160),
.C(n_1165),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1174),
.A2(n_1072),
.B1(n_1075),
.B2(n_1133),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1212),
.B(n_1213),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1221),
.A2(n_1133),
.B1(n_1023),
.B2(n_1120),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1162),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_R g1280 ( 
.A(n_1189),
.B(n_1062),
.Y(n_1280)
);

INVx4_ASAP7_75t_SL g1281 ( 
.A(n_1163),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1254),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1214),
.B(n_1052),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1176),
.B(n_1087),
.Y(n_1284)
);

CKINVDCx16_ASAP7_75t_R g1285 ( 
.A(n_1230),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1177),
.Y(n_1286)
);

AND2x4_ASAP7_75t_SL g1287 ( 
.A(n_1193),
.B(n_1121),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1209),
.Y(n_1288)
);

OR2x6_ASAP7_75t_L g1289 ( 
.A(n_1250),
.B(n_1043),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1198),
.A2(n_1076),
.B(n_1144),
.Y(n_1290)
);

AOI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1189),
.A2(n_1054),
.B1(n_1091),
.B2(n_1078),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1195),
.A2(n_1140),
.B(n_1126),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_R g1293 ( 
.A(n_1199),
.B(n_1071),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_1240),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1188),
.B(n_1082),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1159),
.Y(n_1296)
);

NAND2xp33_ASAP7_75t_SL g1297 ( 
.A(n_1237),
.B(n_1123),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1239),
.B(n_1153),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1181),
.B(n_1145),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1161),
.B(n_1151),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1169),
.B(n_1199),
.Y(n_1301)
);

AND2x2_ASAP7_75t_SL g1302 ( 
.A(n_1266),
.B(n_1071),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1192),
.B(n_1155),
.Y(n_1303)
);

NAND2xp33_ASAP7_75t_R g1304 ( 
.A(n_1236),
.B(n_1117),
.Y(n_1304)
);

BUFx3_ASAP7_75t_L g1305 ( 
.A(n_1171),
.Y(n_1305)
);

CKINVDCx16_ASAP7_75t_R g1306 ( 
.A(n_1204),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1207),
.Y(n_1307)
);

NAND2xp33_ASAP7_75t_R g1308 ( 
.A(n_1243),
.B(n_1173),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1246),
.Y(n_1309)
);

OR2x6_ASAP7_75t_L g1310 ( 
.A(n_1252),
.B(n_1111),
.Y(n_1310)
);

NOR2x1_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_1099),
.Y(n_1311)
);

AO31x2_ASAP7_75t_L g1312 ( 
.A1(n_1267),
.A2(n_1110),
.A3(n_1098),
.B(n_1146),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1258),
.B(n_1106),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1227),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1206),
.B(n_1228),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1235),
.B(n_1051),
.Y(n_1316)
);

NOR3xp33_ASAP7_75t_SL g1317 ( 
.A(n_1238),
.B(n_1066),
.C(n_1039),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1231),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1185),
.A2(n_1164),
.B1(n_1224),
.B2(n_1215),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1259),
.B(n_1255),
.Y(n_1320)
);

NAND3xp33_ASAP7_75t_SL g1321 ( 
.A(n_1211),
.B(n_1184),
.C(n_1261),
.Y(n_1321)
);

NAND4xp25_ASAP7_75t_L g1322 ( 
.A(n_1241),
.B(n_1251),
.C(n_1242),
.D(n_1167),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1232),
.B(n_1182),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1257),
.B(n_1205),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1226),
.Y(n_1325)
);

OAI21xp33_ASAP7_75t_SL g1326 ( 
.A1(n_1265),
.A2(n_1219),
.B(n_1244),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1232),
.B(n_1200),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1248),
.B(n_1203),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1248),
.B(n_1202),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_SL g1330 ( 
.A(n_1200),
.B(n_1253),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1256),
.Y(n_1331)
);

OR2x6_ASAP7_75t_L g1332 ( 
.A(n_1170),
.B(n_1190),
.Y(n_1332)
);

INVxp67_ASAP7_75t_L g1333 ( 
.A(n_1264),
.Y(n_1333)
);

AND2x4_ASAP7_75t_SL g1334 ( 
.A(n_1264),
.B(n_1245),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1164),
.A2(n_1178),
.B1(n_1234),
.B2(n_1180),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1279),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1269),
.B(n_1249),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1272),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1286),
.B(n_1166),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1331),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1275),
.A2(n_1183),
.B1(n_1187),
.B2(n_1175),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1287),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1284),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1307),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1315),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1314),
.B(n_1303),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1298),
.B(n_1300),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1290),
.A2(n_1180),
.B(n_1201),
.Y(n_1348)
);

HB1xp67_ASAP7_75t_L g1349 ( 
.A(n_1320),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1299),
.B(n_1166),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1319),
.B(n_1263),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1283),
.B(n_1263),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1270),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1321),
.A2(n_1222),
.B1(n_1186),
.B2(n_1208),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1313),
.B(n_1210),
.Y(n_1355)
);

INVx2_ASAP7_75t_L g1356 ( 
.A(n_1316),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1277),
.A2(n_1220),
.B1(n_1229),
.B2(n_1233),
.Y(n_1357)
);

INVx2_ASAP7_75t_SL g1358 ( 
.A(n_1334),
.Y(n_1358)
);

BUFx12f_ASAP7_75t_L g1359 ( 
.A(n_1325),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1328),
.B(n_1329),
.Y(n_1360)
);

OAI22xp5_ASAP7_75t_L g1361 ( 
.A1(n_1276),
.A2(n_1197),
.B1(n_1191),
.B2(n_1194),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1322),
.B(n_1216),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1301),
.B(n_1217),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1297),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1332),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1302),
.B(n_1223),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1295),
.B(n_1260),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1344),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1340),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1342),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1340),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1344),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1347),
.B(n_1335),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1352),
.B(n_1324),
.Y(n_1374)
);

OR2x2_ASAP7_75t_L g1375 ( 
.A(n_1345),
.B(n_1285),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1362),
.B(n_1280),
.C(n_1292),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1360),
.B(n_1296),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1347),
.B(n_1268),
.Y(n_1378)
);

INVx3_ASAP7_75t_L g1379 ( 
.A(n_1364),
.Y(n_1379)
);

OAI221xp5_ASAP7_75t_L g1380 ( 
.A1(n_1362),
.A2(n_1278),
.B1(n_1326),
.B2(n_1291),
.C(n_1293),
.Y(n_1380)
);

INVx3_ASAP7_75t_L g1381 ( 
.A(n_1364),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1350),
.B(n_1268),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1350),
.B(n_1317),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1355),
.B(n_1310),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1355),
.B(n_1310),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1336),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1346),
.B(n_1312),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1339),
.B(n_1311),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1383),
.B(n_1339),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1383),
.B(n_1367),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1377),
.B(n_1337),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1373),
.B(n_1367),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1376),
.B(n_1365),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1375),
.B(n_1356),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1378),
.B(n_1384),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1385),
.B(n_1379),
.Y(n_1397)
);

INVx4_ASAP7_75t_L g1398 ( 
.A(n_1370),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1375),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1368),
.B(n_1338),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1372),
.B(n_1343),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1369),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1386),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1385),
.B(n_1366),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_1369),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1381),
.B(n_1374),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1394),
.A2(n_1380),
.B1(n_1341),
.B2(n_1308),
.Y(n_1407)
);

AOI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1399),
.A2(n_1354),
.B1(n_1357),
.B2(n_1365),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1390),
.B(n_1382),
.Y(n_1409)
);

OR2x2_ASAP7_75t_L g1410 ( 
.A(n_1395),
.B(n_1393),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1393),
.B(n_1382),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1405),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_SL g1413 ( 
.A(n_1398),
.B(n_1381),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1406),
.B(n_1397),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1403),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1389),
.B(n_1381),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1403),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1404),
.A2(n_1387),
.B1(n_1388),
.B2(n_1363),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1389),
.B(n_1371),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1402),
.Y(n_1420)
);

AOI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1392),
.A2(n_1365),
.B1(n_1271),
.B2(n_1351),
.Y(n_1421)
);

AOI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1407),
.A2(n_1408),
.B1(n_1421),
.B2(n_1387),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1415),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1420),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1412),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1419),
.B(n_1391),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1408),
.A2(n_1348),
.B(n_1391),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1417),
.Y(n_1428)
);

OAI31xp33_ASAP7_75t_L g1429 ( 
.A1(n_1411),
.A2(n_1404),
.A3(n_1366),
.B(n_1396),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1425),
.B(n_1273),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1424),
.Y(n_1431)
);

NAND2x1p5_ASAP7_75t_L g1432 ( 
.A(n_1422),
.B(n_1398),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1426),
.Y(n_1433)
);

OAI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1422),
.A2(n_1421),
.B1(n_1418),
.B2(n_1409),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1434),
.A2(n_1427),
.B(n_1429),
.Y(n_1435)
);

INVx1_ASAP7_75t_SL g1436 ( 
.A(n_1430),
.Y(n_1436)
);

NOR3xp33_ASAP7_75t_L g1437 ( 
.A(n_1431),
.B(n_1306),
.C(n_1294),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1433),
.B(n_1318),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1432),
.B(n_1398),
.C(n_1401),
.Y(n_1439)
);

OAI21xp33_ASAP7_75t_L g1440 ( 
.A1(n_1433),
.A2(n_1416),
.B(n_1413),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1435),
.A2(n_1428),
.B1(n_1423),
.B2(n_1388),
.Y(n_1441)
);

NOR3xp33_ASAP7_75t_L g1442 ( 
.A(n_1437),
.B(n_1274),
.C(n_1327),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1436),
.A2(n_1353),
.B(n_1305),
.C(n_1361),
.Y(n_1443)
);

OAI31xp33_ASAP7_75t_L g1444 ( 
.A1(n_1441),
.A2(n_1439),
.A3(n_1438),
.B(n_1440),
.Y(n_1444)
);

OAI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1443),
.A2(n_1288),
.B1(n_1370),
.B2(n_1304),
.C(n_1332),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1445),
.B(n_1359),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1446),
.B(n_1444),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1447),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1447),
.Y(n_1449)
);

XOR2xp5_ASAP7_75t_L g1450 ( 
.A(n_1448),
.B(n_1282),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1449),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1451),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1450),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1452),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1453),
.Y(n_1455)
);

XNOR2xp5_ASAP7_75t_L g1456 ( 
.A(n_1453),
.B(n_1442),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1454),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1455),
.A2(n_1359),
.B1(n_1281),
.B2(n_1309),
.Y(n_1458)
);

OAI22x1_ASAP7_75t_L g1459 ( 
.A1(n_1456),
.A2(n_1281),
.B1(n_1330),
.B2(n_1333),
.Y(n_1459)
);

INVx3_ASAP7_75t_L g1460 ( 
.A(n_1454),
.Y(n_1460)
);

OAI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1457),
.A2(n_1289),
.B(n_1323),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1458),
.A2(n_1282),
.B(n_1309),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_1460),
.Y(n_1463)
);

NOR2x1_ASAP7_75t_R g1464 ( 
.A(n_1459),
.B(n_1342),
.Y(n_1464)
);

OAI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1460),
.A2(n_1289),
.B1(n_1358),
.B2(n_1410),
.Y(n_1465)
);

OAI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1463),
.A2(n_1414),
.B1(n_1358),
.B2(n_1400),
.Y(n_1466)
);

OR2x6_ASAP7_75t_L g1467 ( 
.A(n_1466),
.B(n_1462),
.Y(n_1467)
);

AOI211xp5_ASAP7_75t_L g1468 ( 
.A1(n_1467),
.A2(n_1464),
.B(n_1461),
.C(n_1465),
.Y(n_1468)
);


endmodule