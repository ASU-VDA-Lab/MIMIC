module fake_netlist_1_1585_n_673 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_673);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_673;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_522;
wire n_264;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_25), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_45), .Y(n_78) );
BUFx6f_ASAP7_75t_L g79 ( .A(n_46), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_14), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_29), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_22), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_37), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_36), .Y(n_84) );
INVxp67_ASAP7_75t_L g85 ( .A(n_30), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_15), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_39), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_62), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_53), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_52), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_73), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_48), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_21), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_31), .Y(n_94) );
INVx1_ASAP7_75t_SL g95 ( .A(n_0), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_65), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_60), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_33), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_15), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_20), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_70), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_2), .Y(n_102) );
INVxp67_ASAP7_75t_SL g103 ( .A(n_34), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_69), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_57), .B(n_0), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_32), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_9), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_9), .Y(n_109) );
INVxp33_ASAP7_75t_SL g110 ( .A(n_50), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_59), .Y(n_111) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_19), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_61), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_17), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_55), .Y(n_115) );
NOR2xp67_ASAP7_75t_L g116 ( .A(n_58), .B(n_23), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_1), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_44), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_75), .Y(n_119) );
INVx3_ASAP7_75t_L g120 ( .A(n_43), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_47), .Y(n_121) );
CKINVDCx16_ASAP7_75t_R g122 ( .A(n_14), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_27), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_122), .B(n_1), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_104), .B(n_3), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_77), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_120), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_77), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_120), .B(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_78), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_92), .B(n_4), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_88), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_91), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_79), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_80), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_79), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_97), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_123), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_79), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_112), .B(n_4), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_100), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_80), .A2(n_107), .B1(n_109), .B2(n_108), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_101), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_83), .B(n_5), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
XOR2xp5_ASAP7_75t_L g154 ( .A(n_98), .B(n_5), .Y(n_154) );
AND2x4_ASAP7_75t_L g155 ( .A(n_86), .B(n_6), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_87), .B(n_6), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_101), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_123), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_86), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_113), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_87), .B(n_7), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_93), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_121), .B(n_7), .Y(n_164) );
BUFx8_ASAP7_75t_L g165 ( .A(n_93), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_115), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_127), .B(n_90), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_141), .A2(n_102), .B1(n_99), .B2(n_107), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_127), .B(n_94), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_127), .B(n_84), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_127), .B(n_114), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_129), .A2(n_106), .B(n_103), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_126), .B(n_85), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_160), .B(n_108), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_126), .B(n_111), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_128), .B(n_110), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_128), .B(n_82), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_165), .B(n_121), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_129), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_130), .B(n_96), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_165), .B(n_119), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_130), .B(n_96), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_132), .B(n_89), .Y(n_185) );
AO221x1_ASAP7_75t_L g186 ( .A1(n_150), .A2(n_119), .B1(n_118), .B2(n_115), .C(n_117), .Y(n_186) );
NOR3xp33_ASAP7_75t_L g187 ( .A(n_124), .B(n_95), .C(n_117), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_155), .A2(n_114), .B1(n_109), .B2(n_99), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_155), .A2(n_102), .B1(n_118), .B2(n_89), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_125), .A2(n_81), .B1(n_105), .B2(n_116), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_165), .B(n_41), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_165), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_135), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_132), .B(n_8), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_125), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_134), .B(n_42), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_155), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_134), .B(n_10), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_136), .B(n_11), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_136), .B(n_12), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_137), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_155), .B(n_12), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_138), .B(n_13), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_138), .B(n_13), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_137), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_139), .B(n_16), .Y(n_208) );
NAND2xp33_ASAP7_75t_L g209 ( .A(n_139), .B(n_54), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_133), .A2(n_16), .B1(n_17), .B2(n_18), .Y(n_210) );
NAND2xp33_ASAP7_75t_L g211 ( .A(n_143), .B(n_56), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_143), .B(n_18), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_133), .A2(n_24), .B1(n_26), .B2(n_28), .Y(n_214) );
NOR3xp33_ASAP7_75t_L g215 ( .A(n_147), .B(n_35), .C(n_38), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_146), .B(n_40), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_146), .B(n_49), .Y(n_219) );
AOI22xp5_ASAP7_75t_L g220 ( .A1(n_147), .A2(n_51), .B1(n_63), .B2(n_64), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_148), .B(n_66), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_192), .B(n_131), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_204), .Y(n_223) );
AO21x1_ASAP7_75t_L g224 ( .A1(n_209), .A2(n_162), .B(n_156), .Y(n_224) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_173), .A2(n_149), .B(n_161), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_177), .B(n_196), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_192), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_204), .B(n_149), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_181), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_196), .B(n_151), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_212), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_176), .B(n_151), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_168), .Y(n_234) );
OR2x6_ASAP7_75t_L g235 ( .A(n_204), .B(n_166), .Y(n_235) );
HB1xp67_ASAP7_75t_L g236 ( .A(n_175), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_188), .B(n_148), .Y(n_237) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_170), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_175), .B(n_166), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_172), .Y(n_241) );
OR2x6_ASAP7_75t_L g242 ( .A(n_198), .B(n_157), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_170), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_178), .B(n_158), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_180), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_174), .B(n_158), .Y(n_246) );
NOR2xp33_ASAP7_75t_R g247 ( .A(n_209), .B(n_159), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_179), .B(n_157), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_172), .B(n_161), .Y(n_249) );
HB1xp67_ASAP7_75t_L g250 ( .A(n_172), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_189), .B(n_144), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_167), .Y(n_252) );
INVxp67_ASAP7_75t_L g253 ( .A(n_169), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_190), .B(n_152), .Y(n_254) );
BUFx12f_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
BUFx2_ASAP7_75t_L g256 ( .A(n_171), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_180), .Y(n_257) );
AO22x1_ASAP7_75t_L g258 ( .A1(n_215), .A2(n_159), .B1(n_144), .B2(n_164), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_182), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_195), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_183), .B(n_159), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_187), .B(n_159), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_199), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_193), .Y(n_264) );
INVxp67_ASAP7_75t_SL g265 ( .A(n_184), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_185), .B(n_153), .Y(n_266) );
BUFx12f_ASAP7_75t_L g267 ( .A(n_186), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_201), .A2(n_163), .B(n_153), .C(n_145), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_205), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_214), .B(n_163), .Y(n_271) );
AND3x1_ASAP7_75t_L g272 ( .A(n_210), .B(n_154), .C(n_163), .Y(n_272) );
INVx3_ASAP7_75t_L g273 ( .A(n_206), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_208), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_213), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_193), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_218), .B(n_145), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_194), .Y(n_278) );
BUFx2_ASAP7_75t_L g279 ( .A(n_214), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_219), .B(n_145), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_194), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_220), .B(n_140), .Y(n_283) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_236), .A2(n_191), .B(n_221), .C(n_211), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_235), .B(n_220), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_235), .A2(n_223), .B1(n_279), .B2(n_271), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_238), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_262), .A2(n_197), .B(n_211), .C(n_142), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_235), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_239), .B(n_154), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_279), .A2(n_217), .B1(n_216), .B2(n_207), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_235), .A2(n_217), .B(n_216), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_248), .A2(n_142), .B(n_203), .C(n_200), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_238), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_229), .A2(n_207), .B(n_203), .Y(n_297) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_224), .B(n_140), .Y(n_298) );
AOI21xp5_ASAP7_75t_L g299 ( .A1(n_233), .A2(n_140), .B(n_68), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
BUFx3_ASAP7_75t_L g301 ( .A(n_257), .Y(n_301) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_224), .B(n_140), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_238), .Y(n_303) );
A2O1A1Ixp33_ASAP7_75t_SL g304 ( .A1(n_253), .A2(n_140), .B(n_71), .C(n_72), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_259), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_239), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_244), .A2(n_140), .B(n_74), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_234), .Y(n_308) );
AND2x4_ASAP7_75t_L g309 ( .A(n_239), .B(n_67), .Y(n_309) );
OR2x6_ASAP7_75t_L g310 ( .A(n_223), .B(n_76), .Y(n_310) );
NAND2xp33_ASAP7_75t_SL g311 ( .A(n_247), .B(n_257), .Y(n_311) );
BUFx3_ASAP7_75t_L g312 ( .A(n_238), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_243), .Y(n_313) );
BUFx12f_ASAP7_75t_L g314 ( .A(n_234), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_243), .Y(n_315) );
A2O1A1Ixp33_ASAP7_75t_SL g316 ( .A1(n_273), .A2(n_225), .B(n_274), .C(n_263), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_241), .A2(n_271), .B1(n_250), .B2(n_259), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_231), .B(n_260), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_222), .A2(n_261), .B(n_280), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_231), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_241), .Y(n_321) );
INVxp67_ASAP7_75t_SL g322 ( .A(n_243), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_271), .A2(n_249), .B1(n_242), .B2(n_269), .Y(n_323) );
BUFx6f_ASAP7_75t_SL g324 ( .A(n_242), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_252), .B(n_256), .Y(n_325) );
INVx2_ASAP7_75t_SL g326 ( .A(n_275), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_243), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_277), .A2(n_274), .B(n_269), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_254), .B(n_242), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_245), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_252), .B(n_256), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_242), .A2(n_263), .B1(n_270), .B2(n_227), .Y(n_332) );
CKINVDCx5p33_ASAP7_75t_R g333 ( .A(n_255), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_270), .B(n_273), .Y(n_334) );
INVxp33_ASAP7_75t_L g335 ( .A(n_325), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_312), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_328), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_285), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_334), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_334), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_286), .B(n_245), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_301), .Y(n_344) );
CKINVDCx6p67_ASAP7_75t_R g345 ( .A(n_301), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_312), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_290), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_286), .B(n_273), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_288), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_293), .Y(n_352) );
INVxp67_ASAP7_75t_L g353 ( .A(n_318), .Y(n_353) );
INVx1_ASAP7_75t_SL g354 ( .A(n_325), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_309), .Y(n_355) );
INVx3_ASAP7_75t_L g356 ( .A(n_313), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_320), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_293), .Y(n_358) );
OAI21xp5_ASAP7_75t_L g359 ( .A1(n_298), .A2(n_232), .B(n_283), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_321), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_296), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_298), .A2(n_251), .B(n_266), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_286), .B(n_246), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_302), .A2(n_232), .B(n_268), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
AOI21xp33_ASAP7_75t_SL g366 ( .A1(n_333), .A2(n_258), .B(n_272), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_363), .B(n_323), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_363), .B(n_287), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g369 ( .A(n_345), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_363), .B(n_331), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_343), .B(n_329), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_355), .A2(n_324), .B1(n_267), .B2(n_255), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_340), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_349), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_340), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_343), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_345), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_343), .B(n_355), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_355), .B(n_309), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_353), .B(n_317), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_349), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_348), .B(n_309), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_360), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_354), .B(n_306), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_354), .B(n_353), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_336), .Y(n_389) );
INVxp67_ASAP7_75t_SL g390 ( .A(n_344), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_348), .B(n_310), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_365), .A2(n_310), .B1(n_324), .B2(n_292), .Y(n_392) );
INVx3_ASAP7_75t_SL g393 ( .A(n_345), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_348), .A2(n_267), .B1(n_314), .B2(n_308), .Y(n_394) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_392), .A2(n_308), .B1(n_347), .B2(n_344), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_370), .B(n_368), .Y(n_396) );
INVx1_ASAP7_75t_SL g397 ( .A(n_393), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_368), .B(n_335), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_374), .Y(n_399) );
NAND4xp25_ASAP7_75t_L g400 ( .A(n_394), .B(n_366), .C(n_291), .D(n_357), .Y(n_400) );
INVxp33_ASAP7_75t_L g401 ( .A(n_388), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_370), .B(n_357), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_374), .Y(n_403) );
NAND3xp33_ASAP7_75t_L g404 ( .A(n_392), .B(n_366), .C(n_302), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_393), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_372), .B(n_344), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_367), .B(n_338), .Y(n_407) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_390), .Y(n_408) );
AO21x2_ASAP7_75t_L g409 ( .A1(n_371), .A2(n_365), .B(n_359), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_388), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_372), .B(n_338), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_378), .B(n_341), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_376), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_393), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_326), .B1(n_335), .B2(n_350), .C(n_351), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
NAND3xp33_ASAP7_75t_L g418 ( .A(n_373), .B(n_258), .C(n_316), .Y(n_418) );
AOI21x1_ASAP7_75t_L g419 ( .A1(n_371), .A2(n_359), .B(n_364), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_377), .Y(n_420) );
INVx4_ASAP7_75t_SL g421 ( .A(n_379), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_372), .B(n_350), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_381), .A2(n_310), .B1(n_347), .B2(n_342), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_391), .A2(n_314), .B1(n_311), .B2(n_347), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_381), .A2(n_342), .B1(n_341), .B2(n_351), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_367), .B(n_364), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_427), .B(n_371), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_410), .B(n_390), .Y(n_430) );
OA21x2_ASAP7_75t_L g431 ( .A1(n_404), .A2(n_375), .B(n_419), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_427), .B(n_367), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_406), .B(n_375), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_406), .B(n_375), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_407), .B(n_368), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx1_ASAP7_75t_SL g437 ( .A(n_397), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_408), .Y(n_439) );
NOR2x1p5_ASAP7_75t_L g440 ( .A(n_418), .B(n_379), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_413), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_407), .B(n_386), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_413), .B(n_383), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_415), .Y(n_444) );
NAND3xp33_ASAP7_75t_L g445 ( .A(n_400), .B(n_316), .C(n_386), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g446 ( .A(n_395), .B(n_379), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_415), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g448 ( .A(n_405), .B(n_369), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_402), .B(n_385), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_421), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_426), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_417), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_411), .B(n_385), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_409), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_409), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_409), .Y(n_457) );
AOI32xp33_ASAP7_75t_L g458 ( .A1(n_423), .A2(n_391), .A3(n_381), .B1(n_311), .B2(n_384), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_396), .B(n_383), .Y(n_459) );
NAND2x1p5_ASAP7_75t_L g460 ( .A(n_414), .B(n_389), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_416), .A2(n_383), .B(n_304), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_401), .B(n_380), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_411), .B(n_378), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_398), .B(n_401), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_412), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_398), .B(n_380), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_422), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_425), .B(n_380), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_421), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_424), .B(n_391), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_432), .B(n_389), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVxp67_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
OAI31xp33_ASAP7_75t_L g478 ( .A1(n_446), .A2(n_382), .A3(n_384), .B(n_305), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_448), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_432), .B(n_429), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_469), .B(n_382), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_469), .B(n_384), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_429), .B(n_387), .Y(n_484) );
NAND2xp33_ASAP7_75t_L g485 ( .A(n_458), .B(n_389), .Y(n_485) );
INVx1_ASAP7_75t_SL g486 ( .A(n_433), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_429), .B(n_389), .Y(n_487) );
NAND2xp33_ASAP7_75t_L g488 ( .A(n_458), .B(n_389), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_473), .B(n_387), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_465), .B(n_387), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_429), .B(n_389), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
HB1xp67_ASAP7_75t_L g493 ( .A(n_452), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_436), .B(n_389), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_470), .B(n_362), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_470), .B(n_362), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_436), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_438), .B(n_362), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_438), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_444), .Y(n_500) );
CKINVDCx16_ASAP7_75t_R g501 ( .A(n_450), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_442), .B(n_295), .Y(n_502) );
AND2x4_ASAP7_75t_SL g503 ( .A(n_450), .B(n_346), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_462), .B(n_295), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_451), .B(n_361), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_472), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_451), .B(n_361), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_433), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_464), .B(n_300), .Y(n_509) );
INVxp67_ASAP7_75t_L g510 ( .A(n_430), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_454), .B(n_237), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_434), .B(n_361), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_430), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_444), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_434), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_462), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_468), .B(n_289), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_444), .B(n_361), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_468), .B(n_289), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_459), .B(n_435), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_447), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_459), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_463), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_449), .B(n_358), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_471), .B(n_358), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_474), .A2(n_336), .B1(n_346), .B2(n_356), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_471), .B(n_358), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_447), .B(n_358), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_463), .Y(n_529) );
AOI211xp5_ASAP7_75t_L g530 ( .A1(n_474), .A2(n_284), .B(n_299), .C(n_307), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_476), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_480), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_513), .B(n_466), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_492), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_497), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_510), .B(n_522), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_490), .A2(n_445), .B1(n_467), .B2(n_466), .C(n_456), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_516), .B(n_467), .Y(n_538) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_476), .B(n_440), .Y(n_539) );
NAND2xp33_ASAP7_75t_L g540 ( .A(n_489), .B(n_440), .Y(n_540) );
NAND4xp25_ASAP7_75t_L g541 ( .A(n_478), .B(n_445), .C(n_473), .D(n_461), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_486), .B(n_443), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_481), .B(n_456), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_508), .B(n_443), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_493), .B(n_453), .Y(n_545) );
NAND2xp33_ASAP7_75t_SL g546 ( .A(n_501), .B(n_472), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_479), .B(n_472), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_520), .B(n_447), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_481), .B(n_460), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_475), .B(n_460), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_485), .A2(n_488), .B1(n_477), .B2(n_509), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_500), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_515), .B(n_453), .Y(n_553) );
INVxp33_ASAP7_75t_L g554 ( .A(n_512), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_475), .B(n_431), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_487), .B(n_460), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_487), .B(n_431), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_499), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_494), .B(n_431), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_529), .B(n_453), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_505), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_500), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_517), .B(n_441), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_505), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_507), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_507), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_484), .B(n_441), .Y(n_568) );
AND2x4_ASAP7_75t_L g569 ( .A(n_506), .B(n_457), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_519), .B(n_482), .Y(n_570) );
NOR2xp33_ASAP7_75t_R g571 ( .A(n_485), .B(n_336), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_514), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_484), .B(n_431), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_511), .B(n_457), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_506), .B(n_455), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_494), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_504), .B(n_455), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_503), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_514), .Y(n_581) );
NAND3xp33_ASAP7_75t_L g582 ( .A(n_537), .B(n_488), .C(n_530), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_552), .Y(n_583) );
NAND3xp33_ASAP7_75t_L g584 ( .A(n_531), .B(n_506), .C(n_498), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_570), .A2(n_502), .B1(n_483), .B2(n_525), .C(n_527), .Y(n_585) );
AOI322xp5_ASAP7_75t_L g586 ( .A1(n_546), .A2(n_526), .A3(n_498), .B1(n_495), .B2(n_496), .C1(n_521), .C2(n_528), .Y(n_586) );
AOI21xp5_ASAP7_75t_L g587 ( .A1(n_540), .A2(n_503), .B(n_518), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_543), .B(n_521), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_552), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_543), .B(n_579), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_546), .B(n_518), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_532), .Y(n_592) );
AND2x2_ASAP7_75t_SL g593 ( .A(n_540), .B(n_491), .Y(n_593) );
NAND3xp33_ASAP7_75t_L g594 ( .A(n_541), .B(n_491), .C(n_528), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_574), .A2(n_346), .B1(n_336), .B2(n_356), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_539), .A2(n_304), .B(n_346), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_574), .B(n_349), .Y(n_597) );
OAI21xp5_ASAP7_75t_SL g598 ( .A1(n_551), .A2(n_336), .B(n_346), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_534), .Y(n_599) );
NOR2xp67_ASAP7_75t_L g600 ( .A(n_557), .B(n_349), .Y(n_600) );
OAI21xp33_ASAP7_75t_L g601 ( .A1(n_536), .A2(n_356), .B(n_352), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_547), .B(n_356), .C(n_319), .Y(n_603) );
NAND3xp33_ASAP7_75t_SL g604 ( .A(n_571), .B(n_352), .C(n_337), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_577), .B(n_352), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_558), .Y(n_606) );
NOR2xp33_ASAP7_75t_SL g607 ( .A(n_580), .B(n_337), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_549), .B(n_337), .Y(n_608) );
OAI32xp33_ASAP7_75t_L g609 ( .A1(n_554), .A2(n_356), .A3(n_313), .B1(n_327), .B2(n_315), .Y(n_609) );
OAI211xp5_ASAP7_75t_SL g610 ( .A1(n_578), .A2(n_294), .B(n_297), .C(n_281), .Y(n_610) );
NOR4xp25_ASAP7_75t_L g611 ( .A(n_545), .B(n_313), .C(n_315), .D(n_327), .Y(n_611) );
O2A1O1Ixp33_ASAP7_75t_L g612 ( .A1(n_575), .A2(n_322), .B(n_303), .C(n_296), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_562), .B(n_243), .Y(n_613) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_571), .B(n_303), .Y(n_614) );
OAI211xp5_ASAP7_75t_SL g615 ( .A1(n_547), .A2(n_281), .B(n_278), .C(n_276), .Y(n_615) );
OAI31xp33_ASAP7_75t_L g616 ( .A1(n_554), .A2(n_228), .A3(n_278), .B(n_230), .Y(n_616) );
XNOR2x2_ASAP7_75t_L g617 ( .A(n_548), .B(n_226), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_560), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g619 ( .A1(n_582), .A2(n_538), .B1(n_533), .B2(n_573), .C(n_565), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_592), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_590), .B(n_555), .Y(n_621) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_598), .A2(n_564), .B1(n_553), .B2(n_544), .C(n_542), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_616), .A2(n_576), .B1(n_567), .B2(n_566), .C(n_555), .Y(n_623) );
AOI22xp33_ASAP7_75t_L g624 ( .A1(n_594), .A2(n_557), .B1(n_550), .B2(n_559), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_618), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_599), .Y(n_626) );
OR2x2_ASAP7_75t_L g627 ( .A(n_588), .B(n_559), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g628 ( .A(n_586), .B(n_576), .C(n_569), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_608), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_585), .A2(n_556), .B1(n_568), .B2(n_569), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_602), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_593), .A2(n_561), .B1(n_581), .B2(n_569), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g633 ( .A1(n_604), .A2(n_572), .B(n_563), .Y(n_633) );
AOI21xp5_ASAP7_75t_L g634 ( .A1(n_604), .A2(n_572), .B(n_563), .Y(n_634) );
NAND4xp75_ASAP7_75t_L g635 ( .A(n_591), .B(n_228), .C(n_226), .D(n_230), .Y(n_635) );
NOR2x1p5_ASAP7_75t_L g636 ( .A(n_584), .B(n_276), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_606), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_583), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_587), .A2(n_240), .B(n_264), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_589), .B(n_276), .Y(n_640) );
NOR3xp33_ASAP7_75t_L g641 ( .A(n_623), .B(n_615), .C(n_610), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_635), .B(n_615), .Y(n_642) );
NOR2x1_ASAP7_75t_L g643 ( .A(n_636), .B(n_614), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_628), .B(n_612), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_630), .A2(n_612), .B(n_597), .Y(n_645) );
NAND4xp75_ASAP7_75t_L g646 ( .A(n_619), .B(n_600), .C(n_596), .D(n_605), .Y(n_646) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_630), .A2(n_624), .B1(n_622), .B2(n_632), .Y(n_647) );
BUFx3_ASAP7_75t_L g648 ( .A(n_629), .Y(n_648) );
NOR2x1p5_ASAP7_75t_L g649 ( .A(n_621), .B(n_617), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_620), .Y(n_650) );
NAND3xp33_ASAP7_75t_SL g651 ( .A(n_624), .B(n_611), .C(n_607), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_625), .B(n_603), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_626), .Y(n_653) );
NOR3xp33_ASAP7_75t_L g654 ( .A(n_651), .B(n_640), .C(n_610), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_644), .B(n_652), .Y(n_655) );
INVx3_ASAP7_75t_L g656 ( .A(n_648), .Y(n_656) );
NAND4xp25_ASAP7_75t_L g657 ( .A(n_641), .B(n_595), .C(n_633), .D(n_634), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_647), .A2(n_637), .B1(n_631), .B2(n_638), .C(n_627), .Y(n_658) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_647), .A2(n_627), .B1(n_601), .B2(n_603), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_650), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_653), .B(n_613), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_656), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_658), .A2(n_645), .B1(n_649), .B2(n_646), .C(n_609), .Y(n_663) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_654), .B(n_642), .C(n_639), .D(n_643), .E(n_240), .Y(n_664) );
BUFx2_ASAP7_75t_L g665 ( .A(n_660), .Y(n_665) );
OR3x2_ASAP7_75t_L g666 ( .A(n_664), .B(n_662), .C(n_657), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_665), .B(n_655), .Y(n_667) );
XOR2xp5_ASAP7_75t_L g668 ( .A(n_663), .B(n_659), .Y(n_668) );
AO21x1_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_661), .B(n_264), .Y(n_669) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_667), .A2(n_282), .B(n_666), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_669), .Y(n_671) );
INVx1_ASAP7_75t_SL g672 ( .A(n_670), .Y(n_672) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_672), .A2(n_282), .B(n_671), .Y(n_673) );
endmodule