module fake_ariane_2737_n_200 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_200);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_200;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_190;
wire n_160;
wire n_64;
wire n_179;
wire n_180;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_195;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_197;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_187;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_199;
wire n_91;
wire n_159;
wire n_107;
wire n_189;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_94;
wire n_101;
wire n_48;
wire n_134;
wire n_188;
wire n_185;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_162;
wire n_45;
wire n_112;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_198;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_121;
wire n_93;
wire n_118;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_196;
wire n_125;
wire n_168;
wire n_81;
wire n_87;
wire n_43;
wire n_41;
wire n_140;
wire n_55;
wire n_191;
wire n_151;
wire n_136;
wire n_192;
wire n_80;
wire n_146;
wire n_194;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_186;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_193;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_21),
.Y(n_43)
);

INVxp67_ASAP7_75t_SL g44 ( 
.A(n_10),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp67_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_0),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_R g65 ( 
.A(n_52),
.B(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_R g72 ( 
.A(n_47),
.B(n_14),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_64),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2x1p5_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_55),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_55),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

CKINVDCx11_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

OR2x2_ASAP7_75t_SL g88 ( 
.A(n_62),
.B(n_45),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_54),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_70),
.B1(n_46),
.B2(n_45),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_75),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_75),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_73),
.B(n_69),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_60),
.B1(n_71),
.B2(n_69),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_71),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_90),
.Y(n_106)
);

OAI211xp5_ASAP7_75t_L g107 ( 
.A1(n_105),
.A2(n_44),
.B(n_89),
.C(n_76),
.Y(n_107)
);

AO21x2_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_72),
.B(n_53),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

OR2x4_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_93),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_87),
.C(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_74),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_98),
.B1(n_48),
.B2(n_90),
.Y(n_116)
);

AO31x2_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_97),
.A3(n_61),
.B(n_96),
.Y(n_117)
);

AO31x2_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_61),
.A3(n_96),
.B(n_95),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_88),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_115),
.A2(n_98),
.B1(n_106),
.B2(n_109),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_120),
.B(n_106),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g124 ( 
.A(n_116),
.B(n_84),
.Y(n_124)
);

OAI21x1_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_111),
.B(n_113),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_125),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_120),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_84),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_84),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_121),
.A2(n_86),
.B1(n_103),
.B2(n_108),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_117),
.Y(n_136)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_86),
.C(n_54),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_130),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_136),
.B(n_117),
.Y(n_142)
);

OAI21x1_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_91),
.B(n_80),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_140),
.B(n_134),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_135),
.B(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_142),
.B(n_132),
.Y(n_148)
);

OR2x6_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_131),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_132),
.B1(n_128),
.B2(n_131),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_53),
.A3(n_58),
.B1(n_136),
.B2(n_43),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_143),
.A2(n_58),
.A3(n_37),
.B1(n_36),
.B2(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_149),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_126),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_133),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_129),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_129),
.B1(n_146),
.B2(n_112),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_153),
.B(n_58),
.C(n_129),
.Y(n_165)
);

AOI211xp5_ASAP7_75t_SL g166 ( 
.A1(n_161),
.A2(n_133),
.B(n_82),
.C(n_99),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_155),
.A2(n_112),
.B(n_108),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_108),
.B1(n_91),
.B2(n_95),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_156),
.B(n_112),
.Y(n_169)
);

NAND3xp33_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_104),
.C(n_1),
.Y(n_170)
);

AOI221x1_ASAP7_75t_L g171 ( 
.A1(n_158),
.A2(n_104),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_171)
);

OAI211xp5_ASAP7_75t_L g172 ( 
.A1(n_171),
.A2(n_155),
.B(n_159),
.C(n_156),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_159),
.Y(n_173)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_0),
.Y(n_175)
);

OAI221xp5_ASAP7_75t_L g176 ( 
.A1(n_165),
.A2(n_104),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_176)
);

AOI221xp5_ASAP7_75t_L g177 ( 
.A1(n_167),
.A2(n_65),
.B1(n_7),
.B2(n_8),
.C(n_9),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_2),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g179 ( 
.A1(n_168),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_172),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_178),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_179),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_182),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

AOI21xp33_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_176),
.B(n_168),
.Y(n_190)
);

INVxp33_ASAP7_75t_SL g191 ( 
.A(n_186),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_191),
.A2(n_181),
.B(n_185),
.Y(n_193)
);

AOI22x1_ASAP7_75t_L g194 ( 
.A1(n_188),
.A2(n_185),
.B1(n_184),
.B2(n_11),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

OAI322xp33_ASAP7_75t_L g196 ( 
.A1(n_193),
.A2(n_187),
.A3(n_188),
.B1(n_192),
.B2(n_191),
.C1(n_190),
.C2(n_25),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_195),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_117),
.B1(n_118),
.B2(n_197),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_196),
.B(n_197),
.Y(n_200)
);


endmodule