module fake_jpeg_19564_n_177 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_177);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_5),
.B(n_11),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_32),
.Y(n_66)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_16),
.B(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_35),
.B(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_18),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_8),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_32),
.B1(n_33),
.B2(n_17),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_17),
.B1(n_23),
.B2(n_18),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_29),
.B1(n_26),
.B2(n_25),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_59),
.A2(n_63),
.B1(n_19),
.B2(n_14),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_9),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_41),
.B1(n_19),
.B2(n_14),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_62),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_66),
.C(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_73),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_0),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_1),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_88),
.B(n_1),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_62),
.B(n_7),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_92),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_0),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_99),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_64),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_107),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_47),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_79),
.C(n_76),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_74),
.B(n_1),
.C(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_47),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_114),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_57),
.B(n_66),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_113),
.B(n_76),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_68),
.B(n_64),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_105),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_119),
.Y(n_135)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_105),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_98),
.A2(n_90),
.B1(n_87),
.B2(n_77),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_128),
.B1(n_75),
.B2(n_73),
.Y(n_141)
);

AO22x1_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_95),
.B1(n_97),
.B2(n_114),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_93),
.B(n_100),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.C(n_102),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_125),
.B1(n_127),
.B2(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_103),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_98),
.A2(n_80),
.B1(n_86),
.B2(n_70),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_130),
.A2(n_110),
.B(n_129),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_101),
.B(n_97),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_134),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_136),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_100),
.B(n_112),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_138),
.B(n_122),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_108),
.B(n_107),
.Y(n_138)
);

XOR2x2_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_142),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_70),
.B1(n_94),
.B2(n_75),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

XOR2x1_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_111),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_124),
.C(n_116),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_148),
.C(n_121),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_145),
.A2(n_137),
.B(n_139),
.Y(n_156)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_151),
.Y(n_157)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_155),
.B(n_158),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_156),
.A2(n_150),
.B(n_126),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_116),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_140),
.C(n_141),
.Y(n_159)
);

AOI31xp67_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_160),
.A3(n_148),
.B(n_157),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_117),
.B1(n_133),
.B2(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_162),
.B(n_96),
.Y(n_168)
);

AOI31xp67_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_143),
.A3(n_151),
.B(n_150),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_163),
.B(n_159),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_2),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_166),
.B(n_169),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_158),
.B(n_155),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_167),
.B(n_168),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_164),
.B(n_3),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_172),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_173),
.B(n_174),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_2),
.B(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_4),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_6),
.Y(n_177)
);


endmodule