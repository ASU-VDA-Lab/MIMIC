module fake_jpeg_16904_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_0),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_0),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_61),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_56),
.B(n_53),
.CON(n_62),
.SN(n_62)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_11),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_68),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_44),
.B1(n_52),
.B2(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_65),
.A2(n_69),
.B1(n_47),
.B2(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_42),
.B1(n_40),
.B2(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_51),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_71),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_7),
.C(n_10),
.Y(n_81)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_65),
.B1(n_74),
.B2(n_66),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_79),
.B1(n_14),
.B2(n_15),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_79),
.B(n_83),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_85),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_90),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_94),
.A2(n_92),
.B(n_93),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_73),
.Y(n_97)
);

AO21x1_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_12),
.B(n_16),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_98),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_17),
.Y(n_100)
);

NAND4xp25_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_18),
.C(n_22),
.D(n_24),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g102 ( 
.A(n_101),
.Y(n_102)
);

AOI21x1_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_25),
.B(n_29),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_103),
.B(n_30),
.Y(n_104)
);


endmodule