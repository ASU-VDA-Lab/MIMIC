module real_aes_11555_n_266 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_266);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_266;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_733;
wire n_602;
wire n_402;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_1175;
wire n_778;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1280;
wire n_394;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g318 ( .A(n_0), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_0), .A2(n_265), .B1(n_419), .B2(n_424), .Y(n_418) );
OAI222xp33_ASAP7_75t_L g949 ( .A1(n_1), .A2(n_38), .B1(n_163), .B2(n_950), .C1(n_952), .C2(n_954), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g980 ( .A1(n_1), .A2(n_163), .B1(n_981), .B2(n_983), .C(n_984), .Y(n_980) );
INVx1_ASAP7_75t_L g1331 ( .A(n_2), .Y(n_1331) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_3), .A2(n_12), .B1(n_355), .B2(n_1001), .Y(n_1000) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_3), .A2(n_12), .B1(n_1037), .B2(n_1038), .Y(n_1036) );
INVxp67_ASAP7_75t_SL g841 ( .A(n_4), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_4), .A2(n_224), .B1(n_424), .B2(n_818), .Y(n_875) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_5), .Y(n_280) );
AND2x2_ASAP7_75t_L g305 ( .A(n_5), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_5), .B(n_210), .Y(n_334) );
INVx1_ASAP7_75t_L g386 ( .A(n_5), .Y(n_386) );
INVx1_ASAP7_75t_L g487 ( .A(n_6), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_6), .A2(n_81), .B1(n_544), .B2(n_546), .Y(n_543) );
INVxp67_ASAP7_75t_L g353 ( .A(n_7), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_7), .A2(n_78), .B1(n_424), .B2(n_451), .Y(n_450) );
OAI221xp5_ASAP7_75t_L g482 ( .A1(n_8), .A2(n_228), .B1(n_335), .B2(n_483), .C(n_484), .Y(n_482) );
OAI22xp33_ASAP7_75t_L g515 ( .A1(n_8), .A2(n_228), .B1(n_516), .B2(n_517), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g1066 ( .A(n_9), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g565 ( .A1(n_10), .A2(n_106), .B1(n_566), .B2(n_567), .C(n_570), .Y(n_565) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_10), .A2(n_148), .B1(n_595), .B2(n_596), .Y(n_594) );
INVx1_ASAP7_75t_L g1100 ( .A(n_11), .Y(n_1100) );
INVx1_ASAP7_75t_L g1366 ( .A(n_13), .Y(n_1366) );
INVxp67_ASAP7_75t_L g840 ( .A(n_14), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g874 ( .A1(n_14), .A2(n_165), .B1(n_444), .B2(n_447), .C(n_664), .Y(n_874) );
INVx1_ASAP7_75t_L g490 ( .A(n_15), .Y(n_490) );
AOI221xp5_ASAP7_75t_L g535 ( .A1(n_15), .A2(n_238), .B1(n_536), .B2(n_538), .C(n_542), .Y(n_535) );
INVxp33_ASAP7_75t_L g788 ( .A(n_16), .Y(n_788) );
AOI221xp5_ASAP7_75t_L g822 ( .A1(n_16), .A2(n_144), .B1(n_444), .B2(n_823), .C(n_824), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g1140 ( .A1(n_17), .A2(n_233), .B1(n_641), .B2(n_1141), .Y(n_1140) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_17), .A2(n_233), .B1(n_1196), .B2(n_1198), .Y(n_1195) );
OAI221xp5_ASAP7_75t_L g1512 ( .A1(n_18), .A2(n_180), .B1(n_483), .B2(n_859), .C(n_1080), .Y(n_1512) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_18), .A2(n_180), .B1(n_437), .B2(n_668), .Y(n_1537) );
INVx1_ASAP7_75t_L g1067 ( .A(n_19), .Y(n_1067) );
AO221x2_ASAP7_75t_L g1301 ( .A1(n_20), .A2(n_55), .B1(n_1285), .B2(n_1294), .C(n_1302), .Y(n_1301) );
INVxp33_ASAP7_75t_L g867 ( .A(n_21), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_21), .A2(n_101), .B1(n_546), .B2(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g1319 ( .A(n_22), .Y(n_1319) );
INVx2_ASAP7_75t_L g399 ( .A(n_23), .Y(n_399) );
OR2x2_ASAP7_75t_L g430 ( .A(n_23), .B(n_397), .Y(n_430) );
INVx1_ASAP7_75t_L g830 ( .A(n_24), .Y(n_830) );
INVx1_ASAP7_75t_L g475 ( .A(n_25), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_25), .A2(n_129), .B1(n_520), .B2(n_522), .C(n_524), .Y(n_519) );
AOI221xp5_ASAP7_75t_L g729 ( .A1(n_26), .A2(n_45), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_729) );
INVx1_ASAP7_75t_L g773 ( .A(n_26), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g645 ( .A(n_27), .Y(n_645) );
INVx1_ASAP7_75t_L g897 ( .A(n_28), .Y(n_897) );
INVx1_ASAP7_75t_L g1303 ( .A(n_29), .Y(n_1303) );
INVx1_ASAP7_75t_L g304 ( .A(n_30), .Y(n_304) );
OR2x2_ASAP7_75t_L g333 ( .A(n_30), .B(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_L g345 ( .A(n_30), .Y(n_345) );
BUFx2_ASAP7_75t_L g393 ( .A(n_30), .Y(n_393) );
INVxp33_ASAP7_75t_L g866 ( .A(n_31), .Y(n_866) );
AOI21xp33_ASAP7_75t_L g881 ( .A1(n_31), .A2(n_412), .B(n_882), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g1055 ( .A1(n_32), .A2(n_40), .B1(n_824), .B2(n_1056), .C(n_1058), .Y(n_1055) );
INVx1_ASAP7_75t_L g1076 ( .A(n_32), .Y(n_1076) );
INVx1_ASAP7_75t_L g1364 ( .A(n_33), .Y(n_1364) );
INVx1_ASAP7_75t_L g1523 ( .A(n_34), .Y(n_1523) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_35), .A2(n_236), .B1(n_451), .B2(n_826), .Y(n_1064) );
INVx1_ASAP7_75t_L g1089 ( .A(n_35), .Y(n_1089) );
INVx1_ASAP7_75t_L g848 ( .A(n_36), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_37), .A2(n_76), .B1(n_994), .B2(n_996), .Y(n_1002) );
INVx1_ASAP7_75t_L g1035 ( .A(n_37), .Y(n_1035) );
INVx1_ASAP7_75t_L g985 ( .A(n_38), .Y(n_985) );
CKINVDCx16_ASAP7_75t_R g1316 ( .A(n_39), .Y(n_1316) );
INVx1_ASAP7_75t_L g1074 ( .A(n_40), .Y(n_1074) );
OAI22xp33_ASAP7_75t_R g1216 ( .A1(n_41), .A2(n_249), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_41), .A2(n_249), .B1(n_339), .B2(n_483), .C(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1360 ( .A(n_42), .Y(n_1360) );
INVx1_ASAP7_75t_L g804 ( .A(n_43), .Y(n_804) );
AOI22xp33_ASAP7_75t_SL g993 ( .A1(n_44), .A2(n_219), .B1(n_994), .B2(n_996), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g1022 ( .A1(n_44), .A2(n_178), .B1(n_820), .B2(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g776 ( .A(n_45), .Y(n_776) );
INVx1_ASAP7_75t_L g751 ( .A(n_46), .Y(n_751) );
INVx1_ASAP7_75t_L g1230 ( .A(n_47), .Y(n_1230) );
INVxp67_ASAP7_75t_SL g579 ( .A(n_48), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_48), .A2(n_104), .B1(n_615), .B2(n_617), .C(n_619), .Y(n_614) );
INVxp67_ASAP7_75t_L g1507 ( .A(n_49), .Y(n_1507) );
AOI221xp5_ASAP7_75t_L g1535 ( .A1(n_49), .A2(n_145), .B1(n_409), .B2(n_415), .C(n_736), .Y(n_1535) );
INVxp67_ASAP7_75t_SL g583 ( .A(n_50), .Y(n_583) );
OAI211xp5_ASAP7_75t_SL g602 ( .A1(n_50), .A2(n_603), .B(n_606), .C(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g586 ( .A(n_51), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_52), .A2(n_95), .B1(n_599), .B2(n_904), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_52), .A2(n_195), .B1(n_424), .B2(n_925), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_53), .A2(n_204), .B1(n_659), .B2(n_661), .Y(n_658) );
INVx1_ASAP7_75t_L g693 ( .A(n_53), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_54), .A2(n_72), .B1(n_1132), .B2(n_1133), .Y(n_1131) );
INVxp67_ASAP7_75t_L g1181 ( .A(n_54), .Y(n_1181) );
XNOR2x2_ASAP7_75t_L g986 ( .A(n_55), .B(n_987), .Y(n_986) );
INVxp33_ASAP7_75t_L g1515 ( .A(n_56), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_56), .A2(n_222), .B1(n_823), .B2(n_1542), .Y(n_1541) );
INVxp33_ASAP7_75t_L g864 ( .A(n_57), .Y(n_864) );
NAND2xp33_ASAP7_75t_SL g879 ( .A(n_57), .B(n_880), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_58), .Y(n_509) );
OAI222xp33_ASAP7_75t_L g955 ( .A1(n_59), .A2(n_140), .B1(n_218), .B2(n_585), .C1(n_829), .C2(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g961 ( .A(n_59), .Y(n_961) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_60), .Y(n_1011) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_61), .A2(n_139), .B1(n_1132), .B2(n_1211), .C(n_1212), .Y(n_1210) );
INVxp33_ASAP7_75t_L g1235 ( .A(n_61), .Y(n_1235) );
INVx1_ASAP7_75t_L g1264 ( .A(n_62), .Y(n_1264) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_63), .A2(n_178), .B1(n_617), .B2(n_999), .Y(n_998) );
AOI21xp33_ASAP7_75t_L g1025 ( .A1(n_63), .A2(n_742), .B(n_1026), .Y(n_1025) );
CKINVDCx16_ASAP7_75t_R g1278 ( .A(n_64), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_65), .A2(n_471), .B1(n_554), .B2(n_555), .Y(n_470) );
INVx1_ASAP7_75t_L g554 ( .A(n_65), .Y(n_554) );
AOI22xp33_ASAP7_75t_SL g562 ( .A1(n_66), .A2(n_148), .B1(n_451), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_66), .A2(n_106), .B1(n_598), .B2(n_599), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_67), .A2(n_141), .B1(n_424), .B2(n_925), .Y(n_946) );
INVx1_ASAP7_75t_L g978 ( .A(n_67), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_68), .A2(n_89), .B1(n_572), .B2(n_746), .Y(n_943) );
INVx1_ASAP7_75t_L g966 ( .A(n_68), .Y(n_966) );
INVx1_ASAP7_75t_L g887 ( .A(n_69), .Y(n_887) );
INVxp67_ASAP7_75t_L g347 ( .A(n_70), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_70), .A2(n_183), .B1(n_443), .B2(n_444), .C(n_447), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_71), .A2(n_98), .B1(n_563), .B2(n_572), .Y(n_571) );
INVxp67_ASAP7_75t_SL g625 ( .A(n_71), .Y(n_625) );
INVxp67_ASAP7_75t_L g1179 ( .A(n_72), .Y(n_1179) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_73), .A2(n_150), .B1(n_415), .B2(n_451), .C(n_575), .Y(n_574) );
INVxp33_ASAP7_75t_SL g610 ( .A(n_73), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g1225 ( .A1(n_74), .A2(n_235), .B1(n_1226), .B2(n_1228), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1249 ( .A(n_74), .Y(n_1249) );
INVx1_ASAP7_75t_L g1332 ( .A(n_75), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_76), .B(n_460), .Y(n_1017) );
INVx1_ASAP7_75t_L g1014 ( .A(n_77), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_77), .A2(n_132), .B1(n_1023), .B2(n_1026), .Y(n_1030) );
INVxp67_ASAP7_75t_L g359 ( .A(n_78), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g858 ( .A1(n_79), .A2(n_176), .B1(n_326), .B2(n_335), .C(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g883 ( .A(n_79), .Y(n_883) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_80), .A2(n_243), .B1(n_633), .B2(n_635), .C(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g677 ( .A(n_80), .Y(n_677) );
INVx1_ASAP7_75t_L g499 ( .A(n_81), .Y(n_499) );
OA22x2_ASAP7_75t_L g1201 ( .A1(n_82), .A2(n_1202), .B1(n_1203), .B2(n_1253), .Y(n_1201) );
CKINVDCx16_ASAP7_75t_R g1253 ( .A(n_82), .Y(n_1253) );
AOI22xp5_ASAP7_75t_L g1299 ( .A1(n_83), .A2(n_142), .B1(n_1288), .B2(n_1291), .Y(n_1299) );
INVx1_ASAP7_75t_L g397 ( .A(n_84), .Y(n_397) );
INVx1_ASAP7_75t_L g417 ( .A(n_84), .Y(n_417) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_85), .Y(n_1205) );
INVx1_ASAP7_75t_L g1117 ( .A(n_86), .Y(n_1117) );
INVx1_ASAP7_75t_L g1006 ( .A(n_87), .Y(n_1006) );
AOI21xp5_ASAP7_75t_L g1031 ( .A1(n_87), .A2(n_545), .B(n_648), .Y(n_1031) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_88), .A2(n_262), .B1(n_432), .B2(n_517), .Y(n_728) );
INVx1_ASAP7_75t_L g755 ( .A(n_88), .Y(n_755) );
INVx1_ASAP7_75t_L g963 ( .A(n_89), .Y(n_963) );
INVx1_ASAP7_75t_L g1531 ( .A(n_90), .Y(n_1531) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_91), .A2(n_120), .B1(n_326), .B2(n_335), .C(n_339), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_91), .A2(n_120), .B1(n_432), .B2(n_437), .Y(n_431) );
INVxp67_ASAP7_75t_SL g797 ( .A(n_92), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_92), .A2(n_213), .B1(n_447), .B2(n_566), .C(n_664), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g479 ( .A(n_93), .Y(n_479) );
INVx1_ASAP7_75t_L g931 ( .A(n_94), .Y(n_931) );
AOI221xp5_ASAP7_75t_L g921 ( .A1(n_95), .A2(n_170), .B1(n_447), .B2(n_922), .C(n_923), .Y(n_921) );
INVxp33_ASAP7_75t_SL g785 ( .A(n_96), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_96), .A2(n_117), .B1(n_443), .B2(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_97), .A2(n_244), .B1(n_599), .B2(n_908), .Y(n_907) );
INVxp67_ASAP7_75t_L g920 ( .A(n_97), .Y(n_920) );
INVxp33_ASAP7_75t_L g611 ( .A(n_98), .Y(n_611) );
INVxp67_ASAP7_75t_L g1511 ( .A(n_99), .Y(n_1511) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_99), .A2(n_192), .B1(n_732), .B2(n_953), .Y(n_1536) );
INVxp33_ASAP7_75t_SL g899 ( .A(n_100), .Y(n_899) );
AOI21xp33_ASAP7_75t_L g918 ( .A1(n_100), .A2(n_531), .B(n_820), .Y(n_918) );
INVxp33_ASAP7_75t_L g862 ( .A(n_101), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_102), .A2(n_156), .B1(n_444), .B2(n_447), .C(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1085 ( .A(n_102), .Y(n_1085) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_103), .Y(n_477) );
OAI211xp5_ASAP7_75t_SL g560 ( .A1(n_104), .A2(n_465), .B(n_561), .C(n_577), .Y(n_560) );
INVx1_ASAP7_75t_L g1318 ( .A(n_105), .Y(n_1318) );
AO221x2_ASAP7_75t_L g1329 ( .A1(n_107), .A2(n_191), .B1(n_1280), .B2(n_1285), .C(n_1330), .Y(n_1329) );
CKINVDCx5p33_ASAP7_75t_R g637 ( .A(n_108), .Y(n_637) );
INVx1_ASAP7_75t_L g1545 ( .A(n_109), .Y(n_1545) );
OAI22xp33_ASAP7_75t_SL g662 ( .A1(n_110), .A2(n_215), .B1(n_663), .B2(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g696 ( .A(n_110), .Y(n_696) );
INVx1_ASAP7_75t_L g802 ( .A(n_111), .Y(n_802) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_111), .A2(n_177), .B1(n_424), .B2(n_818), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_112), .Y(n_1054) );
INVxp33_ASAP7_75t_SL g1109 ( .A(n_113), .Y(n_1109) );
AOI221xp5_ASAP7_75t_L g1168 ( .A1(n_113), .A2(n_157), .B1(n_770), .B2(n_908), .C(n_1169), .Y(n_1168) );
OAI22xp33_ASAP7_75t_L g1060 ( .A1(n_114), .A2(n_239), .B1(n_668), .B2(n_829), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_114), .A2(n_239), .B1(n_339), .B2(n_1079), .C(n_1080), .Y(n_1078) );
INVx1_ASAP7_75t_L g272 ( .A(n_115), .Y(n_272) );
INVx1_ASAP7_75t_L g851 ( .A(n_116), .Y(n_851) );
INVxp33_ASAP7_75t_SL g789 ( .A(n_117), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g1134 ( .A1(n_118), .A2(n_190), .B1(n_544), .B2(n_1135), .Y(n_1134) );
INVxp67_ASAP7_75t_SL g1191 ( .A(n_118), .Y(n_1191) );
XNOR2x1_ASAP7_75t_L g292 ( .A(n_119), .B(n_293), .Y(n_292) );
INVxp67_ASAP7_75t_SL g893 ( .A(n_121), .Y(n_893) );
OAI221xp5_ASAP7_75t_L g914 ( .A1(n_121), .A2(n_200), .B1(n_437), .B2(n_828), .C(n_915), .Y(n_914) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_122), .A2(n_158), .B1(n_536), .B2(n_641), .C(n_642), .Y(n_640) );
INVx1_ASAP7_75t_L g700 ( .A(n_122), .Y(n_700) );
INVx1_ASAP7_75t_L g368 ( .A(n_123), .Y(n_368) );
INVx1_ASAP7_75t_L g740 ( .A(n_124), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_124), .A2(n_167), .B1(n_769), .B2(n_770), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g1300 ( .A1(n_125), .A2(n_184), .B1(n_1285), .B2(n_1294), .Y(n_1300) );
CKINVDCx5p33_ASAP7_75t_R g646 ( .A(n_126), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g1222 ( .A1(n_127), .A2(n_214), .B1(n_536), .B2(n_1223), .C(n_1224), .Y(n_1222) );
INVxp67_ASAP7_75t_SL g1244 ( .A(n_127), .Y(n_1244) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_128), .Y(n_502) );
INVx1_ASAP7_75t_L g480 ( .A(n_129), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g906 ( .A1(n_130), .A2(n_221), .B1(n_497), .B2(n_595), .Y(n_906) );
INVxp33_ASAP7_75t_L g930 ( .A(n_130), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g944 ( .A1(n_131), .A2(n_186), .B1(n_444), .B2(n_742), .C(n_945), .Y(n_944) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_131), .A2(n_141), .B1(n_973), .B2(n_975), .C(n_977), .Y(n_972) );
INVx1_ASAP7_75t_L g1010 ( .A(n_132), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_133), .A2(n_245), .B1(n_744), .B2(n_746), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_133), .A2(n_143), .B1(n_507), .B2(n_595), .Y(n_764) );
INVx1_ASAP7_75t_L g778 ( .A(n_134), .Y(n_778) );
INVx1_ASAP7_75t_L g854 ( .A(n_135), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_136), .Y(n_508) );
INVx1_ASAP7_75t_L g1304 ( .A(n_137), .Y(n_1304) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_138), .A2(n_153), .B1(n_412), .B2(n_415), .C(n_922), .Y(n_942) );
INVx1_ASAP7_75t_L g964 ( .A(n_138), .Y(n_964) );
INVxp33_ASAP7_75t_L g1237 ( .A(n_139), .Y(n_1237) );
INVx1_ASAP7_75t_L g967 ( .A(n_140), .Y(n_967) );
AOI221xp5_ASAP7_75t_L g741 ( .A1(n_143), .A2(n_149), .B1(n_567), .B2(n_653), .C(n_742), .Y(n_741) );
INVxp33_ASAP7_75t_L g786 ( .A(n_144), .Y(n_786) );
INVxp67_ASAP7_75t_L g1510 ( .A(n_145), .Y(n_1510) );
INVx1_ASAP7_75t_L g379 ( .A(n_146), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_147), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g758 ( .A1(n_149), .A2(n_245), .B1(n_759), .B2(n_761), .Y(n_758) );
OAI21xp33_ASAP7_75t_SL g591 ( .A1(n_150), .A2(n_592), .B(n_593), .Y(n_591) );
INVx1_ASAP7_75t_L g750 ( .A(n_151), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_151), .A2(n_185), .B1(n_595), .B2(n_766), .Y(n_765) );
INVxp33_ASAP7_75t_SL g900 ( .A(n_152), .Y(n_900) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_152), .A2(n_212), .B1(n_425), .B2(n_569), .Y(n_917) );
INVx1_ASAP7_75t_L g971 ( .A(n_153), .Y(n_971) );
CKINVDCx5p33_ASAP7_75t_R g948 ( .A(n_154), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_155), .A2(n_188), .B1(n_567), .B2(n_641), .Y(n_1059) );
INVx1_ASAP7_75t_L g1072 ( .A(n_155), .Y(n_1072) );
INVx1_ASAP7_75t_L g1087 ( .A(n_156), .Y(n_1087) );
INVxp33_ASAP7_75t_SL g1105 ( .A(n_157), .Y(n_1105) );
INVx1_ASAP7_75t_L g702 ( .A(n_158), .Y(n_702) );
AOI22xp33_ASAP7_75t_SL g1137 ( .A1(n_159), .A2(n_168), .B1(n_1135), .B2(n_1138), .Y(n_1137) );
OAI211xp5_ASAP7_75t_SL g1158 ( .A1(n_159), .A2(n_1159), .B(n_1164), .C(n_1170), .Y(n_1158) );
CKINVDCx5p33_ASAP7_75t_R g1051 ( .A(n_160), .Y(n_1051) );
XNOR2xp5_ASAP7_75t_L g1095 ( .A(n_161), .B(n_1096), .Y(n_1095) );
OAI221xp5_ASAP7_75t_L g790 ( .A1(n_162), .A2(n_263), .B1(n_326), .B2(n_336), .C(n_339), .Y(n_790) );
OAI22xp33_ASAP7_75t_L g827 ( .A1(n_162), .A2(n_263), .B1(n_828), .B2(n_829), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g1307 ( .A1(n_164), .A2(n_172), .B1(n_1288), .B2(n_1291), .Y(n_1307) );
INVxp33_ASAP7_75t_L g846 ( .A(n_165), .Y(n_846) );
INVxp67_ASAP7_75t_L g1519 ( .A(n_166), .Y(n_1519) );
AOI221xp5_ASAP7_75t_L g1539 ( .A1(n_166), .A2(n_226), .B1(n_542), .B2(n_573), .C(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g749 ( .A(n_167), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g1175 ( .A1(n_168), .A2(n_1176), .B1(n_1178), .B2(n_1187), .C(n_1194), .Y(n_1175) );
INVx1_ASAP7_75t_L g1215 ( .A(n_169), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_170), .A2(n_195), .B1(n_595), .B2(n_856), .Y(n_905) );
CKINVDCx5p33_ASAP7_75t_R g991 ( .A(n_171), .Y(n_991) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_173), .Y(n_652) );
INVx1_ASAP7_75t_L g780 ( .A(n_174), .Y(n_780) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_175), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g1267 ( .A(n_175), .B(n_272), .Y(n_1267) );
AND3x2_ASAP7_75t_L g1283 ( .A(n_175), .B(n_272), .C(n_1270), .Y(n_1283) );
INVx1_ASAP7_75t_L g884 ( .A(n_176), .Y(n_884) );
INVxp67_ASAP7_75t_SL g796 ( .A(n_177), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g1308 ( .A1(n_179), .A2(n_217), .B1(n_1280), .B2(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1208 ( .A(n_181), .Y(n_1208) );
INVx2_ASAP7_75t_L g285 ( .A(n_182), .Y(n_285) );
INVxp33_ASAP7_75t_L g366 ( .A(n_183), .Y(n_366) );
INVx1_ASAP7_75t_L g727 ( .A(n_185), .Y(n_727) );
INVx1_ASAP7_75t_L g979 ( .A(n_186), .Y(n_979) );
AOI22xp5_ASAP7_75t_L g1293 ( .A1(n_187), .A2(n_197), .B1(n_1285), .B2(n_1294), .Y(n_1293) );
INVxp67_ASAP7_75t_L g1501 ( .A(n_187), .Y(n_1501) );
AOI22xp33_ASAP7_75t_L g1552 ( .A1(n_187), .A2(n_1553), .B1(n_1557), .B2(n_1562), .Y(n_1552) );
INVx1_ASAP7_75t_L g1077 ( .A(n_188), .Y(n_1077) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_189), .Y(n_512) );
INVxp67_ASAP7_75t_SL g1190 ( .A(n_190), .Y(n_1190) );
INVxp67_ASAP7_75t_L g1506 ( .A(n_192), .Y(n_1506) );
INVx1_ASAP7_75t_L g371 ( .A(n_193), .Y(n_371) );
XNOR2xp5_ASAP7_75t_L g1046 ( .A(n_194), .B(n_1047), .Y(n_1046) );
INVx1_ASAP7_75t_L g1270 ( .A(n_196), .Y(n_1270) );
CKINVDCx16_ASAP7_75t_R g1315 ( .A(n_198), .Y(n_1315) );
XNOR2x1_ASAP7_75t_L g889 ( .A(n_199), .B(n_890), .Y(n_889) );
INVx1_ASAP7_75t_L g1362 ( .A(n_199), .Y(n_1362) );
INVxp67_ASAP7_75t_SL g894 ( .A(n_200), .Y(n_894) );
OAI211xp5_ASAP7_75t_SL g580 ( .A1(n_201), .A2(n_581), .B(n_582), .C(n_588), .Y(n_580) );
INVx1_ASAP7_75t_L g622 ( .A(n_201), .Y(n_622) );
INVx1_ASAP7_75t_L g1221 ( .A(n_202), .Y(n_1221) );
AOI22x1_ASAP7_75t_L g834 ( .A1(n_203), .A2(n_835), .B1(n_836), .B2(n_888), .Y(n_834) );
INVx1_ASAP7_75t_L g888 ( .A(n_203), .Y(n_888) );
INVx1_ASAP7_75t_L g695 ( .A(n_204), .Y(n_695) );
INVx1_ASAP7_75t_L g1213 ( .A(n_205), .Y(n_1213) );
INVx1_ASAP7_75t_L g1015 ( .A(n_206), .Y(n_1015) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_206), .A2(n_585), .B(n_1034), .C(n_1039), .Y(n_1033) );
INVx1_ASAP7_75t_L g807 ( .A(n_207), .Y(n_807) );
INVx1_ASAP7_75t_L g1530 ( .A(n_208), .Y(n_1530) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_209), .Y(n_671) );
INVx1_ASAP7_75t_L g287 ( .A(n_210), .Y(n_287) );
INVx2_ASAP7_75t_L g306 ( .A(n_210), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_211), .Y(n_670) );
INVxp33_ASAP7_75t_SL g896 ( .A(n_212), .Y(n_896) );
INVxp67_ASAP7_75t_SL g801 ( .A(n_213), .Y(n_801) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_214), .Y(n_1248) );
INVx1_ASAP7_75t_L g690 ( .A(n_215), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g1287 ( .A1(n_216), .A2(n_237), .B1(n_1288), .B2(n_1291), .Y(n_1287) );
INVx1_ASAP7_75t_L g960 ( .A(n_218), .Y(n_960) );
INVx1_ASAP7_75t_L g1020 ( .A(n_219), .Y(n_1020) );
INVxp33_ASAP7_75t_L g313 ( .A(n_220), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_220), .A2(n_223), .B1(n_409), .B2(n_412), .C(n_415), .Y(n_408) );
INVxp67_ASAP7_75t_L g913 ( .A(n_221), .Y(n_913) );
INVxp67_ASAP7_75t_L g1520 ( .A(n_222), .Y(n_1520) );
INVxp33_ASAP7_75t_L g307 ( .A(n_223), .Y(n_307) );
INVxp33_ASAP7_75t_L g843 ( .A(n_224), .Y(n_843) );
INVx1_ASAP7_75t_L g805 ( .A(n_225), .Y(n_805) );
INVxp33_ASAP7_75t_L g1516 ( .A(n_226), .Y(n_1516) );
INVx1_ASAP7_75t_L g1113 ( .A(n_227), .Y(n_1113) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_229), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g1558 ( .A1(n_230), .A2(n_1559), .B1(n_1560), .B2(n_1561), .Y(n_1558) );
CKINVDCx5p33_ASAP7_75t_R g1559 ( .A(n_230), .Y(n_1559) );
INVx1_ASAP7_75t_L g1272 ( .A(n_231), .Y(n_1272) );
INVx1_ASAP7_75t_L g375 ( .A(n_232), .Y(n_375) );
INVx1_ASAP7_75t_L g1271 ( .A(n_234), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_234), .B(n_1269), .Y(n_1276) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_235), .Y(n_1243) );
INVx1_ASAP7_75t_L g1084 ( .A(n_236), .Y(n_1084) );
INVx1_ASAP7_75t_L g495 ( .A(n_238), .Y(n_495) );
INVx1_ASAP7_75t_L g587 ( .A(n_240), .Y(n_587) );
INVx1_ASAP7_75t_L g1123 ( .A(n_241), .Y(n_1123) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_242), .Y(n_405) );
INVx1_ASAP7_75t_L g686 ( .A(n_243), .Y(n_686) );
INVxp33_ASAP7_75t_L g929 ( .A(n_244), .Y(n_929) );
INVx1_ASAP7_75t_L g1525 ( .A(n_246), .Y(n_1525) );
AOI22x1_ASAP7_75t_L g557 ( .A1(n_247), .A2(n_558), .B1(n_627), .B2(n_628), .Y(n_557) );
INVxp67_ASAP7_75t_L g627 ( .A(n_247), .Y(n_627) );
CKINVDCx5p33_ASAP7_75t_R g1052 ( .A(n_248), .Y(n_1052) );
INVx1_ASAP7_75t_L g1231 ( .A(n_250), .Y(n_1231) );
AOI21xp5_ASAP7_75t_L g735 ( .A1(n_251), .A2(n_531), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g775 ( .A(n_251), .Y(n_775) );
INVx1_ASAP7_75t_L g857 ( .A(n_252), .Y(n_857) );
INVx2_ASAP7_75t_L g284 ( .A(n_253), .Y(n_284) );
XNOR2x1_ASAP7_75t_L g938 ( .A(n_254), .B(n_939), .Y(n_938) );
CKINVDCx5p33_ASAP7_75t_R g1149 ( .A(n_255), .Y(n_1149) );
XNOR2x2_ASAP7_75t_L g629 ( .A(n_256), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g808 ( .A(n_257), .Y(n_808) );
BUFx3_ASAP7_75t_L g402 ( .A(n_258), .Y(n_402) );
INVx1_ASAP7_75t_L g427 ( .A(n_258), .Y(n_427) );
BUFx3_ASAP7_75t_L g404 ( .A(n_259), .Y(n_404) );
INVx1_ASAP7_75t_L g423 ( .A(n_259), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_260), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_261), .Y(n_734) );
INVx1_ASAP7_75t_L g754 ( .A(n_262), .Y(n_754) );
INVx1_ASAP7_75t_L g578 ( .A(n_264), .Y(n_578) );
INVxp33_ASAP7_75t_L g297 ( .A(n_265), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_288), .B(n_1256), .Y(n_266) );
BUFx12f_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_275), .Y(n_269) );
AND2x4_ASAP7_75t_L g1551 ( .A(n_270), .B(n_276), .Y(n_1551) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_SL g1556 ( .A(n_271), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1569 ( .A(n_271), .B(n_273), .Y(n_1569) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_273), .B(n_1556), .Y(n_1555) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g601 ( .A(n_279), .B(n_287), .Y(n_601) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g343 ( .A(n_280), .B(n_344), .Y(n_343) );
OR2x6_ASAP7_75t_L g281 ( .A(n_282), .B(n_286), .Y(n_281) );
INVx2_ASAP7_75t_SL g358 ( .A(n_282), .Y(n_358) );
INVx2_ASAP7_75t_SL g374 ( .A(n_282), .Y(n_374) );
OR2x2_ASAP7_75t_L g390 ( .A(n_282), .B(n_333), .Y(n_390) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_282), .Y(n_501) );
BUFx2_ASAP7_75t_L g605 ( .A(n_282), .Y(n_605) );
INVx1_ASAP7_75t_L g621 ( .A(n_282), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g984 ( .A1(n_282), .A2(n_362), .B1(n_948), .B2(n_985), .Y(n_984) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_L g301 ( .A(n_284), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g311 ( .A(n_284), .Y(n_311) );
AND2x2_ASAP7_75t_L g317 ( .A(n_284), .B(n_285), .Y(n_317) );
INVx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
INVx1_ASAP7_75t_L g365 ( .A(n_284), .Y(n_365) );
INVx2_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
INVx1_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
INVx1_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_285), .B(n_322), .Y(n_352) );
INVx1_ASAP7_75t_L g364 ( .A(n_285), .Y(n_364) );
INVx2_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OAI22xp33_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_1040), .B1(n_1041), .B2(n_1255), .Y(n_288) );
INVx1_ASAP7_75t_L g1255 ( .A(n_289), .Y(n_1255) );
XNOR2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_718), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_556), .B1(n_716), .B2(n_717), .Y(n_290) );
INVxp33_ASAP7_75t_L g717 ( .A(n_291), .Y(n_717) );
XOR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_470), .Y(n_291) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_387), .Y(n_293) );
NOR3xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_325), .C(n_341), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_312), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_298), .B1(n_307), .B2(n_308), .Y(n_296) );
BUFx2_ASAP7_75t_L g476 ( .A(n_298), .Y(n_476) );
BUFx2_ASAP7_75t_L g626 ( .A(n_298), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_298), .A2(n_308), .B1(n_645), .B2(n_700), .Y(n_699) );
BUFx2_ASAP7_75t_L g863 ( .A(n_298), .Y(n_863) );
BUFx2_ASAP7_75t_L g1073 ( .A(n_298), .Y(n_1073) );
AOI22xp33_ASAP7_75t_L g1236 ( .A1(n_298), .A2(n_1213), .B1(n_1237), .B2(n_1238), .Y(n_1236) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
BUFx3_ASAP7_75t_L g507 ( .A(n_299), .Y(n_507) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g370 ( .A(n_300), .Y(n_370) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_300), .Y(n_618) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_301), .Y(n_355) );
INVx1_ASAP7_75t_L g1186 ( .A(n_301), .Y(n_1186) );
AND2x4_ASAP7_75t_L g310 ( .A(n_302), .B(n_311), .Y(n_310) );
AND2x6_ASAP7_75t_L g308 ( .A(n_303), .B(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g314 ( .A(n_303), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_303), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g481 ( .A(n_303), .B(n_320), .Y(n_481) );
AND2x2_ASAP7_75t_L g612 ( .A(n_303), .B(n_320), .Y(n_612) );
AND2x2_ASAP7_75t_L g777 ( .A(n_303), .B(n_320), .Y(n_777) );
AND2x2_ASAP7_75t_L g969 ( .A(n_303), .B(n_970), .Y(n_969) );
AND2x2_ASAP7_75t_L g1009 ( .A(n_303), .B(n_320), .Y(n_1009) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_303), .B(n_370), .Y(n_1013) );
AND2x2_ASAP7_75t_L g1508 ( .A(n_303), .B(n_771), .Y(n_1508) );
AND2x4_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
INVx1_ASAP7_75t_L g383 ( .A(n_304), .Y(n_383) );
OR2x2_ASAP7_75t_L g1104 ( .A(n_304), .B(n_430), .Y(n_1104) );
INVx2_ASAP7_75t_L g1162 ( .A(n_305), .Y(n_1162) );
AND2x4_ASAP7_75t_L g1177 ( .A(n_305), .B(n_760), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_305), .B(n_321), .Y(n_1197) );
INVx1_ASAP7_75t_L g344 ( .A(n_306), .Y(n_344) );
INVx1_ASAP7_75t_L g385 ( .A(n_306), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_308), .A2(n_475), .B1(n_476), .B2(n_477), .Y(n_474) );
INVx1_ASAP7_75t_SL g592 ( .A(n_308), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_308), .A2(n_626), .B1(n_734), .B2(n_773), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_308), .A2(n_626), .B1(n_785), .B2(n_786), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_308), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g895 ( .A1(n_308), .A2(n_863), .B1(n_896), .B2(n_897), .Y(n_895) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_308), .A2(n_777), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_308), .A2(n_1009), .B1(n_1010), .B2(n_1011), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_308), .A2(n_1072), .B1(n_1073), .B2(n_1074), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1238 ( .A(n_308), .Y(n_1238) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_309), .B(n_332), .Y(n_340) );
BUFx2_ASAP7_75t_L g599 ( .A(n_309), .Y(n_599) );
BUFx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx2_ASAP7_75t_L g715 ( .A(n_310), .Y(n_715) );
BUFx6f_ASAP7_75t_L g763 ( .A(n_310), .Y(n_763) );
BUFx6f_ASAP7_75t_L g771 ( .A(n_310), .Y(n_771) );
INVx1_ASAP7_75t_L g997 ( .A(n_310), .Y(n_997) );
BUFx3_ASAP7_75t_L g1163 ( .A(n_310), .Y(n_1163) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_318), .B2(n_319), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_314), .A2(n_479), .B1(n_480), .B2(n_481), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_314), .A2(n_610), .B1(n_611), .B2(n_612), .Y(n_609) );
BUFx2_ASAP7_75t_L g674 ( .A(n_314), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_314), .A2(n_775), .B1(n_776), .B2(n_777), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g787 ( .A1(n_314), .A2(n_777), .B1(n_788), .B2(n_789), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_314), .A2(n_777), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g898 ( .A1(n_314), .A2(n_612), .B1(n_899), .B2(n_900), .Y(n_898) );
NAND2xp5_ASAP7_75t_L g1005 ( .A(n_314), .B(n_1006), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_314), .A2(n_319), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
INVx2_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g598 ( .A(n_316), .Y(n_598) );
INVx2_ASAP7_75t_SL g970 ( .A(n_316), .Y(n_970) );
INVx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
BUFx6f_ASAP7_75t_L g760 ( .A(n_317), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g1234 ( .A1(n_319), .A2(n_674), .B1(n_1215), .B2(n_1235), .Y(n_1234) );
INVx2_ASAP7_75t_SL g616 ( .A(n_320), .Y(n_616) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
BUFx2_ASAP7_75t_L g595 ( .A(n_321), .Y(n_595) );
INVx1_ASAP7_75t_L g974 ( .A(n_321), .Y(n_974) );
INVx1_ASAP7_75t_L g982 ( .A(n_321), .Y(n_982) );
BUFx6f_ASAP7_75t_L g999 ( .A(n_321), .Y(n_999) );
BUFx6f_ASAP7_75t_L g1001 ( .A(n_321), .Y(n_1001) );
AND2x4_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
INVx1_ASAP7_75t_L g338 ( .A(n_322), .Y(n_338) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g483 ( .A(n_327), .Y(n_483) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
HB1xp67_ASAP7_75t_L g1079 ( .A(n_328), .Y(n_1079) );
NAND2x1_ASAP7_75t_SL g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_329), .A2(n_337), .B1(n_586), .B2(n_587), .Y(n_607) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
HB1xp67_ASAP7_75t_L g713 ( .A(n_331), .Y(n_713) );
NAND2x1p5_ASAP7_75t_L g336 ( .A(n_332), .B(n_337), .Y(n_336) );
AOI32xp33_ASAP7_75t_L g593 ( .A1(n_332), .A2(n_594), .A3(n_597), .B1(n_600), .B2(n_602), .Y(n_593) );
AND2x4_ASAP7_75t_L g707 ( .A(n_332), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g712 ( .A(n_332), .B(n_713), .Y(n_712) );
AND2x4_ASAP7_75t_L g714 ( .A(n_332), .B(n_715), .Y(n_714) );
INVx3_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g1156 ( .A(n_334), .Y(n_1156) );
BUFx4f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx4f_ASAP7_75t_L g1080 ( .A(n_336), .Y(n_1080) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x6_ASAP7_75t_L g1174 ( .A(n_338), .B(n_1155), .Y(n_1174) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx2_ASAP7_75t_L g484 ( .A(n_340), .Y(n_484) );
BUFx3_ASAP7_75t_L g859 ( .A(n_340), .Y(n_859) );
OAI33xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_346), .A3(n_356), .B1(n_367), .B2(n_372), .B3(n_380), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g485 ( .A1(n_342), .A2(n_380), .A3(n_486), .B1(n_491), .B2(n_500), .B3(n_505), .Y(n_485) );
OAI33xp33_ASAP7_75t_L g675 ( .A1(n_342), .A2(n_676), .A3(n_682), .B1(n_687), .B2(n_694), .B3(n_697), .Y(n_675) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_342), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g838 ( .A1(n_342), .A2(n_380), .A3(n_839), .B1(n_842), .B2(n_847), .B3(n_852), .Y(n_838) );
OAI33xp33_ASAP7_75t_L g1081 ( .A1(n_342), .A2(n_380), .A3(n_1082), .B1(n_1086), .B2(n_1091), .B3(n_1092), .Y(n_1081) );
OAI33xp33_ASAP7_75t_L g1241 ( .A1(n_342), .A2(n_1242), .A3(n_1245), .B1(n_1250), .B2(n_1251), .B3(n_1252), .Y(n_1241) );
OAI33xp33_ASAP7_75t_L g1513 ( .A1(n_342), .A2(n_1252), .A3(n_1514), .B1(n_1518), .B2(n_1522), .B3(n_1529), .Y(n_1513) );
OR2x6_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
BUFx2_ASAP7_75t_L g469 ( .A(n_345), .Y(n_469) );
INVx2_ASAP7_75t_L g553 ( .A(n_345), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_353), .B2(n_354), .Y(n_346) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_348), .A2(n_368), .B1(n_369), .B2(n_371), .Y(n_367) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g1088 ( .A(n_349), .Y(n_1088) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx2_ASAP7_75t_L g503 ( .A(n_350), .Y(n_503) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx3_ASAP7_75t_L g689 ( .A(n_351), .Y(n_689) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g494 ( .A(n_352), .Y(n_494) );
INVx1_ASAP7_75t_L g685 ( .A(n_352), .Y(n_685) );
INVx2_ASAP7_75t_L g596 ( .A(n_354), .Y(n_596) );
OAI22xp5_ASAP7_75t_L g798 ( .A1(n_354), .A2(n_799), .B1(n_801), .B2(n_802), .Y(n_798) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_354), .A2(n_503), .B1(n_804), .B2(n_805), .Y(n_803) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
BUFx3_ASAP7_75t_L g856 ( .A(n_355), .Y(n_856) );
INVx2_ASAP7_75t_SL g1167 ( .A(n_355), .Y(n_1167) );
OAI22xp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_359), .B1(n_360), .B2(n_366), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g1187 ( .A1(n_357), .A2(n_1188), .B1(n_1190), .B2(n_1191), .C(n_1192), .Y(n_1187) );
OAI22xp33_ASAP7_75t_L g1242 ( .A1(n_357), .A2(n_606), .B1(n_1243), .B2(n_1244), .Y(n_1242) );
OAI22xp33_ASAP7_75t_L g1250 ( .A1(n_357), .A2(n_1180), .B1(n_1208), .B2(n_1230), .Y(n_1250) );
OAI22xp5_ASAP7_75t_SL g1529 ( .A1(n_357), .A2(n_606), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g842 ( .A1(n_360), .A2(n_843), .B1(n_844), .B2(n_846), .Y(n_842) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g606 ( .A(n_361), .Y(n_606) );
INVx2_ASAP7_75t_L g623 ( .A(n_361), .Y(n_623) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_362), .A2(n_605), .B1(n_978), .B2(n_979), .Y(n_977) );
BUFx3_ASAP7_75t_L g1189 ( .A(n_362), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
AND2x2_ASAP7_75t_L g378 ( .A(n_364), .B(n_365), .Y(n_378) );
INVx1_ASAP7_75t_L g709 ( .A(n_365), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_368), .A2(n_408), .B1(n_418), .B2(n_428), .C(n_431), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_369), .A2(n_799), .B1(n_840), .B2(n_841), .Y(n_839) );
INVx2_ASAP7_75t_L g983 ( .A(n_369), .Y(n_983) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g498 ( .A(n_370), .Y(n_498) );
INVx2_ASAP7_75t_L g767 ( .A(n_370), .Y(n_767) );
INVx2_ASAP7_75t_L g976 ( .A(n_370), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_371), .A2(n_375), .B1(n_459), .B2(n_464), .Y(n_458) );
OAI22xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_375), .B1(n_376), .B2(n_379), .Y(n_372) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_373), .A2(n_487), .B1(n_488), .B2(n_490), .Y(n_486) );
INVx3_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g793 ( .A1(n_376), .A2(n_794), .B1(n_796), .B2(n_797), .Y(n_793) );
BUFx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g489 ( .A(n_377), .Y(n_489) );
INVx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g681 ( .A(n_378), .Y(n_681) );
BUFx2_ASAP7_75t_L g850 ( .A(n_378), .Y(n_850) );
INVx2_ASAP7_75t_L g1517 ( .A(n_378), .Y(n_1517) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_379), .A2(n_442), .B1(n_450), .B2(n_453), .C(n_455), .Y(n_441) );
OAI33xp33_ASAP7_75t_L g791 ( .A1(n_380), .A2(n_792), .A3(n_793), .B1(n_798), .B2(n_803), .B3(n_806), .Y(n_791) );
CKINVDCx8_ASAP7_75t_R g380 ( .A(n_381), .Y(n_380) );
INVx5_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx6_ASAP7_75t_L g624 ( .A(n_382), .Y(n_624) );
OR2x6_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g1122 ( .A(n_383), .B(n_395), .Y(n_1122) );
INVx2_ASAP7_75t_L g1004 ( .A(n_384), .Y(n_1004) );
NAND2x1p5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
AOI21xp33_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_405), .B(n_406), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_388), .A2(n_672), .B1(n_725), .B2(n_751), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_388), .A2(n_869), .B1(n_870), .B2(n_887), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_388), .A2(n_869), .B1(n_911), .B2(n_931), .Y(n_910) );
INVx5_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g511 ( .A(n_389), .Y(n_511) );
INVx1_ASAP7_75t_L g831 ( .A(n_389), .Y(n_831) );
INVx2_ASAP7_75t_L g1068 ( .A(n_389), .Y(n_1068) );
INVx2_ASAP7_75t_SL g1544 ( .A(n_389), .Y(n_1544) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx2_ASAP7_75t_L g703 ( .A(n_390), .Y(n_703) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x6_ASAP7_75t_L g1150 ( .A(n_392), .B(n_1151), .Y(n_1150) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_393), .B(n_416), .Y(n_1143) );
INVx2_ASAP7_75t_L g585 ( .A(n_394), .Y(n_585) );
AND2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_400), .Y(n_394) );
AND2x4_ASAP7_75t_L g433 ( .A(n_395), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g438 ( .A(n_395), .B(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g457 ( .A(n_395), .Y(n_457) );
AND2x2_ASAP7_75t_L g518 ( .A(n_395), .B(n_439), .Y(n_518) );
BUFx2_ASAP7_75t_L g656 ( .A(n_395), .Y(n_656) );
AND2x4_ASAP7_75t_L g669 ( .A(n_395), .B(n_434), .Y(n_669) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_395), .B(n_439), .Y(n_1219) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g416 ( .A(n_398), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g449 ( .A(n_399), .B(n_417), .Y(n_449) );
INVx6_ASAP7_75t_L g414 ( .A(n_400), .Y(n_414) );
BUFx2_ASAP7_75t_L g823 ( .A(n_400), .Y(n_823) );
INVx2_ASAP7_75t_L g1057 ( .A(n_400), .Y(n_1057) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g440 ( .A(n_401), .Y(n_440) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g411 ( .A(n_402), .B(n_404), .Y(n_411) );
AND2x4_ASAP7_75t_L g422 ( .A(n_402), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g436 ( .A(n_403), .Y(n_436) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g426 ( .A(n_404), .B(n_427), .Y(n_426) );
AOI31xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_441), .A3(n_458), .B(n_467), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g1034 ( .A1(n_409), .A2(n_429), .B(n_1035), .C(n_1036), .Y(n_1034) );
BUFx2_ASAP7_75t_L g1223 ( .A(n_409), .Y(n_1223) );
BUFx4f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g454 ( .A(n_410), .B(n_429), .Y(n_454) );
BUFx3_ASAP7_75t_L g566 ( .A(n_410), .Y(n_566) );
INVx2_ASAP7_75t_SL g576 ( .A(n_410), .Y(n_576) );
AND2x4_ASAP7_75t_L g927 ( .A(n_410), .B(n_656), .Y(n_927) );
BUFx6f_ASAP7_75t_L g1136 ( .A(n_410), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_411), .Y(n_446) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g745 ( .A(n_413), .Y(n_745) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
INVx1_ASAP7_75t_L g545 ( .A(n_414), .Y(n_545) );
INVx2_ASAP7_75t_L g736 ( .A(n_414), .Y(n_736) );
INVx2_ASAP7_75t_SL g820 ( .A(n_414), .Y(n_820) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_414), .Y(n_926) );
INVx1_ASAP7_75t_L g1139 ( .A(n_414), .Y(n_1139) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g531 ( .A(n_416), .Y(n_531) );
INVx2_ASAP7_75t_SL g648 ( .A(n_416), .Y(n_648) );
INVx1_ASAP7_75t_L g824 ( .A(n_416), .Y(n_824) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g1141 ( .A(n_420), .Y(n_1141) );
INVx2_ASAP7_75t_SL g420 ( .A(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g428 ( .A(n_421), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g521 ( .A(n_421), .Y(n_521) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx2_ASAP7_75t_L g443 ( .A(n_422), .Y(n_443) );
INVx2_ASAP7_75t_SL g537 ( .A(n_422), .Y(n_537) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_422), .Y(n_569) );
BUFx6f_ASAP7_75t_L g573 ( .A(n_422), .Y(n_573) );
BUFx6f_ASAP7_75t_L g664 ( .A(n_422), .Y(n_664) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_422), .Y(n_945) );
BUFx2_ASAP7_75t_L g953 ( .A(n_422), .Y(n_953) );
BUFx3_ASAP7_75t_L g1026 ( .A(n_422), .Y(n_1026) );
INVx1_ASAP7_75t_L g463 ( .A(n_423), .Y(n_463) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g564 ( .A(n_425), .Y(n_564) );
BUFx3_ASAP7_75t_L g641 ( .A(n_425), .Y(n_641) );
INVx1_ASAP7_75t_L g661 ( .A(n_425), .Y(n_661) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g466 ( .A(n_426), .Y(n_466) );
INVx1_ASAP7_75t_L g523 ( .A(n_426), .Y(n_523) );
BUFx6f_ASAP7_75t_L g548 ( .A(n_426), .Y(n_548) );
INVx1_ASAP7_75t_L g1103 ( .A(n_426), .Y(n_1103) );
INVx1_ASAP7_75t_L g462 ( .A(n_427), .Y(n_462) );
AOI211xp5_ASAP7_75t_L g514 ( .A1(n_428), .A2(n_504), .B(n_515), .C(n_519), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_428), .A2(n_459), .B1(n_578), .B2(n_579), .Y(n_577) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_428), .A2(n_459), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_428), .A2(n_459), .B1(n_848), .B2(n_854), .Y(n_885) );
AOI21xp33_ASAP7_75t_L g912 ( .A1(n_428), .A2(n_913), .B(n_914), .Y(n_912) );
HB1xp67_ASAP7_75t_L g1209 ( .A(n_428), .Y(n_1209) );
OAI21xp33_ASAP7_75t_L g657 ( .A1(n_429), .A2(n_658), .B(n_662), .Y(n_657) );
AND2x2_ASAP7_75t_L g814 ( .A(n_429), .B(n_664), .Y(n_814) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_429), .A2(n_459), .B1(n_948), .B2(n_949), .C(n_955), .Y(n_947) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g460 ( .A(n_430), .B(n_461), .Y(n_460) );
OR2x2_ASAP7_75t_L g465 ( .A(n_430), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g516 ( .A(n_433), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g582 ( .A1(n_433), .A2(n_518), .B1(n_583), .B2(n_584), .C1(n_586), .C2(n_587), .Y(n_582) );
AOI322xp5_ASAP7_75t_L g876 ( .A1(n_433), .A2(n_518), .A3(n_877), .B1(n_879), .B2(n_881), .C1(n_883), .C2(n_884), .Y(n_876) );
INVx2_ASAP7_75t_SL g1217 ( .A(n_433), .Y(n_1217) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g1120 ( .A(n_435), .Y(n_1120) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_SL g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_438), .A2(n_667), .B1(n_670), .B2(n_671), .Y(n_666) );
INVx2_ASAP7_75t_L g829 ( .A(n_438), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_438), .A2(n_669), .B1(n_990), .B2(n_991), .Y(n_1039) );
INVx2_ASAP7_75t_L g1126 ( .A(n_439), .Y(n_1126) );
BUFx3_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AND2x4_ASAP7_75t_L g455 ( .A(n_445), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g654 ( .A(n_445), .Y(n_654) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g541 ( .A(n_446), .Y(n_541) );
BUFx6f_ASAP7_75t_L g1540 ( .A(n_446), .Y(n_1540) );
INVx3_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g570 ( .A(n_448), .Y(n_570) );
BUFx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g542 ( .A(n_449), .Y(n_542) );
INVx2_ASAP7_75t_SL g742 ( .A(n_449), .Y(n_742) );
INVx2_ASAP7_75t_L g1130 ( .A(n_449), .Y(n_1130) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g651 ( .A(n_452), .Y(n_651) );
INVx2_ASAP7_75t_L g1227 ( .A(n_452), .Y(n_1227) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g534 ( .A(n_454), .Y(n_534) );
INVx1_ASAP7_75t_L g581 ( .A(n_454), .Y(n_581) );
INVx2_ASAP7_75t_SL g739 ( .A(n_454), .Y(n_739) );
INVx1_ASAP7_75t_L g873 ( .A(n_454), .Y(n_873) );
AOI221xp5_ASAP7_75t_L g1538 ( .A1(n_454), .A2(n_927), .B1(n_1531), .B2(n_1539), .C(n_1541), .Y(n_1538) );
AOI221xp5_ASAP7_75t_L g532 ( .A1(n_455), .A2(n_509), .B1(n_533), .B2(n_535), .C(n_543), .Y(n_532) );
INVx1_ASAP7_75t_L g588 ( .A(n_455), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g737 ( .A1(n_455), .A2(n_738), .B1(n_740), .B2(n_741), .C(n_743), .Y(n_737) );
AOI221xp5_ASAP7_75t_L g815 ( .A1(n_455), .A2(n_738), .B1(n_808), .B2(n_816), .C(n_817), .Y(n_815) );
AOI221xp5_ASAP7_75t_L g871 ( .A1(n_455), .A2(n_851), .B1(n_872), .B2(n_874), .C(n_875), .Y(n_871) );
AOI221xp5_ASAP7_75t_L g1220 ( .A1(n_455), .A2(n_872), .B1(n_1221), .B2(n_1222), .C(n_1225), .Y(n_1220) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_459), .A2(n_464), .B1(n_502), .B2(n_508), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g811 ( .A1(n_459), .A2(n_804), .B1(n_807), .B2(n_812), .Y(n_811) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_459), .A2(n_464), .B1(n_929), .B2(n_930), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1050 ( .A1(n_459), .A2(n_814), .B1(n_1051), .B2(n_1052), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1229 ( .A1(n_459), .A2(n_464), .B1(n_1230), .B2(n_1231), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1543 ( .A1(n_459), .A2(n_464), .B1(n_1525), .B2(n_1530), .Y(n_1543) );
INVx6_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g529 ( .A(n_461), .Y(n_529) );
INVx2_ASAP7_75t_L g660 ( .A(n_461), .Y(n_660) );
BUFx2_ASAP7_75t_L g1214 ( .A(n_461), .Y(n_1214) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x2_ASAP7_75t_L g527 ( .A(n_462), .B(n_463), .Y(n_527) );
AOI211xp5_ASAP7_75t_L g726 ( .A1(n_464), .A2(n_727), .B(n_728), .C(n_729), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_464), .A2(n_805), .B1(n_822), .B2(n_825), .C(n_827), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g886 ( .A(n_464), .B(n_857), .Y(n_886) );
AOI221xp5_ASAP7_75t_L g1053 ( .A1(n_464), .A2(n_1054), .B1(n_1055), .B2(n_1059), .C(n_1060), .Y(n_1053) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g826 ( .A(n_466), .Y(n_826) );
INVx2_ASAP7_75t_L g1024 ( .A(n_466), .Y(n_1024) );
INVx5_ASAP7_75t_L g589 ( .A(n_467), .Y(n_589) );
BUFx8_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g869 ( .A(n_468), .Y(n_869) );
OAI31xp33_ASAP7_75t_L g1157 ( .A1(n_468), .A2(n_1158), .A3(n_1175), .B(n_1195), .Y(n_1157) );
AOI31xp33_ASAP7_75t_L g1206 ( .A1(n_468), .A2(n_1207), .A3(n_1220), .B(n_1229), .Y(n_1206) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g672 ( .A(n_469), .Y(n_672) );
INVx1_ASAP7_75t_L g555 ( .A(n_471), .Y(n_555) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_510), .Y(n_471) );
NOR3xp33_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .C(n_485), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g965 ( .A1(n_476), .A2(n_703), .B1(n_966), .B2(n_967), .Y(n_965) );
OAI221xp5_ASAP7_75t_L g524 ( .A1(n_477), .A2(n_479), .B1(n_525), .B2(n_528), .C(n_530), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g505 ( .A1(n_488), .A2(n_506), .B1(n_508), .B2(n_509), .Y(n_505) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_495), .B1(n_496), .B2(n_499), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OAI22xp33_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_503), .B2(n_504), .Y(n_500) );
INVx1_ASAP7_75t_L g795 ( .A(n_501), .Y(n_795) );
INVx1_ASAP7_75t_L g845 ( .A(n_501), .Y(n_845) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B(n_513), .Y(n_510) );
AOI31xp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_532), .A3(n_549), .B(n_550), .Y(n_513) );
INVx2_ASAP7_75t_SL g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g732 ( .A(n_523), .Y(n_732) );
INVx1_ASAP7_75t_L g1228 ( .A(n_523), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_525), .A2(n_568), .B1(n_637), .B2(n_638), .C(n_639), .Y(n_636) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g665 ( .A(n_526), .Y(n_665) );
BUFx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx4f_ASAP7_75t_L g644 ( .A(n_527), .Y(n_644) );
INVx1_ASAP7_75t_L g951 ( .A(n_527), .Y(n_951) );
INVx2_ASAP7_75t_L g1029 ( .A(n_527), .Y(n_1029) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_528), .A2(n_643), .B1(n_645), .B2(n_646), .C(n_647), .Y(n_642) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OAI221xp5_ASAP7_75t_L g1212 ( .A1(n_530), .A2(n_1021), .B1(n_1213), .B2(n_1214), .C(n_1215), .Y(n_1212) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g882 ( .A(n_531), .Y(n_882) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g878 ( .A(n_537), .Y(n_878) );
INVx1_ASAP7_75t_L g1063 ( .A(n_537), .Y(n_1063) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g639 ( .A(n_542), .Y(n_639) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g634 ( .A(n_545), .Y(n_634) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_548), .Y(n_635) );
INVx2_ASAP7_75t_L g747 ( .A(n_548), .Y(n_747) );
BUFx6f_ASAP7_75t_L g1542 ( .A(n_548), .Y(n_1542) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g1532 ( .A1(n_551), .A2(n_1533), .B1(n_1544), .B2(n_1545), .Y(n_1532) );
CKINVDCx8_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
BUFx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g600 ( .A(n_553), .B(n_601), .Y(n_600) );
AND2x4_ASAP7_75t_L g757 ( .A(n_553), .B(n_601), .Y(n_757) );
AND2x2_ASAP7_75t_L g1003 ( .A(n_553), .B(n_1004), .Y(n_1003) );
OR2x6_ASAP7_75t_L g1129 ( .A(n_553), .B(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1152 ( .A(n_553), .Y(n_1152) );
INVx1_ASAP7_75t_L g716 ( .A(n_556), .Y(n_716) );
XNOR2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_629), .Y(n_556) );
INVx2_ASAP7_75t_SL g628 ( .A(n_558), .Y(n_628) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_590), .Y(n_558) );
OAI21xp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_580), .B(n_589), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .B1(n_571), .B2(n_574), .Y(n_561) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g731 ( .A(n_573), .Y(n_731) );
INVx1_ASAP7_75t_L g1037 ( .A(n_573), .Y(n_1037) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g880 ( .A(n_576), .Y(n_880) );
INVx2_ASAP7_75t_L g922 ( .A(n_576), .Y(n_922) );
INVx1_ASAP7_75t_L g1058 ( .A(n_576), .Y(n_1058) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_578), .A2(n_620), .B1(n_622), .B2(n_623), .Y(n_619) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_589), .A2(n_810), .B1(n_830), .B2(n_831), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_608), .Y(n_590) );
BUFx3_ASAP7_75t_L g769 ( .A(n_598), .Y(n_769) );
INVx1_ASAP7_75t_L g1193 ( .A(n_601), .Y(n_1193) );
OAI22xp33_ASAP7_75t_L g1514 ( .A1(n_603), .A2(n_1515), .B1(n_1516), .B2(n_1517), .Y(n_1514) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_604), .Y(n_1083) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g806 ( .A1(n_606), .A2(n_794), .B1(n_807), .B2(n_808), .Y(n_806) );
OAI22xp33_ASAP7_75t_L g1092 ( .A1(n_606), .A2(n_1051), .B1(n_1066), .B2(n_1083), .Y(n_1092) );
OAI22xp33_ASAP7_75t_L g1251 ( .A1(n_606), .A2(n_1167), .B1(n_1221), .B2(n_1231), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_613), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_612), .A2(n_652), .B1(n_702), .B2(n_703), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_624), .B1(n_625), .B2(n_626), .Y(n_613) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_618), .A2(n_638), .B1(n_683), .B2(n_686), .Y(n_682) );
INVx3_ASAP7_75t_L g692 ( .A(n_618), .Y(n_692) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g678 ( .A(n_621), .Y(n_678) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_623), .A2(n_678), .B1(n_695), .B2(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g697 ( .A(n_624), .Y(n_697) );
AOI33xp33_ASAP7_75t_L g756 ( .A1(n_624), .A2(n_757), .A3(n_758), .B1(n_764), .B2(n_765), .B3(n_768), .Y(n_756) );
AOI33xp33_ASAP7_75t_L g901 ( .A1(n_624), .A2(n_902), .A3(n_903), .B1(n_905), .B2(n_906), .B3(n_907), .Y(n_901) );
AOI222xp33_ASAP7_75t_L g968 ( .A1(n_624), .A2(n_757), .B1(n_969), .B2(n_971), .C1(n_972), .C2(n_980), .Y(n_968) );
INVx1_ASAP7_75t_L g1252 ( .A(n_624), .Y(n_1252) );
NAND4xp25_ASAP7_75t_L g630 ( .A(n_631), .B(n_673), .C(n_698), .D(n_704), .Y(n_630) );
OAI31xp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_640), .A3(n_649), .B(n_672), .Y(n_631) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_SL g954 ( .A(n_635), .Y(n_954) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_637), .A2(n_677), .B1(n_678), .B2(n_679), .Y(n_676) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
INVx2_ASAP7_75t_L g916 ( .A(n_644), .Y(n_916) );
INVx1_ASAP7_75t_L g1021 ( .A(n_644), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g673 ( .A1(n_646), .A2(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_650), .B(n_657), .C(n_666), .Y(n_649) );
A2O1A1Ixp33_ASAP7_75t_SL g650 ( .A1(n_651), .A2(n_652), .B(n_653), .C(n_655), .Y(n_650) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI21xp5_ASAP7_75t_SL g733 ( .A1(n_665), .A2(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx4_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g828 ( .A(n_669), .Y(n_828) );
INVx1_ASAP7_75t_SL g956 ( .A(n_669), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g704 ( .A1(n_670), .A2(n_671), .B1(n_705), .B2(n_710), .C(n_714), .Y(n_704) );
INVx2_ASAP7_75t_L g957 ( .A(n_672), .Y(n_957) );
OAI31xp33_ASAP7_75t_L g1016 ( .A1(n_672), .A2(n_1017), .A3(n_1018), .B(n_1033), .Y(n_1016) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_681), .B(n_1155), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1518 ( .A1(n_683), .A2(n_1519), .B1(n_1520), .B2(n_1521), .Y(n_1518) );
BUFx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx2_ASAP7_75t_L g800 ( .A(n_685), .Y(n_800) );
HB1xp67_ASAP7_75t_L g1247 ( .A(n_685), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_690), .B1(n_691), .B2(n_693), .Y(n_687) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_688), .Y(n_1180) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g853 ( .A(n_689), .Y(n_853) );
INVx2_ASAP7_75t_L g1524 ( .A(n_689), .Y(n_1524) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_701), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_703), .A2(n_1013), .B1(n_1014), .B2(n_1015), .Y(n_1012) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_707), .A2(n_712), .B1(n_714), .B2(n_754), .C(n_755), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_707), .A2(n_712), .B1(n_714), .B2(n_893), .C(n_894), .Y(n_892) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_707), .A2(n_712), .B1(n_714), .B2(n_960), .C(n_961), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_707), .A2(n_712), .B1(n_714), .B2(n_990), .C(n_991), .Y(n_989) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_713), .B(n_1154), .Y(n_1172) );
OAI22xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_720), .B1(n_934), .B2(n_935), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
XNOR2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_832), .Y(n_720) );
XOR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_779), .Y(n_721) );
XNOR2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_778), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_752), .Y(n_723) );
NAND3xp33_ASAP7_75t_SL g725 ( .A(n_726), .B(n_737), .C(n_748), .Y(n_725) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g923 ( .A(n_731), .Y(n_923) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g1065 ( .A(n_739), .Y(n_1065) );
BUFx2_ASAP7_75t_L g1224 ( .A(n_742), .Y(n_1224) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AND4x1_ASAP7_75t_L g752 ( .A(n_753), .B(n_756), .C(n_772), .D(n_774), .Y(n_752) );
BUFx2_ASAP7_75t_L g902 ( .A(n_757), .Y(n_902) );
AOI33xp33_ASAP7_75t_L g992 ( .A1(n_757), .A2(n_993), .A3(n_998), .B1(n_1000), .B2(n_1002), .B3(n_1003), .Y(n_992) );
HB1xp67_ASAP7_75t_L g904 ( .A(n_759), .Y(n_904) );
INVx1_ASAP7_75t_L g909 ( .A(n_759), .Y(n_909) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g995 ( .A(n_760), .Y(n_995) );
INVx2_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1091 ( .A1(n_767), .A2(n_1052), .B1(n_1054), .B2(n_1088), .Y(n_1091) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
XNOR2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_809), .Y(n_781) );
NOR3xp33_ASAP7_75t_L g782 ( .A(n_783), .B(n_790), .C(n_791), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_784), .B(n_787), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g847 ( .A1(n_794), .A2(n_848), .B1(n_849), .B2(n_851), .Y(n_847) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND3xp33_ASAP7_75t_L g810 ( .A(n_811), .B(n_815), .C(n_821), .Y(n_810) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g1534 ( .A1(n_814), .A2(n_1523), .B1(n_1535), .B2(n_1536), .C(n_1537), .Y(n_1534) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_889), .B1(n_932), .B2(n_933), .Y(n_832) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_834), .Y(n_933) );
INVx1_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_868), .Y(n_836) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_838), .B(n_858), .C(n_860), .Y(n_837) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
OAI22xp33_ASAP7_75t_L g1082 ( .A1(n_849), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_854), .B1(n_855), .B2(n_857), .Y(n_852) );
INVx2_ASAP7_75t_L g1166 ( .A(n_853), .Y(n_1166) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_861), .B(n_865), .Y(n_860) );
AOI22xp5_ASAP7_75t_L g1048 ( .A1(n_869), .A2(n_1049), .B1(n_1067), .B2(n_1068), .Y(n_1048) );
NAND4xp25_ASAP7_75t_L g870 ( .A(n_871), .B(n_876), .C(n_885), .D(n_886), .Y(n_870) );
AOI221xp5_ASAP7_75t_L g919 ( .A1(n_872), .A2(n_920), .B1(n_921), .B2(n_924), .C(n_927), .Y(n_919) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
AND2x2_ASAP7_75t_L g1114 ( .A(n_878), .B(n_1112), .Y(n_1114) );
INVx1_ASAP7_75t_L g932 ( .A(n_889), .Y(n_932) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_910), .Y(n_890) );
AND4x1_ASAP7_75t_L g891 ( .A(n_892), .B(n_895), .C(n_898), .D(n_901), .Y(n_891) );
OAI211xp5_ASAP7_75t_L g915 ( .A1(n_897), .A2(n_916), .B(n_917), .C(n_918), .Y(n_915) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_919), .C(n_928), .Y(n_911) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g941 ( .A1(n_927), .A2(n_942), .B1(n_943), .B2(n_944), .C(n_946), .Y(n_941) );
INVx1_ASAP7_75t_L g1032 ( .A(n_927), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g1061 ( .A1(n_927), .A2(n_1062), .B1(n_1064), .B2(n_1065), .C(n_1066), .Y(n_1061) );
INVxp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
HB1xp67_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
XNOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_986), .Y(n_937) );
NOR2x1_ASAP7_75t_L g939 ( .A(n_940), .B(n_958), .Y(n_939) );
AOI21xp5_ASAP7_75t_L g940 ( .A1(n_941), .A2(n_947), .B(n_957), .Y(n_940) );
HB1xp67_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
NAND4xp25_ASAP7_75t_L g958 ( .A(n_959), .B(n_962), .C(n_965), .D(n_968), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g1509 ( .A1(n_969), .A2(n_1009), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_970), .B(n_1154), .Y(n_1153) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g1090 ( .A(n_975), .Y(n_1090) );
INVx2_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g1521 ( .A(n_983), .Y(n_1521) );
NAND3xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_1007), .C(n_1016), .Y(n_987) );
AND3x1_ASAP7_75t_L g988 ( .A(n_989), .B(n_992), .C(n_1005), .Y(n_988) );
INVx2_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
INVx2_ASAP7_75t_SL g1169 ( .A(n_1004), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1012), .Y(n_1007) );
OAI211xp5_ASAP7_75t_L g1027 ( .A1(n_1011), .A2(n_1028), .B(n_1030), .C(n_1031), .Y(n_1027) );
AOI22xp5_ASAP7_75t_L g1505 ( .A1(n_1013), .A2(n_1506), .B1(n_1507), .B2(n_1508), .Y(n_1505) );
NAND3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1027), .C(n_1032), .Y(n_1018) );
OAI211xp5_ASAP7_75t_L g1019 ( .A1(n_1020), .A2(n_1021), .B(n_1022), .C(n_1025), .Y(n_1019) );
BUFx2_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx2_ASAP7_75t_L g1038 ( .A(n_1024), .Y(n_1038) );
BUFx3_ASAP7_75t_L g1132 ( .A(n_1026), .Y(n_1132) );
BUFx3_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
OR2x6_ASAP7_75t_L g1107 ( .A(n_1029), .B(n_1104), .Y(n_1107) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1038), .Y(n_1211) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1043), .B1(n_1200), .B2(n_1254), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
XNOR2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1093), .Y(n_1043) );
INVx1_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_1048), .B(n_1069), .Y(n_1047) );
NAND3xp33_ASAP7_75t_SL g1049 ( .A(n_1050), .B(n_1053), .C(n_1061), .Y(n_1049) );
INVx1_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_1057), .Y(n_1111) );
AOI21xp5_ASAP7_75t_L g1204 ( .A1(n_1068), .A2(n_1205), .B(n_1206), .Y(n_1204) );
NOR3xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1078), .C(n_1081), .Y(n_1069) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_1071), .B(n_1075), .Y(n_1070) );
HB1xp67_ASAP7_75t_L g1240 ( .A(n_1080), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1088), .B1(n_1089), .B2(n_1090), .Y(n_1086) );
INVx1_ASAP7_75t_L g1093 ( .A(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
AND3x1_ASAP7_75t_L g1096 ( .A(n_1097), .B(n_1148), .C(n_1157), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1115), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1098 ( .A(n_1099), .B(n_1108), .Y(n_1098) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1101), .B1(n_1105), .B2(n_1106), .Y(n_1099) );
OAI221xp5_ASAP7_75t_L g1164 ( .A1(n_1100), .A2(n_1113), .B1(n_1165), .B2(n_1167), .C(n_1168), .Y(n_1164) );
CKINVDCx6p67_ASAP7_75t_R g1101 ( .A(n_1102), .Y(n_1101) );
OR2x6_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1104), .Y(n_1102) );
INVx2_ASAP7_75t_L g1133 ( .A(n_1103), .Y(n_1133) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1104), .Y(n_1112) );
CKINVDCx6p67_ASAP7_75t_R g1106 ( .A(n_1107), .Y(n_1106) );
AOI22xp33_ASAP7_75t_L g1108 ( .A1(n_1109), .A2(n_1110), .B1(n_1113), .B2(n_1114), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
NAND3xp33_ASAP7_75t_SL g1115 ( .A(n_1116), .B(n_1127), .C(n_1144), .Y(n_1115) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_1117), .A2(n_1118), .B1(n_1123), .B2(n_1124), .Y(n_1116) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_1117), .A2(n_1123), .B1(n_1171), .B2(n_1173), .Y(n_1170) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
NAND2x1p5_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1121), .Y(n_1119) );
INVx2_ASAP7_75t_SL g1121 ( .A(n_1122), .Y(n_1121) );
OR2x6_ASAP7_75t_L g1125 ( .A(n_1122), .B(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1122), .Y(n_1147) );
INVx2_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
AOI33xp33_ASAP7_75t_L g1127 ( .A1(n_1128), .A2(n_1131), .A3(n_1134), .B1(n_1137), .B2(n_1140), .B3(n_1142), .Y(n_1127) );
CKINVDCx5p33_ASAP7_75t_R g1128 ( .A(n_1129), .Y(n_1128) );
HB1xp67_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1136), .B(n_1147), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
BUFx4f_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
NAND2xp5_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
NOR2xp67_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx8_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
AND2x4_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1163), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1199 ( .A(n_1161), .B(n_1185), .Y(n_1199) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_1167), .A2(n_1246), .B1(n_1248), .B2(n_1249), .Y(n_1245) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
CKINVDCx11_ASAP7_75t_R g1173 ( .A(n_1174), .Y(n_1173) );
CKINVDCx6p67_ASAP7_75t_R g1176 ( .A(n_1177), .Y(n_1176) );
OAI22xp5_ASAP7_75t_SL g1178 ( .A1(n_1179), .A2(n_1180), .B1(n_1181), .B2(n_1182), .Y(n_1178) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1186), .Y(n_1528) );
BUFx3_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx3_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx3_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_SL g1200 ( .A(n_1201), .Y(n_1200) );
HB1xp67_ASAP7_75t_L g1254 ( .A(n_1201), .Y(n_1254) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1204), .B(n_1232), .Y(n_1203) );
AOI211xp5_ASAP7_75t_L g1207 ( .A1(n_1208), .A2(n_1209), .B(n_1210), .C(n_1216), .Y(n_1207) );
INVx3_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
HB1xp67_ASAP7_75t_L g1226 ( .A(n_1227), .Y(n_1226) );
NOR3xp33_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1239), .C(n_1241), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1234), .B(n_1236), .Y(n_1233) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1247), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_1253), .A2(n_1278), .B1(n_1279), .B2(n_1284), .Y(n_1277) );
OAI221xp5_ASAP7_75t_SL g1256 ( .A1(n_1257), .A2(n_1497), .B1(n_1499), .B2(n_1546), .C(n_1552), .Y(n_1256) );
AND5x1_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1407), .C(n_1445), .D(n_1457), .E(n_1480), .Y(n_1257) );
A2O1A1Ixp33_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1261), .B(n_1349), .C(n_1383), .Y(n_1258) );
OAI211xp5_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1295), .B(n_1336), .C(n_1338), .Y(n_1259) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1286), .Y(n_1260) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1261), .Y(n_1347) );
INVx3_ASAP7_75t_L g1369 ( .A(n_1261), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1261), .B(n_1328), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1381 ( .A(n_1261), .B(n_1382), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1261), .B(n_1393), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1261), .B(n_1286), .Y(n_1439) );
INVx3_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1348 ( .A(n_1262), .B(n_1286), .Y(n_1348) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1262), .B(n_1372), .Y(n_1371) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1277), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1263 ( .A1(n_1264), .A2(n_1265), .B1(n_1272), .B2(n_1273), .Y(n_1263) );
OAI22xp5_ASAP7_75t_L g1317 ( .A1(n_1265), .A2(n_1275), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
OAI22xp33_ASAP7_75t_L g1330 ( .A1(n_1265), .A2(n_1275), .B1(n_1331), .B2(n_1332), .Y(n_1330) );
BUFx3_ASAP7_75t_L g1365 ( .A(n_1265), .Y(n_1365) );
BUFx6f_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_1266), .A2(n_1275), .B1(n_1303), .B2(n_1304), .Y(n_1302) );
OR2x2_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1268), .Y(n_1266) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1267), .B(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1267), .Y(n_1290) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1268), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1271), .Y(n_1268) );
HB1xp67_ASAP7_75t_L g1568 ( .A(n_1269), .Y(n_1568) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1271), .Y(n_1282) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_1273), .Y(n_1367) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1276), .Y(n_1292) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1280), .Y(n_1279) );
INVx1_ASAP7_75t_L g1361 ( .A(n_1280), .Y(n_1361) );
AND2x4_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1283), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1281), .B(n_1283), .Y(n_1294) );
HB1xp67_ASAP7_75t_L g1566 ( .A(n_1281), .Y(n_1566) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
AND2x4_ASAP7_75t_L g1285 ( .A(n_1282), .B(n_1283), .Y(n_1285) );
OAI22xp5_ASAP7_75t_L g1313 ( .A1(n_1284), .A2(n_1314), .B1(n_1315), .B2(n_1316), .Y(n_1313) );
INVx1_ASAP7_75t_SL g1284 ( .A(n_1285), .Y(n_1284) );
INVx2_ASAP7_75t_L g1310 ( .A(n_1285), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1344 ( .A(n_1286), .B(n_1328), .Y(n_1344) );
OR2x2_ASAP7_75t_L g1355 ( .A(n_1286), .B(n_1328), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1372 ( .A(n_1286), .B(n_1329), .Y(n_1372) );
INVx2_ASAP7_75t_L g1382 ( .A(n_1286), .Y(n_1382) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1286), .B(n_1329), .Y(n_1393) );
OAI211xp5_ASAP7_75t_L g1421 ( .A1(n_1286), .A2(n_1422), .B(n_1424), .C(n_1427), .Y(n_1421) );
OAI221xp5_ASAP7_75t_L g1447 ( .A1(n_1286), .A2(n_1336), .B1(n_1448), .B2(n_1450), .C(n_1451), .Y(n_1447) );
OAI211xp5_ASAP7_75t_L g1459 ( .A1(n_1286), .A2(n_1460), .B(n_1462), .C(n_1468), .Y(n_1459) );
AND2x4_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1293), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1290), .Y(n_1288) );
AND2x4_ASAP7_75t_L g1291 ( .A(n_1290), .B(n_1292), .Y(n_1291) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1294), .Y(n_1314) );
AOI211xp5_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1305), .B(n_1320), .C(n_1323), .Y(n_1295) );
AOI21xp33_ASAP7_75t_L g1401 ( .A1(n_1296), .A2(n_1402), .B(n_1404), .Y(n_1401) );
AOI21xp5_ASAP7_75t_L g1455 ( .A1(n_1296), .A2(n_1404), .B(n_1441), .Y(n_1455) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1297), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1297), .B(n_1321), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1297), .B(n_1311), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1409 ( .A(n_1297), .B(n_1305), .Y(n_1409) );
NAND2xp5_ASAP7_75t_L g1419 ( .A(n_1297), .B(n_1306), .Y(n_1419) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1301), .Y(n_1297) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_1298), .B(n_1301), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1298), .B(n_1335), .Y(n_1334) );
NOR2xp33_ASAP7_75t_L g1342 ( .A(n_1298), .B(n_1343), .Y(n_1342) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1298), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1298), .B(n_1312), .Y(n_1454) );
AND2x2_ASAP7_75t_L g1298 ( .A(n_1299), .B(n_1300), .Y(n_1298) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1301), .Y(n_1335) );
AND2x2_ASAP7_75t_L g1376 ( .A(n_1301), .B(n_1377), .Y(n_1376) );
AND2x2_ASAP7_75t_L g1392 ( .A(n_1301), .B(n_1311), .Y(n_1392) );
NOR2xp33_ASAP7_75t_L g1403 ( .A(n_1301), .B(n_1311), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1301), .B(n_1305), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1305), .B(n_1376), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1413 ( .A(n_1305), .B(n_1414), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1311), .Y(n_1305) );
INVx4_ASAP7_75t_L g1321 ( .A(n_1306), .Y(n_1321) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1306), .Y(n_1325) );
OR2x2_ASAP7_75t_L g1336 ( .A(n_1306), .B(n_1337), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1390 ( .A(n_1306), .B(n_1322), .Y(n_1390) );
OR2x2_ASAP7_75t_L g1444 ( .A(n_1306), .B(n_1326), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1460 ( .A(n_1306), .B(n_1461), .Y(n_1460) );
NOR2xp33_ASAP7_75t_L g1471 ( .A(n_1306), .B(n_1311), .Y(n_1471) );
AND2x6_ASAP7_75t_L g1306 ( .A(n_1307), .B(n_1308), .Y(n_1306) );
INVx2_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1359 ( .A1(n_1310), .A2(n_1360), .B1(n_1361), .B2(n_1362), .Y(n_1359) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1310), .Y(n_1498) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1311), .B(n_1335), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1374 ( .A(n_1311), .B(n_1335), .Y(n_1374) );
NOR2xp33_ASAP7_75t_L g1418 ( .A(n_1311), .B(n_1419), .Y(n_1418) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1311), .B(n_1376), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1311), .B(n_1353), .Y(n_1449) );
CKINVDCx6p67_ASAP7_75t_R g1311 ( .A(n_1312), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1312), .B(n_1322), .Y(n_1337) );
NAND2xp5_ASAP7_75t_L g1352 ( .A(n_1312), .B(n_1353), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1312), .B(n_1377), .Y(n_1400) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1312), .B(n_1376), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1442 ( .A(n_1312), .B(n_1414), .Y(n_1442) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1312), .B(n_1334), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1479 ( .A(n_1312), .B(n_1377), .Y(n_1479) );
OR2x6_ASAP7_75t_SL g1312 ( .A(n_1313), .B(n_1317), .Y(n_1312) );
NOR2xp33_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1322), .Y(n_1320) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1321), .B(n_1344), .Y(n_1343) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1321), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1321), .B(n_1429), .Y(n_1428) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1321), .B(n_1479), .Y(n_1485) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1322), .Y(n_1414) );
NOR2xp33_ASAP7_75t_L g1323 ( .A(n_1324), .B(n_1333), .Y(n_1323) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1324), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1326), .Y(n_1324) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1325), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1325), .B(n_1392), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1398 ( .A(n_1325), .B(n_1399), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1325), .B(n_1423), .Y(n_1422) );
OAI21xp33_ASAP7_75t_L g1440 ( .A1(n_1325), .A2(n_1402), .B(n_1441), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1325), .B(n_1454), .Y(n_1453) );
NOR2xp33_ASAP7_75t_L g1465 ( .A(n_1325), .B(n_1382), .Y(n_1465) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1327), .Y(n_1346) );
O2A1O1Ixp33_ASAP7_75t_L g1396 ( .A1(n_1327), .A2(n_1397), .B(n_1398), .C(n_1401), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g1477 ( .A(n_1327), .B(n_1478), .Y(n_1477) );
INVx2_ASAP7_75t_SL g1327 ( .A(n_1328), .Y(n_1327) );
INVx2_ASAP7_75t_SL g1328 ( .A(n_1329), .Y(n_1328) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_1329), .Y(n_1412) );
NOR2xp33_ASAP7_75t_L g1435 ( .A(n_1333), .B(n_1436), .Y(n_1435) );
NOR3xp33_ASAP7_75t_L g1443 ( .A(n_1333), .B(n_1369), .C(n_1444), .Y(n_1443) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OAI222xp33_ASAP7_75t_L g1370 ( .A1(n_1337), .A2(n_1371), .B1(n_1373), .B2(n_1375), .C1(n_1378), .C2(n_1380), .Y(n_1370) );
NOR2xp33_ASAP7_75t_L g1456 ( .A(n_1337), .B(n_1371), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1338 ( .A1(n_1339), .A2(n_1342), .B1(n_1345), .B2(n_1348), .Y(n_1338) );
NOR2x1_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1341), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1340), .B(n_1479), .Y(n_1478) );
NOR2x1_ASAP7_75t_R g1491 ( .A(n_1340), .B(n_1492), .Y(n_1491) );
OR2x2_ASAP7_75t_L g1496 ( .A(n_1340), .B(n_1355), .Y(n_1496) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_1344), .A2(n_1389), .B1(n_1391), .B2(n_1393), .C(n_1394), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1344), .B(n_1395), .Y(n_1394) );
A2O1A1Ixp33_ASAP7_75t_L g1451 ( .A1(n_1344), .A2(n_1358), .B(n_1452), .C(n_1455), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1347), .Y(n_1345) );
O2A1O1Ixp33_ASAP7_75t_SL g1407 ( .A1(n_1347), .A2(n_1408), .B(n_1421), .C(n_1430), .Y(n_1407) );
INVxp67_ASAP7_75t_SL g1349 ( .A(n_1350), .Y(n_1349) );
OAI211xp5_ASAP7_75t_L g1383 ( .A1(n_1350), .A2(n_1384), .B(n_1388), .C(n_1396), .Y(n_1383) );
AOI21xp5_ASAP7_75t_L g1350 ( .A1(n_1351), .A2(n_1368), .B(n_1370), .Y(n_1350) );
OAI21xp5_ASAP7_75t_SL g1351 ( .A1(n_1352), .A2(n_1354), .B(n_1356), .Y(n_1351) );
OAI21xp5_ASAP7_75t_SL g1415 ( .A1(n_1354), .A2(n_1416), .B(n_1420), .Y(n_1415) );
OAI21xp33_ASAP7_75t_SL g1431 ( .A1(n_1354), .A2(n_1432), .B(n_1433), .Y(n_1431) );
INVx2_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
NOR2xp33_ASAP7_75t_L g1466 ( .A(n_1355), .B(n_1467), .Y(n_1466) );
CKINVDCx14_ASAP7_75t_R g1356 ( .A(n_1357), .Y(n_1356) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1368 ( .A(n_1358), .B(n_1369), .Y(n_1368) );
CKINVDCx5p33_ASAP7_75t_R g1386 ( .A(n_1358), .Y(n_1386) );
AOI31xp33_ASAP7_75t_L g1430 ( .A1(n_1358), .A2(n_1431), .A3(n_1434), .B(n_1438), .Y(n_1430) );
OR2x6_ASAP7_75t_SL g1358 ( .A(n_1359), .B(n_1363), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1365), .B1(n_1366), .B2(n_1367), .Y(n_1363) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1368), .Y(n_1458) );
INVx1_ASAP7_75t_SL g1387 ( .A(n_1369), .Y(n_1387) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1371), .Y(n_1446) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1372), .Y(n_1429) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1374), .B(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1395 ( .A(n_1375), .Y(n_1395) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1376), .Y(n_1492) );
INVx1_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
AOI221xp5_ASAP7_75t_L g1438 ( .A1(n_1379), .A2(n_1398), .B1(n_1439), .B2(n_1440), .C(n_1443), .Y(n_1438) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1381), .Y(n_1380) );
AOI21xp5_ASAP7_75t_L g1434 ( .A1(n_1381), .A2(n_1397), .B(n_1435), .Y(n_1434) );
NOR2xp33_ASAP7_75t_L g1450 ( .A(n_1381), .B(n_1412), .Y(n_1450) );
A2O1A1Ixp33_ASAP7_75t_L g1408 ( .A1(n_1382), .A2(n_1409), .B(n_1410), .C(n_1415), .Y(n_1408) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1382), .B(n_1386), .Y(n_1476) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1387), .Y(n_1385) );
OAI21xp33_ASAP7_75t_L g1483 ( .A1(n_1386), .A2(n_1412), .B(n_1484), .Y(n_1483) );
AOI21xp5_ASAP7_75t_L g1490 ( .A1(n_1386), .A2(n_1429), .B(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1391), .Y(n_1487) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1393), .B(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1489 ( .A(n_1393), .Y(n_1489) );
INVx1_ASAP7_75t_L g1488 ( .A(n_1398), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_1399), .B(n_1423), .Y(n_1464) );
INVx1_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
AND2x2_ASAP7_75t_L g1473 ( .A(n_1409), .B(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1410), .Y(n_1481) );
OR2x2_ASAP7_75t_L g1410 ( .A(n_1411), .B(n_1413), .Y(n_1410) );
OAI21xp33_ASAP7_75t_L g1468 ( .A1(n_1411), .A2(n_1469), .B(n_1472), .Y(n_1468) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1412), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1470 ( .A(n_1414), .B(n_1471), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1494 ( .A(n_1414), .B(n_1495), .Y(n_1494) );
AOI211xp5_ASAP7_75t_L g1445 ( .A1(n_1416), .A2(n_1446), .B(n_1447), .C(n_1456), .Y(n_1445) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1422), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1425 ( .A(n_1423), .B(n_1426), .Y(n_1425) );
INVxp67_ASAP7_75t_L g1424 ( .A(n_1425), .Y(n_1424) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1449), .Y(n_1448) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
AOI22xp5_ASAP7_75t_L g1457 ( .A1(n_1458), .A2(n_1459), .B1(n_1475), .B2(n_1477), .Y(n_1457) );
INVx1_ASAP7_75t_L g1482 ( .A(n_1460), .Y(n_1482) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1461), .Y(n_1467) );
AOI21xp5_ASAP7_75t_L g1462 ( .A1(n_1463), .A2(n_1465), .B(n_1466), .Y(n_1462) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1469 ( .A(n_1470), .Y(n_1469) );
INVxp67_ASAP7_75t_SL g1472 ( .A(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
OAI321xp33_ASAP7_75t_L g1480 ( .A1(n_1476), .A2(n_1481), .A3(n_1482), .B1(n_1483), .B2(n_1486), .C(n_1493), .Y(n_1480) );
INVxp33_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
A2O1A1Ixp33_ASAP7_75t_L g1486 ( .A1(n_1487), .A2(n_1488), .B(n_1489), .C(n_1490), .Y(n_1486) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx1_ASAP7_75t_L g1495 ( .A(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1498), .Y(n_1497) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
XNOR2x1_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1502), .Y(n_1500) );
HB1xp67_ASAP7_75t_L g1560 ( .A(n_1502), .Y(n_1560) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1503), .B(n_1532), .Y(n_1502) );
NOR3xp33_ASAP7_75t_L g1503 ( .A(n_1504), .B(n_1512), .C(n_1513), .Y(n_1503) );
NAND2xp5_ASAP7_75t_L g1504 ( .A(n_1505), .B(n_1509), .Y(n_1504) );
OAI22xp5_ASAP7_75t_SL g1522 ( .A1(n_1523), .A2(n_1524), .B1(n_1525), .B2(n_1526), .Y(n_1522) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
HB1xp67_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
NAND3xp33_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1538), .C(n_1543), .Y(n_1533) );
INVx1_ASAP7_75t_SL g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
CKINVDCx5p33_ASAP7_75t_R g1554 ( .A(n_1555), .Y(n_1554) );
A2O1A1Ixp33_ASAP7_75t_L g1564 ( .A1(n_1556), .A2(n_1565), .B(n_1567), .C(n_1569), .Y(n_1564) );
INVxp33_ASAP7_75t_SL g1557 ( .A(n_1558), .Y(n_1557) );
INVx1_ASAP7_75t_L g1561 ( .A(n_1560), .Y(n_1561) );
BUFx2_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
HB1xp67_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
endmodule