module fake_jpeg_25292_n_324 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_324);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_324;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_44),
.Y(n_48)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_47),
.A2(n_63),
.B1(n_40),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_44),
.A2(n_25),
.B1(n_17),
.B2(n_27),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_60),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_58),
.Y(n_74)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_64),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_41),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_67),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_53),
.B1(n_57),
.B2(n_64),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_51),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_41),
.B1(n_35),
.B2(n_40),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_85),
.B1(n_21),
.B2(n_22),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_77),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_53),
.A2(n_38),
.B1(n_43),
.B2(n_40),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_76),
.B(n_87),
.Y(n_95)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_54),
.B(n_20),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_79),
.B(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_46),
.B(n_18),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_43),
.B1(n_26),
.B2(n_24),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_31),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_43),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_61),
.B(n_20),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_89),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_43),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_39),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_43),
.B1(n_33),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_23),
.B1(n_31),
.B2(n_30),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_33),
.B1(n_60),
.B2(n_56),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_108),
.B1(n_113),
.B2(n_120),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_24),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_87),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_68),
.B(n_61),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_122),
.B(n_87),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_37),
.C(n_39),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_91),
.C(n_88),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_111),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_108)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_76),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_121),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_81),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_117),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_72),
.A2(n_33),
.B1(n_19),
.B2(n_23),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_80),
.A2(n_30),
.B1(n_39),
.B2(n_36),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_124),
.B1(n_151),
.B2(n_115),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_80),
.B1(n_70),
.B2(n_73),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_131),
.B(n_143),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_128),
.B(n_138),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_129),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_96),
.B(n_82),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_132),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_95),
.A2(n_89),
.B(n_79),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_101),
.Y(n_132)
);

AO21x1_ASAP7_75t_SL g134 ( 
.A1(n_108),
.A2(n_76),
.B(n_87),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_120),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_100),
.B(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_152),
.Y(n_163)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_86),
.A3(n_84),
.B1(n_83),
.B2(n_76),
.Y(n_137)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_91),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_104),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_139),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_142),
.C(n_16),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_76),
.B(n_92),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_148),
.B(n_117),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_75),
.C(n_55),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_100),
.A2(n_77),
.B(n_93),
.C(n_74),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_95),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_146),
.B1(n_149),
.B2(n_144),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_99),
.A2(n_102),
.B1(n_122),
.B2(n_113),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_19),
.B(n_16),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_74),
.B1(n_93),
.B2(n_30),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_36),
.B1(n_39),
.B2(n_37),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_155),
.B(n_159),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_165),
.B1(n_136),
.B2(n_146),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_158),
.B(n_162),
.Y(n_191)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_110),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_168),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_167),
.A2(n_169),
.B1(n_183),
.B2(n_0),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_110),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_112),
.B1(n_103),
.B2(n_105),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_172),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_103),
.B1(n_109),
.B2(n_96),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_171),
.A2(n_173),
.B1(n_131),
.B2(n_148),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_145),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_123),
.A2(n_109),
.B1(n_98),
.B2(n_118),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_174),
.B(n_175),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_115),
.B(n_118),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_126),
.B(n_1),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_125),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_177),
.B(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_138),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_129),
.B(n_121),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_181),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_127),
.B(n_140),
.C(n_142),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_136),
.A2(n_114),
.B1(n_36),
.B2(n_37),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_184),
.Y(n_188)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_214),
.C(n_155),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_189),
.A2(n_194),
.B1(n_199),
.B2(n_200),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_190),
.B(n_212),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_133),
.B1(n_130),
.B2(n_134),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_192),
.A2(n_203),
.B1(n_208),
.B2(n_7),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_170),
.A2(n_151),
.B1(n_128),
.B2(n_126),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_197),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_198),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_36),
.B1(n_37),
.B2(n_16),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_154),
.A2(n_37),
.B1(n_16),
.B2(n_19),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_185),
.A2(n_37),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_213),
.B1(n_183),
.B2(n_167),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_8),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_168),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g213 ( 
.A1(n_157),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_9),
.C(n_14),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_213),
.A2(n_184),
.B1(n_164),
.B2(n_161),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_227),
.B1(n_231),
.B2(n_203),
.Y(n_241)
);

AO22x1_ASAP7_75t_L g216 ( 
.A1(n_207),
.A2(n_158),
.B1(n_163),
.B2(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_221),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_179),
.B(n_182),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_SL g253 ( 
.A(n_218),
.B(n_222),
.C(n_225),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_202),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_206),
.B(n_153),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_190),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_226),
.C(n_232),
.Y(n_242)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_229),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_179),
.B(n_163),
.Y(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_193),
.A2(n_174),
.B1(n_169),
.B2(n_159),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_209),
.B(n_176),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_234),
.C(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_9),
.C(n_14),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_238),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_188),
.Y(n_239)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_193),
.B(n_204),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_240),
.B(n_247),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_199),
.B1(n_201),
.B2(n_200),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_188),
.Y(n_244)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_254),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_187),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_216),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_187),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_227),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_213),
.B(n_2),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_223),
.C(n_233),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_220),
.B1(n_231),
.B2(n_225),
.Y(n_261)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_261),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_259),
.C(n_249),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_265),
.C(n_273),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_226),
.C(n_211),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_267),
.A2(n_270),
.B1(n_255),
.B2(n_248),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_222),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_253),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_243),
.A2(n_220),
.B1(n_234),
.B2(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_218),
.B1(n_213),
.B2(n_196),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_232),
.C(n_197),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_213),
.C(n_9),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_274),
.B(n_252),
.C(n_245),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_240),
.B(n_243),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_279),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_285),
.B1(n_278),
.B2(n_262),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_274),
.B(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_283),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_271),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_289),
.C(n_270),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_250),
.C(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_280),
.C(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_287),
.Y(n_299)
);

NAND2xp33_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_7),
.Y(n_288)
);

OAI321xp33_ASAP7_75t_L g298 ( 
.A1(n_288),
.A2(n_10),
.A3(n_15),
.B1(n_13),
.B2(n_12),
.C(n_11),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_7),
.B(n_13),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_261),
.Y(n_291)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_291),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_292),
.A2(n_298),
.B(n_4),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_263),
.C(n_272),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_3),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_260),
.C(n_268),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_267),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_279),
.B1(n_287),
.B2(n_15),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_302),
.A2(n_309),
.B1(n_306),
.B2(n_290),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_SL g303 ( 
.A(n_293),
.B(n_10),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_306),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_296),
.B(n_1),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_310),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_4),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_297),
.Y(n_312)
);

BUFx24_ASAP7_75t_SL g317 ( 
.A(n_312),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_299),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_299),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_314),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_311),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_311),
.B1(n_319),
.B2(n_315),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_316),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_322),
.B(n_4),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_5),
.B(n_6),
.Y(n_324)
);


endmodule