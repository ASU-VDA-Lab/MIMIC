module fake_netlist_1_6506_n_659 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_659);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_659;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_387;
wire n_476;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_616;
wire n_365;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_187;
wire n_375;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
BUFx2_ASAP7_75t_L g183 ( .A(n_117), .Y(n_183) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_85), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_118), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_100), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_103), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g189 ( .A(n_141), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_64), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_40), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_1), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_72), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g194 ( .A(n_99), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_6), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_131), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g197 ( .A(n_157), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_150), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_97), .Y(n_199) );
INVxp67_ASAP7_75t_SL g200 ( .A(n_142), .Y(n_200) );
BUFx3_ASAP7_75t_L g201 ( .A(n_12), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_110), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_91), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_127), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_36), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_177), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_106), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_82), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_89), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_29), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_169), .B(n_2), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_95), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_134), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_71), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_39), .Y(n_216) );
INVx1_ASAP7_75t_SL g217 ( .A(n_138), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_56), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g219 ( .A(n_43), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_90), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_135), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_11), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_172), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_144), .Y(n_225) );
BUFx3_ASAP7_75t_L g226 ( .A(n_146), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_137), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_18), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_96), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_139), .Y(n_230) );
INVxp67_ASAP7_75t_L g231 ( .A(n_125), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_111), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_87), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_54), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_109), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_70), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_94), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_16), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_101), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_115), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_152), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_163), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_18), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_107), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_86), .Y(n_245) );
INVxp33_ASAP7_75t_SL g246 ( .A(n_128), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_143), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_30), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_116), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_57), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_46), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_92), .Y(n_252) );
CKINVDCx14_ASAP7_75t_R g253 ( .A(n_168), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_98), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_102), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_173), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_108), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_105), .Y(n_258) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_174), .Y(n_259) );
NOR2xp67_ASAP7_75t_L g260 ( .A(n_84), .B(n_30), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_145), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_149), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_56), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_133), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_59), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_121), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_130), .Y(n_267) );
INVxp33_ASAP7_75t_SL g268 ( .A(n_93), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_77), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_171), .Y(n_270) );
BUFx2_ASAP7_75t_L g271 ( .A(n_123), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_129), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_58), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_136), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_57), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_122), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_49), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_11), .Y(n_278) );
CKINVDCx14_ASAP7_75t_R g279 ( .A(n_79), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_51), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_52), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_104), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_73), .Y(n_283) );
INVxp67_ASAP7_75t_SL g284 ( .A(n_80), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_36), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_166), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_37), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_0), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_182), .Y(n_289) );
INVxp33_ASAP7_75t_SL g290 ( .A(n_42), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_8), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_154), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_51), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_183), .B(n_0), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_271), .B(n_1), .Y(n_295) );
AND2x4_ASAP7_75t_L g296 ( .A(n_288), .B(n_3), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_237), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g298 ( .A1(n_290), .A2(n_5), .B1(n_3), .B2(n_4), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_237), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_237), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_237), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_201), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_215), .B(n_4), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_185), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_185), .Y(n_305) );
AND2x6_ASAP7_75t_L g306 ( .A(n_205), .B(n_74), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_290), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_308) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_219), .A2(n_10), .B1(n_7), .B2(n_9), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_233), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_215), .B(n_10), .Y(n_311) );
INVxp67_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_205), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_293), .B(n_12), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_233), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_239), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_201), .Y(n_317) );
BUFx3_ASAP7_75t_L g318 ( .A(n_226), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_190), .B(n_13), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_243), .B(n_13), .Y(n_320) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_236), .Y(n_321) );
OR2x6_ASAP7_75t_L g322 ( .A(n_260), .B(n_75), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_184), .B(n_14), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_236), .Y(n_324) );
BUFx2_ASAP7_75t_L g325 ( .A(n_280), .Y(n_325) );
INVxp33_ASAP7_75t_SL g326 ( .A(n_193), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_280), .Y(n_327) );
AND2x4_ASAP7_75t_L g328 ( .A(n_239), .B(n_14), .Y(n_328) );
AND2x4_ASAP7_75t_L g329 ( .A(n_270), .B(n_15), .Y(n_329) );
BUFx3_ASAP7_75t_L g330 ( .A(n_313), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
INVx4_ASAP7_75t_L g332 ( .A(n_322), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g333 ( .A1(n_296), .A2(n_192), .B1(n_195), .B2(n_191), .Y(n_333) );
BUFx10_ASAP7_75t_L g334 ( .A(n_294), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_313), .Y(n_337) );
INVx4_ASAP7_75t_L g338 ( .A(n_322), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_305), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_322), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_325), .B(n_270), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_325), .B(n_274), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_328), .B(n_274), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_300), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_328), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_321), .B(n_194), .Y(n_350) );
INVx6_ASAP7_75t_L g351 ( .A(n_328), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g352 ( .A(n_321), .B(n_207), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_310), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_312), .B(n_242), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g355 ( .A(n_312), .B(n_259), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_295), .B(n_253), .Y(n_356) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_300), .Y(n_357) );
INVx4_ASAP7_75t_L g358 ( .A(n_322), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_302), .B(n_317), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_315), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_302), .B(n_276), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_302), .B(n_286), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_315), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_302), .B(n_286), .Y(n_365) );
INVx5_ASAP7_75t_L g366 ( .A(n_306), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_317), .B(n_187), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_316), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_326), .B(n_231), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_300), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_332), .A2(n_294), .B1(n_329), .B2(n_328), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_356), .B(n_295), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_331), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_351), .Y(n_375) );
NAND2x1_ASAP7_75t_L g376 ( .A(n_351), .B(n_322), .Y(n_376) );
NAND2xp5_ASAP7_75t_SL g377 ( .A(n_332), .B(n_294), .Y(n_377) );
INVx2_ASAP7_75t_SL g378 ( .A(n_356), .Y(n_378) );
OR2x6_ASAP7_75t_L g379 ( .A(n_350), .B(n_323), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_352), .B(n_345), .Y(n_380) );
NAND2xp5_ASAP7_75t_SL g381 ( .A(n_332), .B(n_294), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_352), .B(n_323), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_345), .B(n_303), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_338), .A2(n_329), .B1(n_296), .B2(n_311), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_338), .B(n_329), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_336), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g387 ( .A(n_338), .B(n_296), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_342), .B(n_296), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_346), .B(n_318), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_342), .A2(n_311), .B1(n_303), .B2(n_317), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
NAND2xp5_ASAP7_75t_SL g392 ( .A(n_342), .B(n_318), .Y(n_392) );
INVxp67_ASAP7_75t_L g393 ( .A(n_369), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_354), .A2(n_320), .B1(n_309), .B2(n_186), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_333), .B(n_317), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_367), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_333), .B(n_327), .Y(n_397) );
NAND2xp5_ASAP7_75t_SL g398 ( .A(n_358), .B(n_188), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_349), .B(n_324), .Y(n_399) );
AND2x4_ASAP7_75t_L g400 ( .A(n_358), .B(n_314), .Y(n_400) );
AND2x4_ASAP7_75t_L g401 ( .A(n_358), .B(n_314), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_349), .B(n_189), .Y(n_402) );
NAND3xp33_ASAP7_75t_L g403 ( .A(n_355), .B(n_308), .C(n_298), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_347), .B(n_319), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_334), .A2(n_319), .B1(n_268), .B2(n_246), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_340), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_367), .B(n_211), .Y(n_407) );
INVx4_ASAP7_75t_L g408 ( .A(n_334), .Y(n_408) );
NAND2x1p5_ASAP7_75t_L g409 ( .A(n_366), .B(n_298), .Y(n_409) );
BUFx8_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_353), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_353), .Y(n_412) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_362), .A2(n_186), .B1(n_214), .B2(n_208), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_330), .B(n_196), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_335), .B(n_307), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_337), .B(n_197), .Y(n_416) );
NAND2xp5_ASAP7_75t_SL g417 ( .A(n_366), .B(n_198), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_337), .B(n_199), .Y(n_418) );
A2O1A1Ixp33_ASAP7_75t_SL g419 ( .A1(n_360), .A2(n_316), .B(n_279), .C(n_204), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_360), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_363), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_361), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
NOR2xp33_ASAP7_75t_SL g424 ( .A(n_366), .B(n_208), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_337), .B(n_199), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_368), .A2(n_306), .B1(n_206), .B2(n_218), .Y(n_426) );
CKINVDCx5p33_ASAP7_75t_R g427 ( .A(n_363), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_368), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_365), .B(n_223), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_359), .B(n_209), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_393), .B(n_308), .Y(n_431) );
NOR2x1_ASAP7_75t_L g432 ( .A(n_400), .B(n_212), .Y(n_432) );
OR2x6_ASAP7_75t_L g433 ( .A(n_379), .B(n_216), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_377), .A2(n_366), .B(n_284), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_383), .B(n_265), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_408), .Y(n_436) );
INVx5_ASAP7_75t_L g437 ( .A(n_379), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_374), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_382), .A2(n_234), .B(n_238), .C(n_228), .Y(n_439) );
AND2x6_ASAP7_75t_L g440 ( .A(n_400), .B(n_226), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_L g441 ( .A1(n_372), .A2(n_250), .B(n_251), .C(n_248), .Y(n_441) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_404), .A2(n_316), .B(n_263), .C(n_273), .Y(n_442) );
O2A1O1Ixp33_ASAP7_75t_SL g443 ( .A1(n_419), .A2(n_210), .B(n_213), .C(n_203), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_429), .B(n_221), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_407), .B(n_227), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_377), .A2(n_200), .B(n_341), .Y(n_446) );
O2A1O1Ixp33_ASAP7_75t_SL g447 ( .A1(n_419), .A2(n_222), .B(n_224), .C(n_220), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_410), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_401), .B(n_229), .Y(n_449) );
O2A1O1Ixp5_ASAP7_75t_SL g450 ( .A1(n_385), .A2(n_230), .B(n_232), .C(n_225), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_405), .B(n_257), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_386), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_371), .A2(n_277), .B(n_278), .C(n_275), .Y(n_453) );
AND2x4_ASAP7_75t_L g454 ( .A(n_381), .B(n_387), .Y(n_454) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_384), .A2(n_285), .B(n_287), .C(n_283), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_394), .B(n_291), .Y(n_456) );
NOR2xp33_ASAP7_75t_R g457 ( .A(n_424), .B(n_262), .Y(n_457) );
A2O1A1Ixp33_ASAP7_75t_L g458 ( .A1(n_395), .A2(n_240), .B(n_241), .C(n_235), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_387), .A2(n_306), .B1(n_245), .B2(n_247), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_413), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g461 ( .A1(n_409), .A2(n_388), .B1(n_397), .B2(n_375), .Y(n_461) );
OAI21xp33_ASAP7_75t_L g462 ( .A1(n_430), .A2(n_269), .B(n_264), .Y(n_462) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_391), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_406), .B(n_282), .Y(n_464) );
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_415), .A2(n_299), .B(n_301), .C(n_297), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_415), .A2(n_249), .B(n_252), .C(n_244), .Y(n_466) );
OAI21x1_ASAP7_75t_L g467 ( .A1(n_392), .A2(n_348), .B(n_343), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_422), .B(n_289), .Y(n_468) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_411), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_412), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_SL g471 ( .A1(n_390), .A2(n_299), .B(n_301), .C(n_297), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_389), .B(n_292), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_428), .A2(n_255), .B1(n_256), .B2(n_254), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_402), .B(n_15), .Y(n_474) );
OAI21xp33_ASAP7_75t_L g475 ( .A1(n_414), .A2(n_217), .B(n_202), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_399), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_398), .A2(n_370), .B(n_261), .Y(n_477) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_420), .A2(n_258), .B1(n_267), .B2(n_266), .Y(n_478) );
AND2x6_ASAP7_75t_L g479 ( .A(n_423), .B(n_272), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_416), .A2(n_301), .B(n_297), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_418), .B(n_357), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_425), .A2(n_357), .B(n_76), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_426), .B(n_17), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_417), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_417), .A2(n_22), .B1(n_23), .B2(n_24), .Y(n_485) );
AOI21x1_ASAP7_75t_L g486 ( .A1(n_376), .A2(n_357), .B(n_78), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_379), .B(n_23), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g488 ( .A1(n_380), .A2(n_25), .B(n_26), .C(n_27), .Y(n_488) );
BUFx6f_ASAP7_75t_L g489 ( .A(n_408), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_421), .A2(n_27), .B1(n_28), .B2(n_29), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_393), .B(n_31), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_379), .B(n_32), .Y(n_492) );
BUFx4f_ASAP7_75t_L g493 ( .A(n_379), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_396), .B(n_32), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g495 ( .A1(n_421), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_377), .A2(n_357), .B(n_81), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_380), .A2(n_33), .B(n_34), .C(n_37), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_378), .B(n_38), .Y(n_498) );
O2A1O1Ixp5_ASAP7_75t_L g499 ( .A1(n_486), .A2(n_120), .B(n_181), .C(n_180), .Y(n_499) );
O2A1O1Ixp33_ASAP7_75t_SL g500 ( .A1(n_471), .A2(n_119), .B(n_179), .C(n_178), .Y(n_500) );
AO31x2_ASAP7_75t_L g501 ( .A1(n_458), .A2(n_41), .A3(n_44), .B(n_45), .Y(n_501) );
AO21x1_ASAP7_75t_L g502 ( .A1(n_488), .A2(n_88), .B(n_83), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_460), .A2(n_46), .B1(n_47), .B2(n_48), .Y(n_503) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_481), .A2(n_124), .B(n_176), .C(n_175), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_489), .B(n_493), .Y(n_505) );
AO31x2_ASAP7_75t_L g506 ( .A1(n_466), .A2(n_48), .A3(n_49), .B(n_50), .Y(n_506) );
OR2x6_ASAP7_75t_L g507 ( .A(n_448), .B(n_50), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_476), .A2(n_53), .B(n_55), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
OAI21xp5_ASAP7_75t_L g510 ( .A1(n_450), .A2(n_132), .B(n_170), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_453), .A2(n_60), .B(n_61), .C(n_62), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_497), .A2(n_63), .B(n_65), .C(n_66), .Y(n_512) );
AO31x2_ASAP7_75t_L g513 ( .A1(n_496), .A2(n_65), .A3(n_67), .B(n_68), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_437), .B(n_69), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
O2A1O1Ixp33_ASAP7_75t_SL g516 ( .A1(n_452), .A2(n_112), .B(n_113), .C(n_114), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_435), .B(n_126), .Y(n_517) );
INVxp67_ASAP7_75t_SL g518 ( .A(n_463), .Y(n_518) );
AO31x2_ASAP7_75t_L g519 ( .A1(n_473), .A2(n_147), .A3(n_148), .B(n_151), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_487), .B(n_153), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_480), .A2(n_156), .B(n_158), .Y(n_521) );
AOI21xp33_ASAP7_75t_L g522 ( .A1(n_451), .A2(n_159), .B(n_160), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_474), .A2(n_161), .B(n_162), .C(n_165), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g524 ( .A(n_436), .B(n_167), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_445), .B(n_444), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_464), .B(n_454), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_454), .A2(n_492), .B1(n_432), .B2(n_440), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_494), .A2(n_475), .B(n_446), .C(n_477), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_443), .B(n_447), .C(n_461), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_434), .A2(n_472), .B(n_468), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_449), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_484), .A2(n_485), .B(n_483), .C(n_462), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_463), .A2(n_469), .B(n_470), .Y(n_533) );
AO31x2_ASAP7_75t_L g534 ( .A1(n_479), .A2(n_469), .A3(n_459), .B(n_457), .Y(n_534) );
NOR2xp33_ASAP7_75t_SL g535 ( .A(n_493), .B(n_410), .Y(n_535) );
AO32x2_ASAP7_75t_L g536 ( .A1(n_490), .A2(n_495), .A3(n_478), .B1(n_473), .B2(n_485), .Y(n_536) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_431), .A2(n_427), .B1(n_421), .B2(n_403), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g538 ( .A1(n_431), .A2(n_456), .B1(n_403), .B2(n_373), .C(n_393), .Y(n_538) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_467), .A2(n_482), .B(n_486), .Y(n_539) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_455), .A2(n_453), .B(n_442), .C(n_458), .Y(n_540) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_489), .Y(n_541) );
INVx5_ASAP7_75t_L g542 ( .A(n_489), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_439), .A2(n_441), .B(n_491), .C(n_404), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_SL g544 ( .A1(n_471), .A2(n_419), .B(n_465), .C(n_458), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_SL g545 ( .A1(n_471), .A2(n_419), .B(n_465), .C(n_458), .Y(n_545) );
A2O1A1Ixp33_ASAP7_75t_L g546 ( .A1(n_439), .A2(n_441), .B(n_491), .C(n_404), .Y(n_546) );
BUFx6f_ASAP7_75t_L g547 ( .A(n_541), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_507), .B(n_509), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_544), .A2(n_545), .B(n_539), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_515), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_538), .B(n_531), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_526), .B(n_525), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_533), .A2(n_500), .B(n_529), .Y(n_553) );
AO21x2_ASAP7_75t_L g554 ( .A1(n_510), .A2(n_529), .B(n_502), .Y(n_554) );
HB1xp67_ASAP7_75t_L g555 ( .A(n_542), .Y(n_555) );
INVx3_ASAP7_75t_L g556 ( .A(n_542), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_507), .Y(n_557) );
BUFx10_ASAP7_75t_L g558 ( .A(n_507), .Y(n_558) );
NAND2x1p5_ASAP7_75t_L g559 ( .A(n_505), .B(n_514), .Y(n_559) );
NOR2x1_ASAP7_75t_SL g560 ( .A(n_541), .B(n_535), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_501), .Y(n_561) );
OA21x2_ASAP7_75t_L g562 ( .A1(n_499), .A2(n_521), .B(n_504), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_508), .A2(n_503), .B1(n_520), .B2(n_524), .Y(n_563) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_508), .A2(n_522), .B(n_516), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_536), .B(n_506), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_534), .B(n_518), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_534), .B(n_511), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_536), .B(n_513), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_519), .Y(n_569) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_502), .A2(n_528), .A3(n_512), .B(n_523), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_537), .B(n_431), .Y(n_571) );
AOI21xp33_ASAP7_75t_L g572 ( .A1(n_532), .A2(n_529), .B(n_540), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_542), .B(n_448), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g576 ( .A1(n_527), .A2(n_537), .B1(n_498), .B2(n_427), .Y(n_576) );
AO31x2_ASAP7_75t_L g577 ( .A1(n_502), .A2(n_528), .A3(n_512), .B(n_523), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_578) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_502), .A2(n_528), .A3(n_512), .B(n_523), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_538), .B(n_531), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_538), .B(n_531), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g582 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_583) );
AOI21xp5_ASAP7_75t_L g584 ( .A1(n_530), .A2(n_528), .B(n_517), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_525), .A2(n_540), .B(n_546), .C(n_543), .Y(n_585) );
INVx5_ASAP7_75t_L g586 ( .A(n_547), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_551), .B(n_580), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_571), .B(n_550), .Y(n_588) );
OR2x6_ASAP7_75t_L g589 ( .A(n_548), .B(n_557), .Y(n_589) );
BUFx3_ASAP7_75t_L g590 ( .A(n_575), .Y(n_590) );
OR2x6_ASAP7_75t_L g591 ( .A(n_548), .B(n_559), .Y(n_591) );
AND2x6_ASAP7_75t_L g592 ( .A(n_566), .B(n_565), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_561), .Y(n_593) );
OA21x2_ASAP7_75t_L g594 ( .A1(n_573), .A2(n_578), .B(n_574), .Y(n_594) );
AOI21xp5_ASAP7_75t_SL g595 ( .A1(n_563), .A2(n_560), .B(n_585), .Y(n_595) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_555), .Y(n_596) );
OA21x2_ASAP7_75t_L g597 ( .A1(n_582), .A2(n_584), .B(n_583), .Y(n_597) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_549), .A2(n_572), .B(n_569), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_556), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_581), .B(n_568), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_552), .B(n_576), .Y(n_601) );
AO21x2_ASAP7_75t_L g602 ( .A1(n_572), .A2(n_553), .B(n_567), .Y(n_602) );
INVx5_ASAP7_75t_L g603 ( .A(n_558), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_564), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_570), .B(n_579), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_593), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_605), .B(n_577), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_605), .B(n_554), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_600), .B(n_562), .Y(n_609) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_595), .B(n_592), .Y(n_610) );
BUFx2_ASAP7_75t_L g611 ( .A(n_592), .Y(n_611) );
BUFx2_ASAP7_75t_L g612 ( .A(n_592), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_602), .B(n_588), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_601), .B(n_587), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_588), .B(n_598), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_613), .B(n_598), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_613), .B(n_604), .Y(n_617) );
NAND2x1p5_ASAP7_75t_L g618 ( .A(n_611), .B(n_603), .Y(n_618) );
INVx3_ASAP7_75t_L g619 ( .A(n_610), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_614), .B(n_596), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_607), .B(n_594), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_607), .B(n_594), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_607), .B(n_597), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_611), .B(n_603), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_606), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_625), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_621), .B(n_615), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_620), .B(n_615), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_622), .B(n_608), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_622), .B(n_608), .Y(n_630) );
NAND2x1_ASAP7_75t_L g631 ( .A(n_619), .B(n_612), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_623), .B(n_609), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_623), .B(n_609), .Y(n_633) );
OR2x2_ASAP7_75t_L g634 ( .A(n_628), .B(n_627), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_626), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_628), .B(n_617), .Y(n_636) );
NOR2xp67_ASAP7_75t_L g637 ( .A(n_632), .B(n_619), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_633), .B(n_616), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_635), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_638), .B(n_629), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_635), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_634), .B(n_630), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_637), .B(n_631), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_636), .B(n_617), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_639), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_641), .Y(n_646) );
NOR2x1p5_ASAP7_75t_L g647 ( .A(n_643), .B(n_642), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_647), .B(n_640), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_645), .B(n_644), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_649), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_648), .B(n_646), .Y(n_651) );
BUFx2_ASAP7_75t_L g652 ( .A(n_650), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_652), .B(n_651), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_653), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_654), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_655), .A2(n_589), .B1(n_591), .B2(n_590), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_656), .Y(n_657) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_657), .A2(n_599), .B(n_624), .C(n_618), .Y(n_658) );
AOI21xp5_ASAP7_75t_L g659 ( .A1(n_658), .A2(n_599), .B(n_586), .Y(n_659) );
endmodule