module fake_jpeg_29208_n_533 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_533);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_17),
.B(n_18),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_SL g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_SL g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_53),
.A2(n_30),
.B1(n_47),
.B2(n_46),
.Y(n_112)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_17),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_56),
.B(n_65),
.Y(n_103)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_57),
.Y(n_137)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_58),
.Y(n_155)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_60),
.Y(n_130)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_89),
.Y(n_102)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_63),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_64),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_26),
.B(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_67),
.Y(n_121)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

INVx11_ASAP7_75t_SL g71 ( 
.A(n_36),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_73),
.Y(n_148)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_85),
.Y(n_114)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_79),
.Y(n_128)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_26),
.B(n_15),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_87),
.Y(n_158)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_21),
.B(n_15),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_15),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_100),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_28),
.B(n_49),
.Y(n_97)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_98),
.Y(n_156)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_0),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_37),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_38),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_30),
.B1(n_45),
.B2(n_43),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_106),
.A2(n_120),
.B1(n_92),
.B2(n_67),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx13_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_55),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_115),
.B(n_123),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_59),
.B(n_24),
.C(n_40),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_119),
.B(n_33),
.C(n_86),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_88),
.A2(n_30),
.B1(n_45),
.B2(n_43),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_93),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_56),
.B(n_47),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_136),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_53),
.A2(n_49),
.B(n_28),
.C(n_40),
.Y(n_135)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_135),
.A2(n_86),
.B(n_63),
.C(n_60),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_46),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_83),
.B(n_38),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_72),
.B(n_37),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_73),
.Y(n_144)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_78),
.B(n_20),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_57),
.B(n_44),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_150),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_44),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_76),
.B(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_153),
.B(n_160),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_51),
.B(n_44),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_78),
.B(n_20),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_82),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_116),
.A2(n_36),
.B(n_40),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_L g256 ( 
.A1(n_165),
.A2(n_110),
.B(n_3),
.C(n_4),
.Y(n_256)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_166),
.Y(n_268)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_167),
.Y(n_230)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_154),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_168),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_105),
.B(n_102),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_133),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_172),
.B(n_178),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_98),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_175),
.B(n_201),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_112),
.A2(n_66),
.B1(n_64),
.B2(n_87),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_176),
.A2(n_159),
.B1(n_157),
.B2(n_151),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_114),
.B(n_74),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_179),
.B(n_191),
.Y(n_265)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_181),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_182),
.Y(n_249)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_109),
.Y(n_183)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_184),
.Y(n_275)
);

CKINVDCx12_ASAP7_75t_R g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_185),
.Y(n_271)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_187),
.Y(n_234)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_189),
.A2(n_195),
.B1(n_107),
.B2(n_154),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_190),
.B(n_210),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_113),
.B(n_76),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_192),
.Y(n_251)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_198),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_106),
.A2(n_58),
.B1(n_69),
.B2(n_23),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_199),
.Y(n_261)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_142),
.B(n_1),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_34),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_141),
.Y(n_203)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_203),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_130),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_204),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_108),
.B(n_50),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_208),
.Y(n_252)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

BUFx6f_ASAP7_75t_SL g247 ( 
.A(n_206),
.Y(n_247)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_104),
.B(n_96),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_135),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_209),
.B(n_225),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_156),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_45),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_213),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_128),
.A2(n_79),
.B1(n_75),
.B2(n_70),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_212),
.A2(n_120),
.B1(n_158),
.B2(n_128),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_125),
.B(n_43),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_214),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_215),
.B(n_14),
.Y(n_262)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_217),
.Y(n_239)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_219),
.Y(n_260)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_119),
.B(n_33),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_163),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_221),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_264)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_223),
.Y(n_263)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_155),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_224),
.B(n_7),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_158),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_231),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_229),
.A2(n_232),
.B1(n_236),
.B2(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_152),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_189),
.A2(n_152),
.B1(n_159),
.B2(n_157),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_237),
.A2(n_269),
.B1(n_203),
.B2(n_182),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_190),
.A2(n_134),
.B1(n_117),
.B2(n_132),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_132),
.C(n_121),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_250),
.C(n_262),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_177),
.B(n_161),
.C(n_134),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_175),
.A2(n_110),
.B1(n_163),
.B2(n_4),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_254),
.A2(n_222),
.B1(n_194),
.B2(n_200),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_259),
.B(n_168),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_258),
.B(n_167),
.Y(n_308)
);

AO22x2_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_264),
.A2(n_168),
.B1(n_172),
.B2(n_198),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_171),
.A2(n_14),
.B1(n_8),
.B2(n_9),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_174),
.B(n_180),
.C(n_170),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_183),
.C(n_217),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_276),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_165),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_277),
.B(n_287),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_279),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_281),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_201),
.B(n_210),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_282),
.A2(n_293),
.B(n_314),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_283),
.A2(n_12),
.B(n_13),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_168),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_284),
.B(n_291),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_263),
.Y(n_286)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_286),
.Y(n_333)
);

AND2x6_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_173),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_238),
.B(n_207),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_304),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_290),
.A2(n_299),
.B1(n_318),
.B2(n_286),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_228),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_241),
.B(n_252),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_292),
.B(n_297),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_274),
.A2(n_192),
.B(n_224),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_294),
.B(n_306),
.Y(n_336)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_230),
.Y(n_295)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_295),
.Y(n_338)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_262),
.B(n_227),
.CI(n_243),
.CON(n_297),
.SN(n_297)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_249),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_261),
.A2(n_184),
.B1(n_219),
.B2(n_181),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_300),
.A2(n_12),
.B1(n_13),
.B2(n_320),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g302 ( 
.A(n_228),
.Y(n_302)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_302),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_231),
.B(n_253),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_261),
.A2(n_204),
.B1(n_214),
.B2(n_257),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_305),
.A2(n_270),
.B1(n_249),
.B2(n_275),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_265),
.B(n_223),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_307),
.B(n_316),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_309),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_216),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_233),
.Y(n_310)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_310),
.Y(n_350)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_235),
.Y(n_311)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_311),
.Y(n_359)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_312),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_188),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_315),
.Y(n_342)
);

O2A1O1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_187),
.B(n_173),
.C(n_206),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_228),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_317),
.B(n_318),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_255),
.B(n_166),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_221),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_322),
.Y(n_361)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_242),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_323),
.Y(n_353)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_8),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_313),
.A2(n_302),
.B(n_277),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_326),
.B(n_282),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

AO21x2_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_259),
.B(n_232),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_331),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_280),
.B(n_272),
.C(n_267),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_334),
.C(n_343),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_226),
.C(n_251),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_293),
.A2(n_229),
.B(n_259),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_345),
.B(n_300),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_297),
.B(n_246),
.C(n_234),
.Y(n_343)
);

OAI32xp33_ASAP7_75t_L g344 ( 
.A1(n_303),
.A2(n_237),
.A3(n_270),
.B1(n_246),
.B2(n_234),
.Y(n_344)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_306),
.A2(n_247),
.B(n_268),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_301),
.A2(n_275),
.B1(n_248),
.B2(n_247),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_355),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_291),
.A2(n_248),
.B1(n_268),
.B2(n_11),
.Y(n_348)
);

BUFx8_ASAP7_75t_L g399 ( 
.A(n_348),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_8),
.C(n_9),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_358),
.Y(n_394)
);

NAND2xp33_ASAP7_75t_SL g389 ( 
.A(n_357),
.B(n_314),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_303),
.B(n_12),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_320),
.A2(n_12),
.B1(n_309),
.B2(n_308),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_360),
.B(n_323),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_364),
.A2(n_290),
.B1(n_287),
.B2(n_283),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_324),
.B(n_292),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_365),
.B(n_371),
.Y(n_428)
);

XNOR2x2_ASAP7_75t_SL g366 ( 
.A(n_342),
.B(n_304),
.Y(n_366)
);

OA21x2_ASAP7_75t_L g424 ( 
.A1(n_366),
.A2(n_331),
.B(n_338),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_367),
.A2(n_325),
.B(n_345),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_334),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_370),
.B(n_397),
.C(n_349),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_330),
.Y(n_373)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_373),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_374),
.A2(n_353),
.B1(n_335),
.B2(n_327),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_375),
.A2(n_338),
.B(n_340),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_352),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_376),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_363),
.B(n_289),
.Y(n_377)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_377),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_278),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_379),
.B(n_398),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_333),
.B(n_279),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_380),
.B(n_386),
.Y(n_405)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_362),
.Y(n_381)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_381),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_294),
.Y(n_382)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_382),
.Y(n_423)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_330),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_384),
.A2(n_395),
.B1(n_360),
.B2(n_355),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_333),
.B(n_321),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_288),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_387),
.B(n_388),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_329),
.B(n_281),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g425 ( 
.A(n_389),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_322),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

XOR2x2_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_299),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_391),
.B(n_384),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_354),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_392),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_354),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_393),
.B(n_396),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_337),
.A2(n_295),
.B1(n_296),
.B2(n_310),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_312),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_335),
.B(n_315),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_317),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_400),
.A2(n_410),
.B1(n_414),
.B2(n_369),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_370),
.B(n_326),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_401),
.B(n_407),
.Y(n_440)
);

AO22x1_ASAP7_75t_SL g402 ( 
.A1(n_369),
.A2(n_331),
.B1(n_344),
.B2(n_364),
.Y(n_402)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_402),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_404),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_408),
.B(n_371),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_332),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_409),
.B(n_411),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_368),
.A2(n_341),
.B1(n_339),
.B2(n_331),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_372),
.B(n_351),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_358),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_422),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_368),
.A2(n_341),
.B1(n_331),
.B2(n_349),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_367),
.B(n_325),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_427),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_347),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_395),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_415),
.A2(n_425),
.B(n_369),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_432),
.A2(n_433),
.B(n_431),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_416),
.A2(n_365),
.B1(n_385),
.B2(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_434),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_392),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g469 ( 
.A(n_436),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_438),
.A2(n_449),
.B1(n_450),
.B2(n_454),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_439),
.A2(n_448),
.B1(n_429),
.B2(n_407),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_400),
.A2(n_385),
.B1(n_378),
.B2(n_376),
.Y(n_441)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_442),
.B(n_446),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_417),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_443),
.B(n_444),
.Y(n_476)
);

OA22x2_ASAP7_75t_L g444 ( 
.A1(n_414),
.A2(n_391),
.B1(n_378),
.B2(n_366),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_402),
.Y(n_472)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_406),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_447),
.B(n_451),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_410),
.A2(n_398),
.B1(n_366),
.B2(n_378),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_405),
.A2(n_393),
.B1(n_373),
.B2(n_383),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_423),
.A2(n_399),
.B1(n_389),
.B2(n_381),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_413),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_427),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_425),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_418),
.A2(n_399),
.B1(n_340),
.B2(n_350),
.Y(n_454)
);

BUFx24_ASAP7_75t_SL g455 ( 
.A(n_411),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_455),
.B(n_394),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_443),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_457),
.B(n_474),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_458),
.A2(n_453),
.B1(n_438),
.B2(n_444),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_409),
.C(n_401),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_459),
.B(n_460),
.C(n_461),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_430),
.B(n_422),
.C(n_415),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_404),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_412),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_462),
.B(n_464),
.C(n_468),
.Y(n_485)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_463),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_431),
.C(n_445),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_424),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_SL g470 ( 
.A(n_433),
.B(n_435),
.Y(n_470)
);

OAI322xp33_ASAP7_75t_L g492 ( 
.A1(n_470),
.A2(n_475),
.A3(n_394),
.B1(n_444),
.B2(n_432),
.C1(n_359),
.C2(n_403),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_472),
.B(n_402),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_473),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_448),
.B(n_424),
.Y(n_474)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_476),
.Y(n_478)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_478),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_453),
.Y(n_479)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_479),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_456),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_482),
.B(n_490),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_484),
.A2(n_493),
.B1(n_420),
.B2(n_350),
.Y(n_505)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_476),
.Y(n_486)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_486),
.Y(n_504)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_465),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_489),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_488),
.B(n_491),
.Y(n_501)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_463),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_467),
.A2(n_439),
.B1(n_444),
.B2(n_426),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_473),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_492),
.Y(n_498)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

OAI21xp33_ASAP7_75t_L g494 ( 
.A1(n_480),
.A2(n_470),
.B(n_466),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_494),
.B(n_497),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_481),
.B(n_460),
.C(n_459),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_496),
.C(n_485),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_464),
.C(n_461),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_477),
.A2(n_472),
.B1(n_458),
.B2(n_468),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_478),
.A2(n_469),
.B1(n_399),
.B2(n_420),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_500),
.B(n_505),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_485),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_509),
.B(n_513),
.C(n_479),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_501),
.A2(n_487),
.B1(n_493),
.B2(n_491),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_510),
.B(n_514),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g518 ( 
.A(n_511),
.B(n_462),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_503),
.A2(n_489),
.B(n_477),
.Y(n_512)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_502),
.B(n_504),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_488),
.C(n_490),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_506),
.B(n_483),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_486),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_497),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_517),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_518),
.B(n_521),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_519),
.B(n_520),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_508),
.A2(n_498),
.B1(n_499),
.B2(n_479),
.Y(n_521)
);

NOR2x1_ASAP7_75t_L g523 ( 
.A(n_516),
.B(n_494),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_523),
.A2(n_516),
.B(n_507),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g528 ( 
.A1(n_526),
.A2(n_527),
.B(n_525),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_524),
.B(n_511),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_528),
.B(n_522),
.C(n_513),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_523),
.B1(n_508),
.B2(n_362),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_399),
.B(n_346),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_531),
.B(n_346),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_298),
.B(n_526),
.Y(n_533)
);


endmodule