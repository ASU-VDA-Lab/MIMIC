module fake_jpeg_7750_n_320 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_28),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_38),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_0),
.Y(n_37)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_37),
.B(n_41),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_46),
.Y(n_58)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_50),
.Y(n_80)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_60),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_32),
.B1(n_25),
.B2(n_29),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_53),
.A2(n_59),
.B(n_20),
.Y(n_93)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_22),
.B1(n_20),
.B2(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_29),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_38),
.Y(n_73)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_64),
.A2(n_69),
.B1(n_40),
.B2(n_41),
.Y(n_98)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_71),
.B(n_81),
.Y(n_107)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_94),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_46),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_84),
.B(n_88),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_85),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_38),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_40),
.B1(n_45),
.B2(n_22),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_39),
.B1(n_54),
.B2(n_56),
.Y(n_122)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_35),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_63),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_63),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_99),
.B(n_82),
.C(n_79),
.Y(n_132)
);

AO22x1_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_41),
.B1(n_63),
.B2(n_65),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_102),
.A2(n_123),
.B(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_121),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_19),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_97),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_110),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_122),
.B1(n_125),
.B2(n_90),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_39),
.A3(n_42),
.B1(n_19),
.B2(n_45),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_114),
.Y(n_147)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_113),
.B(n_33),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_39),
.A3(n_42),
.B1(n_45),
.B2(n_34),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_85),
.A2(n_45),
.B1(n_54),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_80),
.B1(n_76),
.B2(n_87),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_87),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_118),
.A2(n_72),
.B1(n_71),
.B2(n_86),
.Y(n_135)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_77),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_78),
.A2(n_56),
.B(n_54),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_50),
.B1(n_28),
.B2(n_17),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_34),
.B(n_24),
.Y(n_157)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_102),
.A2(n_83),
.B1(n_81),
.B2(n_84),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_129),
.A2(n_133),
.B1(n_140),
.B2(n_141),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_130),
.B(n_134),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_152),
.C(n_153),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_126),
.B(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_139),
.B(n_142),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_120),
.A2(n_96),
.B1(n_86),
.B2(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_144),
.B(n_100),
.Y(n_163)
);

NAND2xp33_ASAP7_75t_SL g144 ( 
.A(n_102),
.B(n_33),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_74),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_145),
.B(n_100),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_120),
.A2(n_80),
.B1(n_64),
.B2(n_69),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_156),
.B1(n_117),
.B2(n_116),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_149),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_101),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_74),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_154),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_34),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_103),
.B(n_79),
.C(n_55),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_112),
.A2(n_69),
.B1(n_64),
.B2(n_70),
.Y(n_156)
);

OA21x2_ASAP7_75t_L g182 ( 
.A1(n_157),
.A2(n_55),
.B(n_24),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_151),
.A2(n_116),
.B1(n_106),
.B2(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_160),
.A2(n_188),
.B1(n_106),
.B2(n_124),
.Y(n_202)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_166),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_183),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_111),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_172),
.C(n_175),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_111),
.Y(n_168)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_171),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_134),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_132),
.B(n_26),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_138),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_174),
.B(n_177),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_26),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_141),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI22xp33_ASAP7_75t_R g216 ( 
.A1(n_182),
.A2(n_21),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_130),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_210),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_147),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_197),
.C(n_201),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_186),
.A2(n_139),
.B(n_142),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_175),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_137),
.B(n_136),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_208),
.B1(n_209),
.B2(n_216),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_179),
.A2(n_129),
.B1(n_155),
.B2(n_157),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_196),
.A2(n_169),
.B1(n_183),
.B2(n_174),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_26),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_26),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_202),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_164),
.A2(n_33),
.B(n_0),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_70),
.B1(n_49),
.B2(n_31),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_165),
.Y(n_210)
);

AOI322xp5_ASAP7_75t_L g211 ( 
.A1(n_178),
.A2(n_21),
.A3(n_17),
.B1(n_33),
.B2(n_49),
.C1(n_5),
.C2(n_6),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_180),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_1),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_187),
.Y(n_219)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_214),
.B(n_204),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_221),
.Y(n_253)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_166),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_232),
.B1(n_224),
.B2(n_225),
.Y(n_252)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_225),
.B(n_238),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_198),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_227),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_172),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_228),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_164),
.B1(n_162),
.B2(n_171),
.Y(n_230)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_184),
.B1(n_196),
.B2(n_200),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_233),
.B(n_235),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_236),
.Y(n_255)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g241 ( 
.A(n_237),
.Y(n_241)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_170),
.B(n_190),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_221),
.A2(n_191),
.B(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_195),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_205),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_197),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_257),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_218),
.A2(n_208),
.B1(n_212),
.B2(n_176),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_256),
.A2(n_219),
.B1(n_238),
.B2(n_220),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_229),
.C(n_232),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_262),
.C(n_264),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_255),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_205),
.C(n_233),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_222),
.C(n_223),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_237),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_201),
.C(n_168),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_271),
.C(n_240),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_235),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_182),
.Y(n_271)
);

NOR4xp25_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_9),
.C(n_3),
.D(n_4),
.Y(n_272)
);

NOR2x1_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_13),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_244),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_273),
.A2(n_253),
.B1(n_5),
.B2(n_6),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_251),
.B1(n_254),
.B2(n_242),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_275),
.A2(n_280),
.B1(n_285),
.B2(n_10),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_266),
.A2(n_254),
.B(n_253),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_277),
.A2(n_16),
.B(n_13),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_10),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_251),
.B1(n_258),
.B2(n_245),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_10),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_241),
.C(n_6),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_7),
.C(n_8),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_265),
.A2(n_270),
.B1(n_263),
.B2(n_262),
.Y(n_285)
);

INVx11_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_286),
.A2(n_1),
.B1(n_7),
.B2(n_8),
.Y(n_289)
);

XNOR2x1_ASAP7_75t_L g287 ( 
.A(n_261),
.B(n_11),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_7),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_288),
.Y(n_301)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_283),
.Y(n_303)
);

INVx6_ASAP7_75t_L g291 ( 
.A(n_287),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_292),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_280),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_297),
.B(n_298),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_SL g298 ( 
.A(n_277),
.B(n_14),
.C(n_15),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_294),
.A2(n_274),
.B(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_297),
.C(n_276),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_289),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_281),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_305),
.B(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_308),
.C(n_309),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_275),
.B(n_286),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_284),
.B(n_276),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_291),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_312),
.Y(n_314)
);

O2A1O1Ixp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_301),
.C(n_278),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_313),
.B(n_304),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_299),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule