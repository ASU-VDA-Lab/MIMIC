module fake_jpeg_16902_n_68 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_68);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_68;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_44;
wire n_38;
wire n_26;
wire n_28;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_5),
.B(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_9),
.A2(n_0),
.B(n_1),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_20),
.A2(n_26),
.B(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_24),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_3),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_22),
.A2(n_11),
.B(n_15),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_17),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_16),
.B1(n_6),
.B2(n_4),
.Y(n_29)
);

OR2x4_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_17),
.Y(n_27)
);

AOI21x1_ASAP7_75t_SL g41 ( 
.A1(n_29),
.A2(n_12),
.B(n_39),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_35),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_22),
.B(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g48 ( 
.A(n_34),
.B(n_32),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_22),
.A2(n_15),
.B(n_13),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_20),
.B(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_13),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_8),
.B1(n_12),
.B2(n_19),
.Y(n_39)
);

OAI22x1_ASAP7_75t_SL g44 ( 
.A1(n_39),
.A2(n_35),
.B1(n_29),
.B2(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_32),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_44),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_28),
.Y(n_51)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_30),
.Y(n_55)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_48),
.C(n_42),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_28),
.B(n_53),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_45),
.C(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_40),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_61),
.B(n_49),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_44),
.B(n_41),
.C(n_59),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_65),
.A2(n_59),
.B1(n_46),
.B2(n_54),
.Y(n_67)
);

AOI322xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_66),
.A3(n_54),
.B1(n_58),
.B2(n_40),
.C1(n_49),
.C2(n_52),
.Y(n_68)
);


endmodule