module fake_netlist_6_1423_n_346 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_92, n_42, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_346);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_92;
input n_42;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_346;

wire n_326;
wire n_256;
wire n_209;
wire n_223;
wire n_278;
wire n_341;
wire n_226;
wire n_148;
wire n_161;
wire n_208;
wire n_316;
wire n_304;
wire n_212;
wire n_144;
wire n_168;
wire n_125;
wire n_297;
wire n_342;
wire n_106;
wire n_160;
wire n_131;
wire n_188;
wire n_310;
wire n_186;
wire n_245;
wire n_142;
wire n_143;
wire n_180;
wire n_233;
wire n_255;
wire n_284;
wire n_140;
wire n_337;
wire n_214;
wire n_246;
wire n_289;
wire n_181;
wire n_182;
wire n_238;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_280;
wire n_287;
wire n_230;
wire n_141;
wire n_200;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_229;
wire n_305;
wire n_173;
wire n_250;
wire n_111;
wire n_314;
wire n_183;
wire n_338;
wire n_119;
wire n_235;
wire n_147;
wire n_191;
wire n_340;
wire n_344;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_153;
wire n_156;
wire n_145;
wire n_133;
wire n_96;
wire n_189;
wire n_213;
wire n_294;
wire n_302;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_155;
wire n_109;
wire n_122;
wire n_218;
wire n_234;
wire n_236;
wire n_112;
wire n_172;
wire n_270;
wire n_239;
wire n_126;
wire n_97;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_107;
wire n_103;
wire n_272;
wire n_185;
wire n_293;
wire n_334;
wire n_232;
wire n_163;
wire n_330;
wire n_298;
wire n_281;
wire n_258;
wire n_154;
wire n_98;
wire n_260;
wire n_265;
wire n_313;
wire n_279;
wire n_252;
wire n_228;
wire n_166;
wire n_184;
wire n_216;
wire n_323;
wire n_152;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_102;
wire n_204;
wire n_261;
wire n_312;
wire n_130;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_291;
wire n_219;
wire n_150;
wire n_264;
wire n_263;
wire n_325;
wire n_329;
wire n_237;
wire n_244;
wire n_243;
wire n_124;
wire n_94;
wire n_282;
wire n_116;
wire n_211;
wire n_117;
wire n_175;
wire n_322;
wire n_345;
wire n_231;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_273;
wire n_95;
wire n_311;
wire n_253;
wire n_123;
wire n_136;
wire n_249;
wire n_201;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_241;
wire n_128;
wire n_275;
wire n_276;
wire n_221;
wire n_146;
wire n_318;
wire n_303;
wire n_306;
wire n_193;
wire n_269;
wire n_277;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_268;
wire n_271;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_206;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_317;
wire n_149;
wire n_328;
wire n_195;
wire n_285;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_324;
wire n_335;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_110;
wire n_151;
wire n_267;
wire n_339;
wire n_315;
wire n_288;
wire n_135;
wire n_165;
wire n_259;
wire n_177;
wire n_295;
wire n_190;
wire n_262;
wire n_187;
wire n_170;
wire n_332;
wire n_336;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_3),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_26),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_12),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_19),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_2),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_4),
.Y(n_110)
);

NOR2xp67_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_83),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_21),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_76),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_15),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_0),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_80),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_39),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_2),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_54),
.Y(n_126)
);

CKINVDCx5p33_ASAP7_75t_R g127 ( 
.A(n_22),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_30),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_9),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_24),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_34),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_1),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_48),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_43),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_32),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_20),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_69),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_38),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_63),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_5),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_25),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_31),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_44),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_40),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_35),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_0),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_3),
.Y(n_159)
);

OAI21x1_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_50),
.B(n_91),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_4),
.Y(n_161)
);

OA21x2_ASAP7_75t_L g162 ( 
.A1(n_94),
.A2(n_5),
.B(n_6),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_6),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_7),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_97),
.B(n_7),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_123),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_145),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_95),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_104),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_8),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_105),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_96),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_10),
.Y(n_178)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_99),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_117),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_180)
);

AND2x6_ASAP7_75t_L g181 ( 
.A(n_116),
.B(n_16),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_101),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_165),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_171),
.Y(n_188)
);

OAI22x1_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_102),
.B1(n_103),
.B2(n_152),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_174),
.B(n_106),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_175),
.Y(n_193)
);

AO22x2_ASAP7_75t_L g194 ( 
.A1(n_180),
.A2(n_107),
.B1(n_108),
.B2(n_113),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_177),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_155),
.A2(n_159),
.B1(n_161),
.B2(n_167),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_158),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_163),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_112),
.Y(n_202)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_181),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

OR2x6_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_167),
.Y(n_205)
);

NAND2xp33_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_153),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_118),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_120),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g213 ( 
.A(n_166),
.B(n_154),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_159),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_198),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_187),
.Y(n_220)
);

OR2x6_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_180),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_141),
.B1(n_119),
.B2(n_143),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g223 ( 
.A1(n_206),
.A2(n_183),
.B(n_179),
.C(n_162),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_186),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_195),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

O2A1O1Ixp33_ASAP7_75t_L g228 ( 
.A1(n_210),
.A2(n_179),
.B(n_162),
.C(n_138),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_127),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_131),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_134),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_139),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_137),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

NAND2x1p5_ASAP7_75t_L g237 ( 
.A(n_192),
.B(n_160),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_201),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_191),
.A2(n_151),
.B1(n_150),
.B2(n_149),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_122),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

OR2x6_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_189),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_213),
.B1(n_111),
.B2(n_146),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_211),
.Y(n_247)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_111),
.B(n_147),
.C(n_144),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_241),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_L g254 ( 
.A1(n_223),
.A2(n_148),
.B(n_126),
.C(n_128),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_234),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_125),
.B1(n_130),
.B2(n_132),
.Y(n_260)
);

INVx2_ASAP7_75t_SL g261 ( 
.A(n_236),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_229),
.B(n_230),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_227),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

OR2x6_ASAP7_75t_L g265 ( 
.A(n_221),
.B(n_184),
.Y(n_265)
);

AO21x2_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_228),
.B(n_235),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_243),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_258),
.B(n_257),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_264),
.A2(n_224),
.B(n_231),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_263),
.Y(n_271)
);

AO32x2_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_260),
.A3(n_261),
.B1(n_248),
.B2(n_221),
.Y(n_272)
);

OAI221xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_222),
.B1(n_185),
.B2(n_196),
.C(n_227),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_247),
.A2(n_203),
.B(n_227),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_17),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g276 ( 
.A1(n_262),
.A2(n_23),
.B(n_27),
.Y(n_276)
);

AOI21xp33_ASAP7_75t_SL g277 ( 
.A1(n_255),
.A2(n_36),
.B(n_37),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_242),
.Y(n_279)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_93),
.B(n_46),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_45),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_278),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_253),
.Y(n_284)
);

BUFx8_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

OR2x6_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_256),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_281),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_272),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_287),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_289),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_266),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_282),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_266),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_277),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_270),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_283),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_270),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_290),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_293),
.Y(n_304)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_280),
.B(n_291),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_296),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_291),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_276),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_294),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_276),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_280),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_300),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_275),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_312),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

AND2x4_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_274),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_313),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_314),
.B(n_305),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_322),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_306),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_319),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_329),
.Y(n_332)
);

OAI331xp33_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_328),
.A3(n_320),
.B1(n_319),
.B2(n_316),
.B3(n_325),
.C1(n_324),
.Y(n_333)
);

HB1xp67_ASAP7_75t_SL g334 ( 
.A(n_332),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_333),
.Y(n_335)
);

NOR3xp33_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_306),
.C(n_57),
.Y(n_336)
);

NAND4xp75_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_323),
.C(n_58),
.D(n_59),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_336),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_R g339 ( 
.A(n_337),
.B(n_55),
.Y(n_339)
);

OR4x2_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_67),
.C(n_70),
.D(n_72),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_338),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_342),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_73),
.B1(n_77),
.B2(n_78),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_344),
.Y(n_345)
);

AOI222xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_84),
.B1(n_86),
.B2(n_87),
.C1(n_88),
.C2(n_89),
.Y(n_346)
);


endmodule