module fake_jpeg_11252_n_121 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_121);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_121;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_28),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_16),
.B(n_0),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_53),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_0),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_1),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_51),
.B1(n_47),
.B2(n_41),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_2),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_52),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_63),
.A2(n_43),
.B1(n_5),
.B2(n_6),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_64),
.B(n_75),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_48),
.B1(n_51),
.B2(n_38),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_8),
.B(n_11),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_50),
.C(n_49),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_81),
.C(n_86),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_56),
.B1(n_53),
.B2(n_43),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_56),
.C(n_43),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_87),
.B1(n_88),
.B2(n_19),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_65),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_90),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_87)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_11),
.B(n_12),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_27),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_72),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_24),
.A3(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_20),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_99),
.C(n_101),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_68),
.B1(n_67),
.B2(n_12),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_94),
.A2(n_103),
.B1(n_104),
.B2(n_100),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_95),
.B(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_22),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_23),
.B(n_26),
.Y(n_100)
);

A2O1A1O1Ixp25_ASAP7_75t_L g108 ( 
.A1(n_100),
.A2(n_102),
.B(n_105),
.C(n_97),
.D(n_101),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_77),
.A2(n_30),
.B(n_33),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_86),
.A2(n_81),
.B1(n_76),
.B2(n_87),
.Y(n_104)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.Y(n_113)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_111),
.B(n_102),
.C(n_105),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_114),
.B(n_107),
.C(n_109),
.Y(n_116)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_112),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_116),
.B1(n_108),
.B2(n_97),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_117),
.Y(n_118)
);

OAI21x1_ASAP7_75t_SL g119 ( 
.A1(n_118),
.A2(n_113),
.B(n_112),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_106),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_103),
.Y(n_121)
);


endmodule