module fake_jpeg_45_n_36 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_SL g8 ( 
.A(n_6),
.B(n_2),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_3),
.B(n_4),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_5),
.B(n_0),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_2),
.Y(n_13)
);

AOI22xp33_ASAP7_75t_SL g14 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_18),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_13),
.B(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_19),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_8),
.C(n_10),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_7),
.A2(n_4),
.B1(n_6),
.B2(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_19),
.B1(n_17),
.B2(n_16),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_19),
.B1(n_15),
.B2(n_16),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_21),
.A2(n_18),
.B1(n_17),
.B2(n_14),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_27),
.C(n_17),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_30),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_22),
.B(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_26),
.Y(n_33)
);

OAI21x1_ASAP7_75t_SL g34 ( 
.A1(n_33),
.A2(n_32),
.B(n_30),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g36 ( 
.A(n_35),
.Y(n_36)
);


endmodule