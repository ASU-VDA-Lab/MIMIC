module fake_jpeg_32117_n_34 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_0),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_0),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_21),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_15),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_20),
.A2(n_16),
.B(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_4),
.Y(n_26)
);

OAI32xp33_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_24),
.A3(n_16),
.B1(n_17),
.B2(n_8),
.Y(n_27)
);

AND2x6_ASAP7_75t_L g24 ( 
.A(n_21),
.B(n_14),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_4),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_7),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_9),
.B(n_10),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_11),
.B(n_13),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_30),
.B(n_28),
.Y(n_33)
);

BUFx24_ASAP7_75t_SL g34 ( 
.A(n_33),
.Y(n_34)
);


endmodule