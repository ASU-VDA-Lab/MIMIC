module fake_jpeg_28972_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_15),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_54),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_19),
.B(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_55),
.B(n_59),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_58),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_19),
.B(n_5),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_5),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_62),
.B(n_65),
.Y(n_157)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_33),
.A2(n_5),
.B1(n_13),
.B2(n_2),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_64),
.A2(n_48),
.B1(n_45),
.B2(n_39),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_4),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_25),
.B(n_4),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_49),
.C(n_48),
.Y(n_152)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_31),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_72),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_74),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_75),
.Y(n_160)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_93),
.Y(n_115)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_85),
.Y(n_162)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_24),
.Y(n_87)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g132 ( 
.A(n_88),
.Y(n_132)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_90),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_35),
.Y(n_96)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_96),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_22),
.B(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_103),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g98 ( 
.A(n_36),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_104),
.Y(n_120)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_36),
.Y(n_99)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_4),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_40),
.Y(n_105)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_105),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_16),
.B1(n_44),
.B2(n_43),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_148),
.B1(n_149),
.B2(n_134),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_62),
.B(n_30),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_137),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g128 ( 
.A(n_68),
.B(n_41),
.CON(n_128),
.SN(n_128)
);

NAND2xp67_ASAP7_75t_SL g201 ( 
.A(n_128),
.B(n_28),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_40),
.B1(n_44),
.B2(n_43),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_134),
.A2(n_98),
.B1(n_101),
.B2(n_75),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_65),
.B(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_64),
.B(n_26),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_139),
.B(n_165),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_50),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_147),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_87),
.B(n_49),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_99),
.A2(n_44),
.B1(n_43),
.B2(n_21),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_52),
.A2(n_21),
.B1(n_47),
.B2(n_38),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_26),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_167),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_23),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g184 ( 
.A1(n_164),
.A2(n_42),
.B1(n_23),
.B2(n_20),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_53),
.B(n_37),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_69),
.B(n_39),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_116),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_38),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_170),
.B(n_171),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_42),
.Y(n_171)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_183),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_174),
.B(n_181),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_153),
.B1(n_141),
.B2(n_131),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_175),
.A2(n_178),
.B1(n_161),
.B2(n_146),
.Y(n_246)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_105),
.B1(n_96),
.B2(n_91),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g181 ( 
.A(n_128),
.B(n_0),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_110),
.Y(n_182)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_182),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_120),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_127),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_187),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_56),
.B1(n_82),
.B2(n_77),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_186),
.A2(n_190),
.B1(n_161),
.B2(n_160),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_151),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g188 ( 
.A1(n_163),
.A2(n_73),
.B1(n_58),
.B2(n_21),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g252 ( 
.A1(n_188),
.A2(n_112),
.B1(n_125),
.B2(n_118),
.Y(n_252)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_113),
.A2(n_93),
.A3(n_45),
.B1(n_37),
.B2(n_30),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_189),
.B(n_191),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_192),
.Y(n_241)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_20),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_210),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_121),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_197),
.Y(n_226)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_136),
.B(n_47),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_203),
.Y(n_237)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_200),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_202),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_119),
.B(n_28),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_132),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_204),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_151),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_205),
.B(n_206),
.Y(n_238)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_93),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_207),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_208),
.Y(n_250)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_209),
.A2(n_212),
.B1(n_214),
.B2(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_123),
.B(n_28),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_10),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_211),
.B(n_215),
.Y(n_245)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_129),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_108),
.B(n_28),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_125),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_109),
.A2(n_28),
.B1(n_10),
.B2(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_149),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_215),
.A2(n_106),
.B1(n_158),
.B2(n_160),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_224),
.A2(n_246),
.B1(n_252),
.B2(n_112),
.Y(n_276)
);

OAI32xp33_ASAP7_75t_L g229 ( 
.A1(n_180),
.A2(n_114),
.A3(n_148),
.B1(n_107),
.B2(n_135),
.Y(n_229)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_132),
.B1(n_122),
.B2(n_158),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_232),
.B(n_155),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_234),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_170),
.B(n_140),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_140),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_251),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_178),
.B1(n_175),
.B2(n_190),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_173),
.A2(n_109),
.B1(n_118),
.B2(n_155),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_242),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_194),
.B(n_146),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_231),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_259),
.Y(n_286)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_241),
.Y(n_256)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_258),
.A2(n_264),
.B1(n_269),
.B2(n_271),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_191),
.C(n_181),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_279),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_222),
.A2(n_202),
.B(n_210),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_261),
.A2(n_237),
.B(n_246),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_263),
.B(n_267),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_244),
.A2(n_213),
.B1(n_184),
.B2(n_188),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_266),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g269 ( 
.A1(n_232),
.A2(n_169),
.B1(n_188),
.B2(n_184),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_243),
.A2(n_216),
.B1(n_212),
.B2(n_204),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_270),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_244),
.A2(n_184),
.B1(n_189),
.B2(n_196),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_274),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_247),
.A2(n_230),
.B1(n_245),
.B2(n_236),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_273),
.A2(n_282),
.B1(n_243),
.B2(n_253),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_237),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_245),
.B1(n_252),
.B2(n_229),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_220),
.B(n_195),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_277),
.B(n_278),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_220),
.B(n_181),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_222),
.A2(n_202),
.B1(n_191),
.B2(n_182),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_236),
.B1(n_251),
.B2(n_263),
.Y(n_293)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_222),
.A2(n_192),
.B1(n_200),
.B2(n_193),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_197),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_226),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_284),
.Y(n_287)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_218),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_253),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_294),
.A2(n_301),
.B1(n_293),
.B2(n_303),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_300),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_255),
.B(n_267),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_297),
.B(n_298),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_239),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_299),
.B(n_260),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_283),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_262),
.A2(n_236),
.B1(n_233),
.B2(n_252),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_303),
.A2(n_313),
.B(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_310),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_225),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_306),
.B(n_299),
.C(n_308),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_284),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_309),
.A2(n_276),
.B1(n_275),
.B2(n_257),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_266),
.B(n_225),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_312),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_262),
.A2(n_221),
.B(n_252),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_254),
.A2(n_219),
.B1(n_250),
.B2(n_249),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_314),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_302),
.B(n_277),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_318),
.B(n_334),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_338),
.B1(n_345),
.B2(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_321),
.Y(n_350)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_322),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_324),
.B(n_332),
.Y(n_353)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_327),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_290),
.A2(n_264),
.B(n_282),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_335),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_329),
.A2(n_313),
.B1(n_296),
.B2(n_304),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_330),
.B(n_347),
.C(n_298),
.Y(n_360)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_290),
.B(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_331),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g332 ( 
.A1(n_288),
.A2(n_258),
.B1(n_268),
.B2(n_280),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_297),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_312),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_306),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_285),
.Y(n_337)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_288),
.A2(n_257),
.B1(n_275),
.B2(n_270),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_287),
.A2(n_261),
.B(n_278),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_340),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_307),
.A2(n_250),
.B(n_249),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_289),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_344),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g343 ( 
.A(n_300),
.B(n_302),
.Y(n_343)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g344 ( 
.A(n_286),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_219),
.B1(n_281),
.B2(n_256),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_223),
.C(n_226),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_305),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_348),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_355),
.B(n_360),
.C(n_365),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_323),
.Y(n_356)
);

BUFx12f_ASAP7_75t_L g395 ( 
.A(n_356),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_322),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_357),
.B(n_358),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_343),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_361),
.A2(n_362),
.B1(n_366),
.B2(n_372),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_316),
.B1(n_308),
.B2(n_314),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_334),
.B1(n_345),
.B2(n_319),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_304),
.C(n_296),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_338),
.A2(n_313),
.B1(n_289),
.B2(n_311),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_336),
.B(n_223),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_367),
.B(n_376),
.Y(n_389)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_337),
.Y(n_370)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_291),
.C(n_228),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_371),
.B(n_340),
.C(n_326),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_328),
.A2(n_291),
.B1(n_256),
.B2(n_281),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_343),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_374),
.B(n_375),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_319),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_339),
.B(n_179),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_329),
.B(n_317),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_378),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_317),
.B(n_132),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_351),
.B(n_331),
.Y(n_381)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_381),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_331),
.B(n_333),
.Y(n_383)
);

AO21x1_ASAP7_75t_L g418 ( 
.A1(n_383),
.A2(n_394),
.B(n_403),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_323),
.Y(n_384)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_384),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_356),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_386),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_373),
.Y(n_387)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_376),
.B(n_335),
.Y(n_388)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_388),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_390),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_379),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_396),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_354),
.A2(n_346),
.B(n_326),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_380),
.Y(n_396)
);

OA22x2_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_327),
.B1(n_321),
.B2(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_399),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_344),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_400),
.A2(n_401),
.B1(n_369),
.B2(n_368),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_355),
.B(n_342),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_360),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_368),
.A2(n_364),
.B(n_353),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_405),
.C(n_408),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_367),
.B(n_342),
.C(n_320),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_352),
.Y(n_406)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_406),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_365),
.B(n_332),
.C(n_325),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_409),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_411),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_371),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_426),
.C(n_430),
.Y(n_435)
);

A2O1A1Ixp33_ASAP7_75t_L g413 ( 
.A1(n_403),
.A2(n_353),
.B(n_350),
.C(n_363),
.Y(n_413)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_394),
.A2(n_383),
.B(n_398),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_416),
.A2(n_219),
.B(n_265),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_366),
.C(n_378),
.Y(n_426)
);

BUFx4f_ASAP7_75t_SL g427 ( 
.A(n_395),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_427),
.Y(n_448)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_395),
.Y(n_428)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_428),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_361),
.B1(n_372),
.B2(n_332),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_429),
.B(n_241),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_332),
.C(n_324),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_341),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_431),
.B(n_407),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_408),
.B(n_341),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_432),
.B(n_407),
.C(n_405),
.Y(n_438)
);

FAx1_ASAP7_75t_SL g436 ( 
.A(n_433),
.B(n_384),
.CI(n_402),
.CON(n_436),
.SN(n_436)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_436),
.B(n_441),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_439),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_389),
.C(n_391),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_433),
.B(n_399),
.CI(n_386),
.CON(n_442),
.SN(n_442)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_443),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_422),
.B(n_399),
.C(n_382),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_415),
.A2(n_382),
.B1(n_393),
.B2(n_406),
.Y(n_444)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_444),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_425),
.A2(n_409),
.B1(n_385),
.B2(n_399),
.Y(n_445)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_445),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_423),
.B(n_395),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_446),
.B(n_452),
.Y(n_469)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_447),
.Y(n_465)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_420),
.Y(n_449)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_450),
.A2(n_451),
.B1(n_420),
.B2(n_421),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_419),
.A2(n_228),
.B1(n_172),
.B2(n_248),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_414),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_235),
.C(n_248),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_431),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_419),
.A2(n_235),
.B1(n_227),
.B2(n_187),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_454),
.A2(n_421),
.B1(n_428),
.B2(n_413),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_432),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_464),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_434),
.A2(n_418),
.B(n_416),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_460),
.B(n_473),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_468),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_462),
.A2(n_463),
.B1(n_467),
.B2(n_457),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_434),
.A2(n_417),
.B1(n_424),
.B2(n_430),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_450),
.A2(n_418),
.B1(n_414),
.B2(n_426),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_437),
.Y(n_468)
);

INVx13_ASAP7_75t_L g470 ( 
.A(n_448),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_470),
.B(n_448),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_454),
.A2(n_411),
.B1(n_427),
.B2(n_227),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_471),
.A2(n_451),
.B1(n_447),
.B2(n_449),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_443),
.A2(n_427),
.B(n_227),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_442),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_475),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_477),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_460),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_SL g479 ( 
.A(n_468),
.B(n_435),
.C(n_441),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_479),
.A2(n_483),
.B(n_489),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_480),
.B(n_3),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_458),
.B(n_438),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_481),
.B(n_482),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_442),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_471),
.B(n_436),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_458),
.B(n_453),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_SL g501 ( 
.A(n_485),
.B(n_486),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_440),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_487),
.B(n_473),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_440),
.B1(n_436),
.B2(n_168),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_488),
.A2(n_206),
.B1(n_198),
.B2(n_130),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_176),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_483),
.B(n_455),
.CI(n_462),
.CON(n_490),
.SN(n_490)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_490),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_SL g492 ( 
.A1(n_477),
.A2(n_465),
.B(n_470),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g507 ( 
.A1(n_492),
.A2(n_497),
.B(n_3),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_493),
.B(n_494),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_474),
.A2(n_459),
.B1(n_209),
.B2(n_166),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_495),
.B(n_502),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_476),
.A2(n_130),
.B(n_117),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_0),
.C(n_1),
.Y(n_499)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_499),
.B(n_484),
.Y(n_505)
);

NOR2xp67_ASAP7_75t_SL g504 ( 
.A(n_491),
.B(n_484),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g512 ( 
.A1(n_504),
.A2(n_500),
.B(n_498),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_511),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_496),
.B(n_3),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_506),
.A2(n_509),
.B(n_11),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_SL g516 ( 
.A1(n_507),
.A2(n_497),
.B(n_492),
.C(n_502),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_490),
.B(n_10),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_501),
.B(n_11),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_515),
.B(n_514),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_516),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_493),
.B(n_499),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_517),
.A2(n_519),
.B(n_503),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_512),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_518),
.A2(n_507),
.B(n_510),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_520),
.B(n_521),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_12),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_12),
.C(n_14),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_524),
.A2(n_12),
.B1(n_0),
.B2(n_1),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_525),
.B(n_1),
.Y(n_526)
);


endmodule