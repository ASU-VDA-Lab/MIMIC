module fake_jpeg_21675_n_182 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_182);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_13),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR3xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_0),
.C(n_1),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_22),
.B1(n_11),
.B2(n_20),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_12),
.B(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_31),
.Y(n_39)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_28),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_17),
.B1(n_20),
.B2(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_36),
.A2(n_41),
.B1(n_26),
.B2(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_31),
.A2(n_17),
.B1(n_20),
.B2(n_16),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_51),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_52),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_39),
.A2(n_38),
.B(n_23),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_48),
.B(n_38),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_25),
.C(n_27),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_27),
.C(n_25),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_50),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_23),
.B(n_30),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_53),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_39),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_56),
.Y(n_67)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_26),
.B1(n_17),
.B2(n_14),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_51),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_60),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_50),
.B(n_25),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_64),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_44),
.B(n_25),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_27),
.C(n_40),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_29),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_41),
.Y(n_71)
);

AO21x2_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_67),
.B(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_77),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_65),
.A2(n_53),
.B(n_54),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_83),
.B(n_59),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_44),
.B1(n_48),
.B2(n_45),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_68),
.B1(n_70),
.B2(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_72),
.A2(n_43),
.B1(n_56),
.B2(n_45),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_78),
.A2(n_68),
.B1(n_37),
.B2(n_40),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_88),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_71),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_86),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_69),
.B(n_55),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_42),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_R g89 ( 
.A1(n_80),
.A2(n_71),
.B(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_95),
.B1(n_86),
.B2(n_84),
.Y(n_110)
);

XNOR2x1_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_57),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_96),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_82),
.A2(n_42),
.B1(n_61),
.B2(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_102),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_34),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_104),
.C(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_34),
.C(n_19),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_19),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_83),
.Y(n_124)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_116),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_121),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_83),
.C(n_80),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_99),
.C(n_105),
.Y(n_127)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_78),
.B1(n_75),
.B2(n_104),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_21),
.B1(n_18),
.B2(n_22),
.Y(n_133)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_115),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_118),
.B(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_106),
.B(n_73),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_81),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_125),
.B(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_135),
.C(n_109),
.Y(n_140)
);

OAI321xp33_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_80),
.A3(n_96),
.B1(n_87),
.B2(n_81),
.C(n_14),
.Y(n_129)
);

AOI31xp67_ASAP7_75t_L g143 ( 
.A1(n_129),
.A2(n_131),
.A3(n_133),
.B(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_133),
.Y(n_147)
);

OAI321xp33_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_15),
.A3(n_14),
.B1(n_18),
.B2(n_21),
.C(n_6),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_19),
.C(n_15),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_22),
.B1(n_15),
.B2(n_14),
.Y(n_138)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_15),
.B1(n_19),
.B2(n_2),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_145),
.C(n_114),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_146),
.B(n_136),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_119),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_135),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_109),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_116),
.B(n_115),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_124),
.Y(n_148)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_136),
.B1(n_134),
.B2(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_150),
.A2(n_154),
.B1(n_147),
.B2(n_2),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_151),
.B(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_136),
.B1(n_112),
.B2(n_137),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_139),
.C(n_3),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_3),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_163),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_10),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_165),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_155),
.C(n_157),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_5),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_161),
.B(n_153),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_168),
.A2(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_159),
.B(n_160),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_5),
.B(n_7),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_169),
.A2(n_5),
.B(n_8),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_166),
.B(n_9),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_177),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_178),
.A2(n_9),
.B(n_10),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_9),
.C(n_2),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_179),
.Y(n_182)
);


endmodule