module real_aes_17615_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AND2x4_ASAP7_75t_L g860 ( .A(n_0), .B(n_861), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_1), .A2(n_32), .B1(n_139), .B2(n_231), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g583 ( .A1(n_2), .A2(n_9), .B1(n_536), .B2(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g861 ( .A(n_3), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g550 ( .A(n_4), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_5), .A2(n_11), .B1(n_537), .B2(n_573), .Y(n_572) );
OR2x2_ASAP7_75t_L g112 ( .A(n_6), .B(n_28), .Y(n_112) );
BUFx2_ASAP7_75t_L g856 ( .A(n_6), .Y(n_856) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_7), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_8), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g863 ( .A(n_10), .Y(n_863) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_12), .B(n_154), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_13), .A2(n_97), .B1(n_184), .B2(n_536), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_14), .A2(n_29), .B1(n_554), .B2(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_15), .B(n_154), .Y(n_551) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_16), .A2(n_46), .B(n_135), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_17), .B(n_235), .Y(n_234) );
CKINVDCx5p33_ASAP7_75t_R g609 ( .A(n_18), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_19), .A2(n_36), .B1(n_191), .B2(n_206), .Y(n_562) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_20), .Y(n_259) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_21), .A2(n_43), .B1(n_206), .B2(n_536), .Y(n_592) );
CKINVDCx5p33_ASAP7_75t_R g528 ( .A(n_22), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_23), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_24), .B(n_214), .Y(n_233) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_25), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_26), .B(n_132), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_27), .Y(n_183) );
HB1xp67_ASAP7_75t_L g855 ( .A(n_28), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_30), .A2(n_81), .B1(n_139), .B2(n_522), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_31), .A2(n_35), .B1(n_139), .B2(n_539), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_33), .A2(n_49), .B1(n_536), .B2(n_591), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g263 ( .A(n_34), .Y(n_263) );
XOR2xp5_ASAP7_75t_L g113 ( .A(n_37), .B(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_38), .Y(n_832) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_39), .B(n_154), .Y(n_202) );
INVx2_ASAP7_75t_L g107 ( .A(n_40), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_41), .B(n_187), .Y(n_229) );
BUFx3_ASAP7_75t_L g110 ( .A(n_42), .Y(n_110) );
INVx1_ASAP7_75t_L g827 ( .A(n_42), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_44), .B(n_173), .Y(n_237) );
XOR2x2_ASAP7_75t_L g121 ( .A(n_45), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g265 ( .A(n_47), .B(n_173), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_48), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_50), .B(n_214), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_51), .B(n_191), .Y(n_190) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_52), .A2(n_68), .B1(n_191), .B2(n_591), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_53), .A2(n_71), .B1(n_139), .B2(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_54), .B(n_295), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_55), .A2(n_143), .B(n_152), .C(n_258), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g535 ( .A1(n_56), .A2(n_94), .B1(n_536), .B2(n_537), .Y(n_535) );
INVx1_ASAP7_75t_L g135 ( .A(n_57), .Y(n_135) );
AND2x4_ASAP7_75t_L g157 ( .A(n_58), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_59), .A2(n_60), .B1(n_206), .B2(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_61), .B(n_132), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_62), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g264 ( .A(n_63), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_64), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g158 ( .A(n_65), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_66), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_67), .B(n_132), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_69), .B(n_139), .Y(n_290) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_70), .B(n_187), .C(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_72), .B(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_73), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g165 ( .A(n_74), .B(n_166), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_75), .B(n_154), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_76), .B(n_148), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_77), .A2(n_93), .B1(n_152), .B2(n_206), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g828 ( .A1(n_78), .A2(n_121), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g830 ( .A(n_78), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_79), .Y(n_594) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_80), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_82), .A2(n_88), .B1(n_213), .B2(n_214), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_83), .B(n_154), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_84), .Y(n_846) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_85), .B(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_86), .B(n_185), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_87), .B(n_132), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g576 ( .A(n_89), .Y(n_576) );
INVx1_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
NOR2xp33_ASAP7_75t_L g825 ( .A(n_90), .B(n_826), .Y(n_825) );
NAND2xp33_ASAP7_75t_L g555 ( .A(n_91), .B(n_154), .Y(n_555) );
NAND2xp33_ASAP7_75t_L g141 ( .A(n_92), .B(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_95), .B(n_173), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g167 ( .A(n_96), .B(n_142), .C(n_166), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_98), .B(n_139), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_99), .B(n_214), .Y(n_293) );
AOI21xp5_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_851), .B(n_862), .Y(n_100) );
OR2x6_ASAP7_75t_L g101 ( .A(n_102), .B(n_845), .Y(n_101) );
OAI21x1_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_113), .B(n_821), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
BUFx12f_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x6_ASAP7_75t_SL g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
AND2x2_ASAP7_75t_L g822 ( .A(n_107), .B(n_823), .Y(n_822) );
NOR2xp33_ASAP7_75t_L g835 ( .A(n_107), .B(n_836), .Y(n_835) );
INVx3_ASAP7_75t_L g843 ( .A(n_107), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NOR2x1_ASAP7_75t_L g838 ( .A(n_110), .B(n_112), .Y(n_838) );
AND2x6_ASAP7_75t_SL g824 ( .A(n_111), .B(n_825), .Y(n_824) );
AND3x2_ASAP7_75t_L g848 ( .A(n_111), .B(n_849), .C(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_121), .B(n_510), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_116), .Y(n_115) );
AND2x2_ASAP7_75t_L g510 ( .A(n_116), .B(n_511), .Y(n_510) );
INVx8_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
BUFx12f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
AND2x2_ASAP7_75t_L g837 ( .A(n_119), .B(n_838), .Y(n_837) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_L g850 ( .A(n_120), .Y(n_850) );
INVx1_ASAP7_75t_L g829 ( .A(n_121), .Y(n_829) );
OR2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_442), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_317), .C(n_357), .D(n_406), .Y(n_123) );
NOR2xp67_ASAP7_75t_L g124 ( .A(n_125), .B(n_266), .Y(n_124) );
OAI22xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_176), .B1(n_238), .B2(n_247), .Y(n_125) );
INVx1_ASAP7_75t_L g438 ( .A(n_126), .Y(n_438) );
INVx1_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_127), .B(n_285), .Y(n_354) );
AND2x2_ASAP7_75t_L g385 ( .A(n_127), .B(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_159), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_128), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g309 ( .A(n_128), .Y(n_309) );
AND2x2_ASAP7_75t_L g484 ( .A(n_128), .B(n_352), .Y(n_484) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
BUFx2_ASAP7_75t_L g249 ( .A(n_129), .Y(n_249) );
AND2x2_ASAP7_75t_L g337 ( .A(n_129), .B(n_299), .Y(n_337) );
AND2x2_ASAP7_75t_L g381 ( .A(n_129), .B(n_286), .Y(n_381) );
OR2x2_ASAP7_75t_L g399 ( .A(n_129), .B(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g303 ( .A(n_130), .B(n_286), .Y(n_303) );
BUFx2_ASAP7_75t_L g360 ( .A(n_130), .Y(n_360) );
OR2x2_ASAP7_75t_L g368 ( .A(n_130), .B(n_326), .Y(n_368) );
INVx1_ASAP7_75t_L g423 ( .A(n_130), .Y(n_423) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
INVx2_ASAP7_75t_L g563 ( .A(n_132), .Y(n_563) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_SL g155 ( .A(n_133), .B(n_156), .Y(n_155) );
INVx1_ASAP7_75t_SL g162 ( .A(n_133), .Y(n_162) );
INVx2_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
BUFx3_ASAP7_75t_L g519 ( .A(n_133), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_133), .B(n_543), .Y(n_542) );
INVx2_ASAP7_75t_SL g547 ( .A(n_133), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_133), .B(n_565), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_133), .B(n_586), .Y(n_585) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
OAI21x1_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_146), .B(n_155), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_143), .Y(n_137) );
OAI22xp33_ASAP7_75t_L g262 ( .A1(n_139), .A2(n_206), .B1(n_263), .B2(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g537 ( .A(n_139), .Y(n_537) );
INVx4_ASAP7_75t_L g539 ( .A(n_139), .Y(n_539) );
INVx1_ASAP7_75t_L g591 ( .A(n_139), .Y(n_591) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_140), .Y(n_142) );
INVx1_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
INVx1_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx1_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_140), .Y(n_206) );
INVx1_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
INVx1_ASAP7_75t_L g218 ( .A(n_140), .Y(n_218) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_140), .Y(n_231) );
INVx2_ASAP7_75t_L g260 ( .A(n_140), .Y(n_260) );
INVx2_ASAP7_75t_L g191 ( .A(n_142), .Y(n_191) );
INVx1_ASAP7_75t_L g554 ( .A(n_142), .Y(n_554) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_143), .A2(n_169), .B(n_171), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_143), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_143), .A2(n_290), .B(n_291), .Y(n_289) );
BUFx4f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx2_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
INVx1_ASAP7_75t_L g166 ( .A(n_145), .Y(n_166) );
BUFx8_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_149), .B1(n_151), .B2(n_153), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_148), .A2(n_189), .B(n_190), .Y(n_188) );
INVx2_ASAP7_75t_SL g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g220 ( .A(n_150), .Y(n_220) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g164 ( .A1(n_154), .A2(n_165), .B(n_167), .Y(n_164) );
INVx1_ASAP7_75t_L g235 ( .A(n_154), .Y(n_235) );
INVx3_ASAP7_75t_L g536 ( .A(n_154), .Y(n_536) );
OAI21x1_ASAP7_75t_L g163 ( .A1(n_156), .A2(n_164), .B(n_168), .Y(n_163) );
OAI21x1_ASAP7_75t_L g181 ( .A1(n_156), .A2(n_182), .B(n_188), .Y(n_181) );
OAI21x1_ASAP7_75t_L g199 ( .A1(n_156), .A2(n_200), .B(n_203), .Y(n_199) );
OAI21x1_ASAP7_75t_L g227 ( .A1(n_156), .A2(n_228), .B(n_232), .Y(n_227) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_156), .A2(n_289), .B(n_292), .Y(n_288) );
BUFx10_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx10_ASAP7_75t_L g222 ( .A(n_157), .Y(n_222) );
INVx1_ASAP7_75t_L g526 ( .A(n_157), .Y(n_526) );
AND2x2_ASAP7_75t_L g250 ( .A(n_159), .B(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g362 ( .A(n_159), .B(n_339), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_159), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx1_ASAP7_75t_L g400 ( .A(n_160), .Y(n_400) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_160), .Y(n_405) );
AND2x2_ASAP7_75t_L g422 ( .A(n_160), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g312 ( .A(n_161), .B(n_252), .Y(n_312) );
INVx1_ASAP7_75t_L g326 ( .A(n_161), .Y(n_326) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_172), .Y(n_161) );
INVx1_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
INVx1_ASAP7_75t_L g524 ( .A(n_166), .Y(n_524) );
INVx1_ASAP7_75t_SL g540 ( .A(n_166), .Y(n_540) );
INVx1_ASAP7_75t_L g582 ( .A(n_170), .Y(n_582) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx2_ASAP7_75t_L g180 ( .A(n_174), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_174), .B(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_174), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g221 ( .A(n_175), .Y(n_221) );
INVx2_ASAP7_75t_L g225 ( .A(n_175), .Y(n_225) );
NAND2x1_ASAP7_75t_L g176 ( .A(n_177), .B(n_193), .Y(n_176) );
AND2x4_ASAP7_75t_L g487 ( .A(n_177), .B(n_415), .Y(n_487) );
INVxp67_ASAP7_75t_SL g177 ( .A(n_178), .Y(n_177) );
INVxp67_ASAP7_75t_SL g246 ( .A(n_178), .Y(n_246) );
BUFx3_ASAP7_75t_L g281 ( .A(n_178), .Y(n_281) );
INVx1_ASAP7_75t_L g347 ( .A(n_178), .Y(n_347) );
AND2x2_ASAP7_75t_L g350 ( .A(n_178), .B(n_196), .Y(n_350) );
AND2x2_ASAP7_75t_L g375 ( .A(n_178), .B(n_226), .Y(n_375) );
INVx1_ASAP7_75t_L g378 ( .A(n_178), .Y(n_378) );
AND2x2_ASAP7_75t_L g410 ( .A(n_178), .B(n_275), .Y(n_410) );
INVx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_192), .Y(n_179) );
OAI21xp5_ASAP7_75t_L g276 ( .A1(n_180), .A2(n_181), .B(n_192), .Y(n_276) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_180), .A2(n_288), .B(n_297), .Y(n_287) );
OAI21xp33_ASAP7_75t_SL g315 ( .A1(n_180), .A2(n_288), .B(n_297), .Y(n_315) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_186), .C(n_187), .Y(n_182) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_187), .A2(n_204), .B(n_205), .Y(n_203) );
INVx6_ASAP7_75t_L g216 ( .A(n_187), .Y(n_216) );
O2A1O1Ixp5_ASAP7_75t_L g549 ( .A1(n_187), .A2(n_539), .B(n_550), .C(n_551), .Y(n_549) );
AND2x4_ASAP7_75t_L g193 ( .A(n_194), .B(n_208), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g319 ( .A(n_195), .B(n_305), .Y(n_319) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_L g345 ( .A(n_197), .B(n_332), .Y(n_345) );
AND2x2_ASAP7_75t_L g374 ( .A(n_197), .B(n_210), .Y(n_374) );
OR2x2_ASAP7_75t_L g470 ( .A(n_197), .B(n_210), .Y(n_470) );
OAI21x1_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_197) );
OA21x2_ASAP7_75t_L g226 ( .A1(n_198), .A2(n_227), .B(n_237), .Y(n_226) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_244) );
OAI21x1_ASAP7_75t_L g275 ( .A1(n_198), .A2(n_227), .B(n_237), .Y(n_275) );
INVx2_ASAP7_75t_L g213 ( .A(n_206), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_206), .A2(n_229), .B(n_230), .Y(n_228) );
AND2x2_ASAP7_75t_L g349 ( .A(n_208), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g498 ( .A(n_208), .Y(n_498) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_209), .Y(n_240) );
OR2x2_ASAP7_75t_L g432 ( .A(n_209), .B(n_242), .Y(n_432) );
INVx1_ASAP7_75t_L g454 ( .A(n_209), .Y(n_454) );
OR2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_226), .Y(n_209) );
AND2x2_ASAP7_75t_L g270 ( .A(n_210), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_275), .Y(n_305) );
INVx1_ASAP7_75t_L g332 ( .A(n_210), .Y(n_332) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_210), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_210), .B(n_226), .Y(n_419) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_221), .A3(n_222), .B(n_223), .Y(n_210) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_216), .B1(n_217), .B2(n_219), .Y(n_211) );
INVx1_ASAP7_75t_L g573 ( .A(n_214), .Y(n_573) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_216), .A2(n_521), .B1(n_523), .B2(n_524), .Y(n_520) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_216), .A2(n_535), .B1(n_538), .B2(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_216), .A2(n_553), .B(n_555), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_216), .A2(n_219), .B1(n_561), .B2(n_562), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_216), .A2(n_540), .B1(n_572), .B2(n_574), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_216), .A2(n_219), .B1(n_581), .B2(n_583), .Y(n_580) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_216), .A2(n_219), .B1(n_590), .B2(n_592), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_216), .A2(n_219), .B1(n_606), .B2(n_607), .Y(n_605) );
INVx1_ASAP7_75t_L g584 ( .A(n_218), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_219), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g296 ( .A(n_220), .Y(n_296) );
INVx2_ASAP7_75t_L g254 ( .A(n_221), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_221), .B(n_528), .Y(n_527) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_221), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g255 ( .A(n_222), .Y(n_255) );
AO31x2_ASAP7_75t_L g559 ( .A1(n_222), .A2(n_560), .A3(n_563), .B(n_564), .Y(n_559) );
AO31x2_ASAP7_75t_L g570 ( .A1(n_222), .A2(n_533), .A3(n_571), .B(n_575), .Y(n_570) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_222), .A2(n_519), .A3(n_580), .B(n_585), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_224), .B(n_225), .Y(n_223) );
BUFx2_ASAP7_75t_L g533 ( .A(n_225), .Y(n_533) );
AND2x2_ASAP7_75t_L g356 ( .A(n_226), .B(n_276), .Y(n_356) );
INVx2_ASAP7_75t_L g295 ( .A(n_231), .Y(n_295) );
AOI21x1_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_236), .Y(n_232) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NOR3x1_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .C(n_245), .Y(n_239) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_242), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g304 ( .A(n_242), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g355 ( .A(n_242), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g395 ( .A(n_242), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_242), .B(n_418), .Y(n_450) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_243), .B(n_331), .Y(n_391) );
AND2x2_ASAP7_75t_L g415 ( .A(n_243), .B(n_275), .Y(n_415) );
BUFx3_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g271 ( .A(n_244), .Y(n_271) );
BUFx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g426 ( .A(n_246), .B(n_305), .Y(n_426) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_250), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_249), .B(n_312), .Y(n_491) );
AND2x4_ASAP7_75t_L g483 ( .A(n_250), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_250), .B(n_303), .Y(n_497) );
INVx2_ASAP7_75t_L g299 ( .A(n_251), .Y(n_299) );
INVx1_ASAP7_75t_L g302 ( .A(n_251), .Y(n_302) );
INVx2_ASAP7_75t_L g387 ( .A(n_251), .Y(n_387) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g371 ( .A(n_252), .Y(n_371) );
AOI21x1_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_256), .B(n_265), .Y(n_252) );
NOR2xp67_ASAP7_75t_SL g253 ( .A(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g588 ( .A(n_254), .Y(n_588) );
INVx1_ASAP7_75t_L g541 ( .A(n_255), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_261), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
INVx2_ASAP7_75t_SL g522 ( .A(n_260), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_306), .Y(n_266) );
AOI22xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_282), .B1(n_300), .B2(n_304), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_277), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g334 ( .A(n_270), .B(n_281), .Y(n_334) );
AND2x2_ASAP7_75t_L g494 ( .A(n_270), .B(n_375), .Y(n_494) );
BUFx2_ASAP7_75t_L g365 ( .A(n_271), .Y(n_365) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g364 ( .A(n_274), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g279 ( .A(n_275), .Y(n_279) );
INVx1_ASAP7_75t_L g331 ( .A(n_275), .Y(n_331) );
INVx1_ASAP7_75t_L g456 ( .A(n_276), .Y(n_456) );
AOI31xp33_ASAP7_75t_L g474 ( .A1(n_277), .A2(n_475), .A3(n_476), .B(n_477), .Y(n_474) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_278), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_279), .B(n_374), .Y(n_473) );
INVx2_ASAP7_75t_L g501 ( .A(n_279), .Y(n_501) );
INVxp67_ASAP7_75t_SL g316 ( .A(n_280), .Y(n_316) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g329 ( .A(n_281), .B(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_281), .B(n_391), .Y(n_390) );
OR2x2_ASAP7_75t_L g459 ( .A(n_281), .B(n_419), .Y(n_459) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_298), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g370 ( .A(n_286), .B(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B(n_296), .Y(n_292) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
HB1xp67_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
INVx1_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
INVx1_ASAP7_75t_L g343 ( .A(n_303), .Y(n_343) );
AND2x2_ASAP7_75t_L g404 ( .A(n_303), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g460 ( .A(n_303), .B(n_387), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_304), .A2(n_377), .B(n_379), .Y(n_376) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_316), .Y(n_306) );
NAND3x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .C(n_313), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g478 ( .A(n_309), .B(n_398), .Y(n_478) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NOR2x1_ASAP7_75t_SL g431 ( .A(n_311), .B(n_343), .Y(n_431) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g351 ( .A(n_312), .B(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_313), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_313), .B(n_422), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_313), .B(n_422), .Y(n_495) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g398 ( .A(n_315), .B(n_371), .Y(n_398) );
AND2x2_ASAP7_75t_L g318 ( .A(n_316), .B(n_319), .Y(n_318) );
AOI221x1_ASAP7_75t_SL g317 ( .A1(n_318), .A2(n_320), .B1(n_327), .B2(n_336), .C(n_340), .Y(n_317) );
AOI32xp33_ASAP7_75t_L g499 ( .A1(n_319), .A2(n_500), .A3(n_505), .B1(n_506), .B2(n_508), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_324), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_324), .B(n_478), .Y(n_477) );
BUFx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g338 ( .A(n_326), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_326), .Y(n_342) );
OR2x2_ASAP7_75t_L g455 ( .A(n_326), .B(n_456), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g327 ( .A(n_328), .B(n_333), .C(n_335), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g377 ( .A(n_330), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g394 ( .A(n_330), .B(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_333), .A2(n_430), .B1(n_432), .B2(n_433), .Y(n_429) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g507 ( .A(n_337), .Y(n_507) );
INVx2_ASAP7_75t_L g352 ( .A(n_339), .Y(n_352) );
OAI21xp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B(n_348), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g476 ( .A(n_345), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_346), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B1(n_353), .B2(n_355), .Y(n_348) );
AND2x4_ASAP7_75t_L g445 ( .A(n_351), .B(n_360), .Y(n_445) );
INVx1_ASAP7_75t_L g504 ( .A(n_352), .Y(n_504) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g383 ( .A(n_356), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_356), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_356), .B(n_384), .Y(n_475) );
AOI211x1_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_364), .B(n_366), .C(n_392), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OR3x2_ASAP7_75t_L g467 ( .A(n_360), .B(n_362), .C(n_363), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_361), .A2(n_383), .B1(n_385), .B2(n_388), .Y(n_382) );
NOR2x1p5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g500 ( .A1(n_362), .A2(n_501), .B1(n_502), .B2(n_503), .Y(n_500) );
INVx2_ASAP7_75t_L g384 ( .A(n_365), .Y(n_384) );
OAI211xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_372), .B(n_376), .C(n_382), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_374), .B(n_378), .Y(n_389) );
INVx1_ASAP7_75t_L g416 ( .A(n_374), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_374), .B(n_481), .Y(n_489) );
OAI32xp33_ASAP7_75t_L g464 ( .A1(n_375), .A2(n_420), .A3(n_465), .B1(n_467), .B2(n_468), .Y(n_464) );
INVx1_ASAP7_75t_L g481 ( .A(n_375), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_375), .B(n_395), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g447 ( .A(n_378), .B(n_412), .Y(n_447) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g425 ( .A(n_384), .B(n_410), .Y(n_425) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g434 ( .A(n_387), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g402 ( .A(n_390), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_401), .B2(n_403), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g440 ( .A(n_397), .Y(n_440) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g421 ( .A(n_398), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_398), .B(n_405), .Y(n_509) );
INVx1_ASAP7_75t_SL g435 ( .A(n_399), .Y(n_435) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx3_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
NOR3xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_429), .C(n_436), .Y(n_406) );
OAI21xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_420), .B(n_424), .Y(n_407) );
NOR2xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_413), .Y(n_408) );
INVxp67_ASAP7_75t_L g441 ( .A(n_409), .Y(n_441) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_416), .C(n_417), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g428 ( .A(n_422), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g437 ( .A(n_425), .Y(n_437) );
OAI221xp5_ASAP7_75t_L g480 ( .A1(n_430), .A2(n_481), .B1(n_482), .B2(n_485), .C(n_486), .Y(n_480) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI32xp33_ASAP7_75t_L g436 ( .A1(n_433), .A2(n_437), .A3(n_438), .B1(n_439), .B2(n_441), .Y(n_436) );
INVx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OAI221xp5_ASAP7_75t_L g448 ( .A1(n_439), .A2(n_449), .B1(n_450), .B2(n_451), .C(n_457), .Y(n_448) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND3xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_461), .C(n_479), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_446), .B(n_448), .Y(n_443) );
AOI211x1_ASAP7_75t_L g461 ( .A1(n_444), .A2(n_462), .B(n_464), .C(n_471), .Y(n_461) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NOR2x1_ASAP7_75t_SL g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g463 ( .A(n_454), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AO21x1_ASAP7_75t_L g471 ( .A1(n_460), .A2(n_472), .B(n_474), .Y(n_471) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVxp67_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g505 ( .A(n_476), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g479 ( .A(n_480), .B(n_492), .Y(n_479) );
INVx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI21xp33_ASAP7_75t_SL g486 ( .A1(n_487), .A2(n_488), .B(n_490), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_496), .Y(n_493) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
INVx1_ASAP7_75t_L g502 ( .A(n_501), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND4xp75_ASAP7_75t_L g511 ( .A(n_512), .B(n_661), .C(n_737), .D(n_789), .Y(n_511) );
AND3x1_ASAP7_75t_L g512 ( .A(n_513), .B(n_634), .C(n_647), .Y(n_512) );
AOI221x1_ASAP7_75t_SL g513 ( .A1(n_514), .A2(n_566), .B1(n_595), .B2(n_599), .C(n_611), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g634 ( .A1(n_514), .A2(n_635), .B(n_637), .C(n_638), .Y(n_634) );
AND2x4_ASAP7_75t_L g514 ( .A(n_515), .B(n_529), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx2_ASAP7_75t_L g598 ( .A(n_518), .Y(n_598) );
BUFx2_ASAP7_75t_L g616 ( .A(n_518), .Y(n_616) );
OR2x2_ASAP7_75t_L g658 ( .A(n_518), .B(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g665 ( .A(n_518), .B(n_532), .Y(n_665) );
AND2x4_ASAP7_75t_L g700 ( .A(n_518), .B(n_531), .Y(n_700) );
OR2x2_ASAP7_75t_L g743 ( .A(n_518), .B(n_559), .Y(n_743) );
AO31x2_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .A3(n_525), .B(n_527), .Y(n_518) );
AO31x2_ASAP7_75t_L g587 ( .A1(n_525), .A2(n_588), .A3(n_589), .B(n_593), .Y(n_587) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_SL g556 ( .A(n_526), .Y(n_556) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_544), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_531), .B(n_614), .Y(n_613) );
HB1xp67_ASAP7_75t_L g630 ( .A(n_531), .Y(n_630) );
INVx2_ASAP7_75t_L g657 ( .A(n_531), .Y(n_657) );
INVx3_ASAP7_75t_L g670 ( .A(n_531), .Y(n_670) );
AND2x2_ASAP7_75t_L g788 ( .A(n_531), .B(n_617), .Y(n_788) );
INVx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g597 ( .A(n_532), .B(n_598), .Y(n_597) );
BUFx2_ASAP7_75t_L g653 ( .A(n_532), .Y(n_653) );
AO31x2_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .A3(n_541), .B(n_542), .Y(n_532) );
AO31x2_ASAP7_75t_L g604 ( .A1(n_541), .A2(n_588), .A3(n_605), .B(n_608), .Y(n_604) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g673 ( .A(n_545), .Y(n_673) );
INVx1_ASAP7_75t_L g800 ( .A(n_545), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_558), .Y(n_545) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_559), .Y(n_596) );
INVx1_ASAP7_75t_L g659 ( .A(n_546), .Y(n_659) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_557), .Y(n_546) );
OAI21x1_ASAP7_75t_L g618 ( .A1(n_547), .A2(n_548), .B(n_557), .Y(n_618) );
OAI21x1_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_552), .B(n_556), .Y(n_548) );
INVx2_ASAP7_75t_L g614 ( .A(n_558), .Y(n_614) );
AND2x2_ASAP7_75t_L g666 ( .A(n_558), .B(n_617), .Y(n_666) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g628 ( .A(n_559), .Y(n_628) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_559), .Y(n_688) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_568), .A2(n_660), .B1(n_664), .B2(n_667), .Y(n_663) );
AND2x4_ASAP7_75t_L g568 ( .A(n_569), .B(n_577), .Y(n_568) );
INVx1_ASAP7_75t_L g681 ( .A(n_569), .Y(n_681) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g601 ( .A(n_570), .B(n_579), .Y(n_601) );
AND2x2_ASAP7_75t_L g632 ( .A(n_570), .B(n_587), .Y(n_632) );
INVx4_ASAP7_75t_SL g643 ( .A(n_570), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_570), .B(n_677), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_570), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g714 ( .A(n_578), .B(n_692), .Y(n_714) );
OR2x2_ASAP7_75t_L g747 ( .A(n_578), .B(n_729), .Y(n_747) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_587), .Y(n_578) );
INVx2_ASAP7_75t_L g621 ( .A(n_579), .Y(n_621) );
INVx1_ASAP7_75t_L g626 ( .A(n_579), .Y(n_626) );
AND2x2_ASAP7_75t_L g633 ( .A(n_579), .B(n_603), .Y(n_633) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_579), .Y(n_649) );
INVx1_ASAP7_75t_L g677 ( .A(n_579), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_579), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g610 ( .A(n_587), .Y(n_610) );
AND2x4_ASAP7_75t_L g620 ( .A(n_587), .B(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g646 ( .A(n_587), .Y(n_646) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_587), .Y(n_723) );
INVx1_ASAP7_75t_L g816 ( .A(n_587), .Y(n_816) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_596), .B(n_669), .Y(n_736) );
AND2x2_ASAP7_75t_L g749 ( .A(n_596), .B(n_665), .Y(n_749) );
AND2x2_ASAP7_75t_L g819 ( .A(n_596), .B(n_670), .Y(n_819) );
AND2x4_ASAP7_75t_L g654 ( .A(n_598), .B(n_617), .Y(n_654) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g721 ( .A(n_601), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g735 ( .A(n_601), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_601), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g637 ( .A(n_602), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_602), .B(n_675), .Y(n_674) );
AOI211xp5_ASAP7_75t_L g731 ( .A1(n_602), .A2(n_732), .B(n_735), .C(n_736), .Y(n_731) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_610), .Y(n_602) );
AND2x2_ASAP7_75t_L g702 ( .A(n_603), .B(n_643), .Y(n_702) );
INVx3_ASAP7_75t_L g729 ( .A(n_603), .Y(n_729) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g624 ( .A(n_604), .Y(n_624) );
AND2x4_ASAP7_75t_L g650 ( .A(n_604), .B(n_610), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g746 ( .A(n_610), .B(n_643), .Y(n_746) );
OAI22xp5_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_619), .B1(n_627), .B2(n_631), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
INVx1_ASAP7_75t_L g768 ( .A(n_613), .Y(n_768) );
AND2x4_ASAP7_75t_L g679 ( .A(n_614), .B(n_659), .Y(n_679) );
INVx1_ASAP7_75t_L g699 ( .A(n_614), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_616), .A2(n_672), .B1(n_682), .B2(n_684), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_616), .B(n_673), .Y(n_730) );
NAND2x1_ASAP7_75t_L g787 ( .A(n_616), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g802 ( .A(n_616), .Y(n_802) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g741 ( .A(n_618), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g660 ( .A(n_620), .B(n_642), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_620), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g701 ( .A(n_620), .B(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_620), .Y(n_775) );
NAND2x1p5_ASAP7_75t_L g782 ( .A(n_620), .B(n_683), .Y(n_782) );
AND2x4_ASAP7_75t_L g805 ( .A(n_620), .B(n_733), .Y(n_805) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx3_ASAP7_75t_L g683 ( .A(n_623), .Y(n_683) );
AND2x2_ASAP7_75t_L g695 ( .A(n_623), .B(n_688), .Y(n_695) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g645 ( .A(n_624), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g693 ( .A(n_624), .Y(n_693) );
INVx1_ASAP7_75t_L g636 ( .A(n_625), .Y(n_636) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g793 ( .A(n_626), .B(n_643), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
AND2x2_ASAP7_75t_L g719 ( .A(n_628), .B(n_700), .Y(n_719) );
INVx2_ASAP7_75t_L g760 ( .A(n_628), .Y(n_760) );
AND2x4_ASAP7_75t_L g761 ( .A(n_628), .B(n_654), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_629), .B(n_679), .Y(n_809) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_632), .B(n_692), .Y(n_691) );
AND2x4_ASAP7_75t_L g704 ( .A(n_632), .B(n_649), .Y(n_704) );
INVx1_ASAP7_75t_L g796 ( .A(n_632), .Y(n_796) );
AND2x2_ASAP7_75t_L g795 ( .A(n_633), .B(n_722), .Y(n_795) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI22xp33_ASAP7_75t_L g766 ( .A1(n_637), .A2(n_767), .B1(n_769), .B2(n_771), .Y(n_766) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_641), .B(n_644), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AND2x4_ASAP7_75t_L g675 ( .A(n_643), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g711 ( .A(n_643), .Y(n_711) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_643), .Y(n_717) );
INVx2_ASAP7_75t_L g734 ( .A(n_643), .Y(n_734) );
OR2x2_ASAP7_75t_L g755 ( .A(n_643), .B(n_718), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_643), .B(n_713), .Y(n_765) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g732 ( .A(n_645), .B(n_733), .Y(n_732) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_645), .Y(n_786) );
INVx1_ASAP7_75t_L g713 ( .A(n_646), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B(n_655), .Y(n_647) );
AND2x4_ASAP7_75t_L g648 ( .A(n_649), .B(n_650), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_650), .B(n_681), .Y(n_680) );
INVx3_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
AND2x2_ASAP7_75t_L g792 ( .A(n_650), .B(n_793), .Y(n_792) );
AOI211x1_ASAP7_75t_SL g720 ( .A1(n_651), .A2(n_721), .B(n_724), .C(n_731), .Y(n_720) );
AND2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x4_ASAP7_75t_L g777 ( .A(n_653), .B(n_654), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_654), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g770 ( .A(n_654), .Y(n_770) );
AND2x2_ASAP7_75t_L g655 ( .A(n_656), .B(n_660), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx1_ASAP7_75t_L g685 ( .A(n_657), .Y(n_685) );
NOR2x1p5_ASAP7_75t_L g742 ( .A(n_657), .B(n_743), .Y(n_742) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_658), .B(n_687), .Y(n_686) );
NOR2xp67_ASAP7_75t_SL g759 ( .A(n_658), .B(n_760), .Y(n_759) );
AND2x2_ASAP7_75t_L g820 ( .A(n_660), .B(n_728), .Y(n_820) );
NOR2x1_ASAP7_75t_L g661 ( .A(n_662), .B(n_705), .Y(n_661) );
NAND3xp33_ASAP7_75t_SL g662 ( .A(n_663), .B(n_671), .C(n_689), .Y(n_662) );
AND2x2_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_665), .Y(n_696) );
AND2x2_ASAP7_75t_L g703 ( .A(n_665), .B(n_699), .Y(n_703) );
AND2x4_ASAP7_75t_SL g817 ( .A(n_665), .B(n_679), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_666), .B(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OAI22xp5_ASAP7_75t_L g781 ( .A1(n_668), .A2(n_710), .B1(n_782), .B2(n_783), .Y(n_781) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g799 ( .A(n_670), .B(n_800), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B1(n_678), .B2(n_680), .Y(n_672) );
NAND2x1_ASAP7_75t_L g748 ( .A(n_675), .B(n_728), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g758 ( .A(n_675), .B(n_722), .Y(n_758) );
INVx1_ASAP7_75t_L g785 ( .A(n_675), .Y(n_785) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OAI21xp5_ASAP7_75t_L g803 ( .A1(n_678), .A2(n_804), .B(n_807), .Y(n_803) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI21xp5_ASAP7_75t_L g690 ( .A1(n_679), .A2(n_691), .B(n_694), .Y(n_690) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx2_ASAP7_75t_L g764 ( .A(n_683), .Y(n_764) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
INVx1_ASAP7_75t_L g708 ( .A(n_686), .Y(n_708) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AOI222xp33_ASAP7_75t_L g689 ( .A1(n_690), .A2(n_696), .B1(n_697), .B2(n_701), .C1(n_703), .C2(n_704), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g724 ( .A1(n_691), .A2(n_725), .B(n_730), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_692), .B(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g806 ( .A(n_692), .Y(n_806) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_693), .Y(n_812) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_700), .Y(n_697) );
AND2x2_ASAP7_75t_L g776 ( .A(n_698), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OR2x2_ASAP7_75t_L g769 ( .A(n_699), .B(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_720), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_709), .B1(n_715), .B2(n_719), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_714), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_L g726 ( .A(n_712), .Y(n_726) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx4_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OR2x2_ASAP7_75t_L g754 ( .A(n_729), .B(n_746), .Y(n_754) );
OR2x2_ASAP7_75t_L g814 ( .A(n_729), .B(n_815), .Y(n_814) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND5xp2_ASAP7_75t_L g790 ( .A(n_735), .B(n_782), .C(n_791), .D(n_794), .E(n_796), .Y(n_790) );
NOR2x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_773), .Y(n_737) );
NAND2xp67_ASAP7_75t_SL g738 ( .A(n_739), .B(n_756), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_744), .B1(n_749), .B2(n_750), .Y(n_739) );
AND2x2_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
NAND3xp33_ASAP7_75t_SL g744 ( .A(n_745), .B(n_747), .C(n_748), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g779 ( .A(n_748), .Y(n_779) );
NAND3xp33_ASAP7_75t_SL g750 ( .A(n_751), .B(n_754), .C(n_755), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g772 ( .A(n_753), .Y(n_772) );
O2A1O1Ixp33_ASAP7_75t_SL g784 ( .A1(n_754), .A2(n_785), .B(n_786), .C(n_787), .Y(n_784) );
AOI221xp5_ASAP7_75t_L g756 ( .A1(n_757), .A2(n_759), .B1(n_761), .B2(n_762), .C(n_766), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_763), .B(n_811), .Y(n_810) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_765), .Y(n_763) );
INVx1_ASAP7_75t_L g780 ( .A(n_767), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g783 ( .A(n_777), .Y(n_783) );
AOI211xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_781), .C(n_784), .Y(n_778) );
AOI211x1_ASAP7_75t_L g789 ( .A1(n_790), .A2(n_797), .B(n_803), .C(n_818), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2x1p5_ASAP7_75t_L g798 ( .A(n_799), .B(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2x1_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_808), .A2(n_810), .B1(n_813), .B2(n_817), .Y(n_807) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
AND2x2_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_828), .B(n_831), .Y(n_821) );
INVx5_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_827), .Y(n_849) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_839), .B2(n_844), .Y(n_831) );
INVx6_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
BUFx10_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx4_ASAP7_75t_SL g839 ( .A(n_840), .Y(n_839) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
CKINVDCx11_ASAP7_75t_R g841 ( .A(n_842), .Y(n_841) );
BUFx6f_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVxp67_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
NOR2x1_ASAP7_75t_R g845 ( .A(n_846), .B(n_847), .Y(n_845) );
INVx4_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
NAND2xp5_ASAP7_75t_L g857 ( .A(n_849), .B(n_858), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_850), .B(n_860), .Y(n_859) );
BUFx12f_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
BUFx8_ASAP7_75t_SL g864 ( .A(n_852), .Y(n_864) );
BUFx12f_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
NOR2x1p5_ASAP7_75t_L g853 ( .A(n_854), .B(n_857), .Y(n_853) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_855), .B(n_856), .Y(n_854) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_864), .Y(n_862) );
endmodule