module real_jpeg_16391_n_29 (n_17, n_8, n_0, n_21, n_2, n_185, n_180, n_10, n_175, n_9, n_178, n_12, n_24, n_176, n_6, n_28, n_183, n_177, n_179, n_23, n_11, n_14, n_172, n_25, n_7, n_22, n_18, n_3, n_174, n_5, n_4, n_173, n_181, n_1, n_26, n_27, n_20, n_19, n_182, n_184, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_2;
input n_185;
input n_180;
input n_10;
input n_175;
input n_9;
input n_178;
input n_12;
input n_24;
input n_176;
input n_6;
input n_28;
input n_183;
input n_177;
input n_179;
input n_23;
input n_11;
input n_14;
input n_172;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_174;
input n_5;
input n_4;
input n_173;
input n_181;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_182;
input n_184;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_0),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_0),
.B(n_54),
.Y(n_157)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_1),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_SL g136 ( 
.A1(n_1),
.A2(n_88),
.A3(n_101),
.B1(n_104),
.B2(n_137),
.C1(n_139),
.C2(n_183),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_2),
.B(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_4),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_5),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_43),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_83),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_8),
.B(n_134),
.CON(n_133),
.SN(n_133)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_9),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g107 ( 
.A(n_10),
.B(n_108),
.C(n_130),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_11),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_12),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_12),
.B(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_13),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_41),
.C(n_168),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_16),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_17),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_17),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_18),
.Y(n_169)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_19),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_20),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_22),
.B(n_76),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_24),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_26),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_27),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_27),
.B(n_112),
.C(n_118),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_28),
.A2(n_110),
.B(n_120),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_28),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_40),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_35),
.B(n_169),
.Y(n_168)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_46),
.C(n_167),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_160),
.B(n_166),
.Y(n_46)
);

OAI31xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_72),
.A3(n_142),
.B(n_146),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_59),
.C(n_65),
.Y(n_48)
);

AOI321xp33_ASAP7_75t_L g146 ( 
.A1(n_49),
.A2(n_59),
.A3(n_147),
.B1(n_148),
.B2(n_151),
.C(n_184),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_53),
.Y(n_49)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_50),
.A2(n_60),
.A3(n_152),
.B1(n_157),
.B2(n_158),
.C1(n_159),
.C2(n_185),
.Y(n_151)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_51),
.Y(n_158)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_53),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_56),
.B(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_58),
.Y(n_115)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_61),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_65),
.B(n_153),
.C(n_154),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_71),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_71),
.Y(n_147)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI31xp67_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_81),
.A3(n_107),
.B(n_132),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_87),
.C(n_96),
.Y(n_81)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_82),
.B(n_98),
.C(n_138),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_85),
.B(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

OAI321xp33_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_96),
.A3(n_133),
.B1(n_135),
.B2(n_136),
.C(n_182),
.Y(n_132)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_101),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_105),
.B(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_126),
.C(n_127),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_116),
.C(n_117),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_133),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_165),
.Y(n_166)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_172),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_173),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_174),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_175),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_176),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_177),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_178),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_179),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_180),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_181),
.Y(n_131)
);


endmodule