module fake_jpeg_9694_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_5),
.B(n_4),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_10),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_20),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_28),
.A2(n_22),
.B1(n_21),
.B2(n_11),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_10),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_16),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_36),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_46),
.C(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_39),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_37),
.A2(n_8),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_42),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_48),
.A2(n_49),
.B1(n_37),
.B2(n_42),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_51),
.B(n_1),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_26),
.B1(n_17),
.B2(n_19),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_51),
.B(n_4),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_2),
.Y(n_55)
);


endmodule