module real_jpeg_11222_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_153;
wire n_64;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_0),
.A2(n_1),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_0),
.A2(n_48),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_1),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_1),
.B(n_43),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_1),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_21),
.B1(n_24),
.B2(n_30),
.Y(n_32)
);

AOI21xp33_ASAP7_75t_L g92 ( 
.A1(n_4),
.A2(n_9),
.B(n_21),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_6),
.B1(n_34),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_46),
.B(n_51),
.C(n_54),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g54 ( 
.A(n_5),
.B(n_46),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g114 ( 
.A1(n_5),
.A2(n_6),
.A3(n_46),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g29 ( 
.A1(n_6),
.A2(n_30),
.B(n_31),
.C(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_6),
.B(n_30),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_6),
.A2(n_9),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_6),
.A2(n_30),
.B(n_35),
.C(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_7),
.Y(n_43)
);

HAxp5_ASAP7_75t_SL g48 ( 
.A(n_7),
.B(n_35),
.CON(n_48),
.SN(n_48)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_21),
.B1(n_24),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_9),
.A2(n_46),
.B(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_9),
.B(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_9),
.A2(n_21),
.B1(n_24),
.B2(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_9),
.B(n_132),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_10),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_82),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_81),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_74),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_74),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_37),
.B1(n_63),
.B2(n_64),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_17),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_28),
.B2(n_36),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_26),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_61),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_20),
.A2(n_22),
.B(n_61),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_22),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_22),
.B(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_24),
.B(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_28),
.A2(n_36),
.B1(n_60),
.B2(n_77),
.Y(n_76)
);

AOI211xp5_ASAP7_75t_SL g79 ( 
.A1(n_28),
.A2(n_57),
.B(n_73),
.C(n_80),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_28),
.A2(n_36),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_28),
.A2(n_36),
.B1(n_91),
.B2(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_28),
.B(n_72),
.C(n_95),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_28),
.A2(n_36),
.B1(n_49),
.B2(n_58),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_28),
.A2(n_36),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_28),
.B(n_126),
.C(n_135),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_32),
.B(n_35),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_34),
.B(n_52),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_36),
.B(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_36),
.B(n_91),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_36),
.A2(n_58),
.B(n_120),
.C(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_59),
.B2(n_62),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_38),
.A2(n_39),
.B1(n_67),
.B2(n_68),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_58),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_40),
.A2(n_57),
.B1(n_118),
.B2(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_45),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_49),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_49),
.A2(n_58),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_49),
.B(n_72),
.C(n_130),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_55),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_59),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_60),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_73),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_72),
.B1(n_97),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_69),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_72),
.A2(n_94),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_72),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_72),
.B(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_72),
.A2(n_97),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_72),
.A2(n_97),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_72),
.B(n_114),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.C(n_78),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_75),
.B(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_76),
.Y(n_155)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_83),
.B(n_156),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_151),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_138),
.B(n_150),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_122),
.B(n_137),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_110),
.B(n_121),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_99),
.B(n_109),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_93),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_94),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_97),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_106),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_112),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_118),
.B1(n_119),
.B2(n_120),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_113),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_125),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_133),
.B2(n_134),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_139),
.B(n_140),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_141),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_146),
.C(n_147),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);


endmodule