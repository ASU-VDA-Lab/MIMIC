module fake_aes_10666_n_664 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_664);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_664;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g89 ( .A(n_88), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_82), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_16), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_29), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_44), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_43), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_0), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_76), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_52), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_8), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
BUFx8_ASAP7_75t_SL g100 ( .A(n_20), .Y(n_100) );
INVx1_ASAP7_75t_SL g101 ( .A(n_57), .Y(n_101) );
BUFx10_ASAP7_75t_L g102 ( .A(n_1), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_39), .Y(n_104) );
BUFx5_ASAP7_75t_L g105 ( .A(n_54), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_58), .Y(n_106) );
INVx4_ASAP7_75t_R g107 ( .A(n_46), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_21), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_64), .Y(n_110) );
BUFx2_ASAP7_75t_SL g111 ( .A(n_9), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_22), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_17), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_77), .Y(n_116) );
INVxp33_ASAP7_75t_L g117 ( .A(n_10), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_83), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_32), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_6), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_66), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_19), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_68), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_10), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_86), .Y(n_127) );
INVxp67_ASAP7_75t_SL g128 ( .A(n_27), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_87), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_100), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_105), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_100), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_117), .B(n_0), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_114), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_114), .B(n_1), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_117), .B(n_3), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_104), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_105), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_121), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_94), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_91), .B(n_3), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_96), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_99), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_105), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_104), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_108), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_106), .B(n_4), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_110), .B(n_4), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_95), .B(n_5), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_112), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_98), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_98), .B(n_5), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_131), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_136), .B(n_93), .Y(n_159) );
BUFx3_ASAP7_75t_L g160 ( .A(n_138), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_157), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_136), .B(n_92), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_140), .B(n_120), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_157), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_140), .B(n_122), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_142), .B(n_92), .Y(n_169) );
BUFx3_ASAP7_75t_L g170 ( .A(n_138), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_142), .B(n_97), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_139), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVxp33_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_138), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_147), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_145), .B(n_108), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_145), .B(n_97), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_146), .B(n_123), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_155), .B(n_102), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_157), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
AND3x4_ASAP7_75t_L g186 ( .A(n_135), .B(n_113), .C(n_126), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_150), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_150), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_146), .B(n_124), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_148), .B(n_125), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_148), .B(n_127), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_179), .B(n_133), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_187), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g194 ( .A1(n_186), .A2(n_133), .B1(n_137), .B2(n_135), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_181), .B(n_137), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_159), .B(n_154), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_165), .Y(n_197) );
OAI22xp5_ASAP7_75t_SL g198 ( .A1(n_186), .A2(n_126), .B1(n_130), .B2(n_132), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_182), .B(n_135), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_185), .B(n_123), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_165), .Y(n_201) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_186), .A2(n_156), .B1(n_154), .B2(n_152), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_182), .B(n_175), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_161), .B(n_180), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_187), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_161), .B(n_156), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_185), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_188), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_163), .Y(n_209) );
NOR3xp33_ASAP7_75t_L g210 ( .A(n_169), .B(n_153), .C(n_144), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_185), .Y(n_211) );
NOR2xp33_ASAP7_75t_R g212 ( .A(n_167), .B(n_119), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_185), .Y(n_213) );
AOI22xp5_ASAP7_75t_L g214 ( .A1(n_167), .A2(n_151), .B1(n_119), .B2(n_118), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_161), .B(n_150), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_167), .B(n_113), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_167), .A2(n_128), .B(n_129), .Y(n_217) );
HB1xp67_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_171), .Y(n_219) );
BUFx8_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_160), .Y(n_221) );
BUFx4f_ASAP7_75t_L g222 ( .A(n_183), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_161), .B(n_150), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_180), .B(n_101), .Y(n_226) );
BUFx2_ASAP7_75t_L g227 ( .A(n_180), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_189), .B(n_102), .Y(n_228) );
INVx2_ASAP7_75t_SL g229 ( .A(n_189), .Y(n_229) );
AND2x6_ASAP7_75t_L g230 ( .A(n_183), .B(n_190), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_134), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_190), .B(n_109), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_160), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_178), .B(n_115), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_164), .B(n_134), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_168), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_223), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_201), .B(n_191), .Y(n_238) );
INVx6_ASAP7_75t_L g239 ( .A(n_220), .Y(n_239) );
BUFx12f_ASAP7_75t_L g240 ( .A(n_220), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_229), .B(n_162), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_207), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_194), .A2(n_162), .B(n_177), .C(n_172), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_194), .A2(n_172), .B1(n_177), .B2(n_174), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_196), .A2(n_174), .B(n_158), .C(n_184), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_202), .A2(n_218), .B1(n_199), .B2(n_230), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_234), .B(n_184), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_198), .B(n_111), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_198), .B(n_111), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_204), .A2(n_184), .B(n_158), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_SL g253 ( .A1(n_231), .A2(n_158), .B(n_173), .C(n_166), .Y(n_253) );
INVx4_ASAP7_75t_L g254 ( .A(n_207), .Y(n_254) );
BUFx3_ASAP7_75t_L g255 ( .A(n_197), .Y(n_255) );
BUFx4f_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_206), .A2(n_173), .B(n_166), .Y(n_257) );
INVx4_ASAP7_75t_L g258 ( .A(n_207), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_234), .B(n_173), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_233), .Y(n_260) );
NOR2xp67_ASAP7_75t_L g261 ( .A(n_202), .B(n_6), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_192), .A2(n_166), .B(n_170), .C(n_160), .Y(n_262) );
O2A1O1Ixp5_ASAP7_75t_SL g263 ( .A1(n_232), .A2(n_176), .B(n_107), .C(n_149), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_215), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_224), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_228), .B(n_102), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_236), .B(n_7), .Y(n_267) );
AOI21x1_ASAP7_75t_L g268 ( .A1(n_226), .A2(n_170), .B(n_176), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_233), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_212), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_199), .B(n_7), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
OAI22xp5_ASAP7_75t_SL g273 ( .A1(n_219), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_214), .B(n_11), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_222), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_205), .Y(n_276) );
BUFx12f_ASAP7_75t_L g277 ( .A(n_209), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_208), .Y(n_278) );
O2A1O1Ixp5_ASAP7_75t_L g279 ( .A1(n_217), .A2(n_170), .B(n_176), .C(n_149), .Y(n_279) );
AOI22x1_ASAP7_75t_L g280 ( .A1(n_221), .A2(n_176), .B1(n_149), .B2(n_138), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_253), .A2(n_195), .B(n_235), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
BUFx4f_ASAP7_75t_SL g283 ( .A(n_240), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_262), .A2(n_200), .B(n_210), .Y(n_284) );
INVx4_ASAP7_75t_L g285 ( .A(n_260), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_263), .A2(n_216), .B(n_214), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_239), .Y(n_287) );
AND2x4_ASAP7_75t_L g288 ( .A(n_264), .B(n_211), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_260), .Y(n_289) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_239), .Y(n_290) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_253), .A2(n_176), .B(n_230), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_261), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_268), .A2(n_216), .B(n_230), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_260), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_265), .B(n_213), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_279), .A2(n_216), .B(n_230), .Y(n_296) );
BUFx12f_ASAP7_75t_L g297 ( .A(n_239), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_279), .A2(n_216), .B(n_105), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_260), .Y(n_299) );
OAI221xp5_ASAP7_75t_L g300 ( .A1(n_247), .A2(n_222), .B1(n_227), .B2(n_213), .C(n_149), .Y(n_300) );
OAI21x1_ASAP7_75t_L g301 ( .A1(n_280), .A2(n_105), .B(n_176), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_233), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_269), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_247), .B(n_105), .Y(n_304) );
INVx3_ASAP7_75t_L g305 ( .A(n_269), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_251), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_254), .B(n_149), .Y(n_307) );
OAI221xp5_ASAP7_75t_L g308 ( .A1(n_243), .A2(n_138), .B1(n_13), .B2(n_14), .C(n_15), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_277), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_276), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_278), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_257), .A2(n_50), .B(n_84), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_237), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_252), .A2(n_49), .B(n_81), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_243), .A2(n_12), .B(n_13), .C(n_14), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_242), .A2(n_53), .B(n_18), .Y(n_316) );
OAI22xp33_ASAP7_75t_L g317 ( .A1(n_292), .A2(n_249), .B1(n_250), .B2(n_270), .Y(n_317) );
AOI221xp5_ASAP7_75t_L g318 ( .A1(n_292), .A2(n_266), .B1(n_271), .B2(n_267), .C(n_238), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_294), .Y(n_319) );
INVx4_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
BUFx4f_ASAP7_75t_L g321 ( .A(n_297), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g322 ( .A1(n_304), .A2(n_249), .B1(n_250), .B2(n_271), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_306), .Y(n_323) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_291), .A2(n_262), .B(n_246), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_294), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_306), .B(n_249), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_310), .Y(n_327) );
INVx6_ASAP7_75t_L g328 ( .A(n_297), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_302), .B(n_250), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_310), .B(n_267), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_311), .B(n_245), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_311), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_313), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_283), .Y(n_334) );
AND2x4_ASAP7_75t_L g335 ( .A(n_288), .B(n_275), .Y(n_335) );
AOI21xp33_ASAP7_75t_L g336 ( .A1(n_300), .A2(n_270), .B(n_248), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_294), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g339 ( .A1(n_315), .A2(n_244), .B(n_241), .C(n_259), .Y(n_339) );
INVxp67_ASAP7_75t_L g340 ( .A(n_282), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_285), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_302), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g343 ( .A1(n_281), .A2(n_246), .B(n_241), .Y(n_343) );
OAI221xp5_ASAP7_75t_L g344 ( .A1(n_308), .A2(n_256), .B1(n_273), .B2(n_272), .C(n_242), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_304), .B(n_272), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_342), .B(n_284), .Y(n_346) );
AND2x4_ASAP7_75t_L g347 ( .A(n_341), .B(n_285), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_319), .Y(n_348) );
INVx2_ASAP7_75t_SL g349 ( .A(n_321), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_331), .B(n_284), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_327), .B(n_281), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_332), .B(n_284), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_333), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_338), .B(n_345), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_345), .B(n_284), .Y(n_357) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_341), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_331), .B(n_285), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_325), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_329), .B(n_285), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_329), .B(n_315), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_341), .B(n_289), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_324), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_329), .B(n_295), .Y(n_367) );
INVx6_ASAP7_75t_L g368 ( .A(n_320), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_325), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_321), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_295), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_348), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_353), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_368), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_346), .B(n_326), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_357), .B(n_326), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_346), .B(n_337), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_351), .B(n_291), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_357), .B(n_322), .Y(n_383) );
OA21x2_ASAP7_75t_L g384 ( .A1(n_366), .A2(n_343), .B(n_298), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_291), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_354), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_352), .B(n_291), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_352), .B(n_322), .Y(n_388) );
AOI221x1_ASAP7_75t_L g389 ( .A1(n_366), .A2(n_336), .B1(n_330), .B2(n_335), .C(n_305), .Y(n_389) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_354), .A2(n_303), .B(n_294), .Y(n_390) );
INVx5_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_355), .B(n_289), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_355), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_373), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_373), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_350), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_368), .B(n_334), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_340), .Y(n_398) );
BUFx2_ASAP7_75t_L g399 ( .A(n_361), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
BUFx3_ASAP7_75t_L g402 ( .A(n_368), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_350), .B(n_289), .Y(n_403) );
AO21x2_ASAP7_75t_L g404 ( .A1(n_372), .A2(n_298), .B(n_308), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_372), .B(n_318), .C(n_344), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
INVx3_ASAP7_75t_L g407 ( .A(n_359), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_378), .B(n_361), .Y(n_409) );
INVx5_ASAP7_75t_SL g410 ( .A(n_391), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_378), .B(n_369), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_396), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_396), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_382), .B(n_364), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_382), .B(n_364), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_393), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_394), .Y(n_418) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_405), .A2(n_317), .B1(n_356), .B2(n_290), .C(n_287), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_385), .B(n_362), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_385), .B(n_362), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_380), .B(n_367), .Y(n_422) );
AND2x4_ASAP7_75t_L g423 ( .A(n_381), .B(n_387), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_391), .B(n_349), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_398), .B(n_334), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_381), .B(n_367), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_387), .B(n_371), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_396), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_386), .B(n_371), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_386), .B(n_363), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_375), .B(n_363), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_405), .A2(n_300), .B(n_349), .Y(n_432) );
NAND4xp25_ASAP7_75t_L g433 ( .A(n_398), .B(n_360), .C(n_320), .D(n_339), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_401), .Y(n_434) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_397), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_394), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_395), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_375), .B(n_359), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_380), .B(n_359), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_379), .B(n_359), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_395), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_383), .B(n_347), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_383), .B(n_347), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_379), .B(n_347), .Y(n_444) );
INVx2_ASAP7_75t_SL g445 ( .A(n_391), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_388), .B(n_347), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_401), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_388), .B(n_368), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_401), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_406), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_400), .B(n_365), .Y(n_452) );
INVx1_ASAP7_75t_SL g453 ( .A(n_377), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_406), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_406), .B(n_365), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_407), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_374), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_407), .B(n_365), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_408), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_412), .Y(n_460) );
OR2x2_ASAP7_75t_L g461 ( .A(n_409), .B(n_376), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_409), .B(n_376), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_412), .Y(n_463) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_457), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_417), .B(n_374), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_427), .B(n_399), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_427), .B(n_426), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_410), .Y(n_469) );
NAND2xp33_ASAP7_75t_SL g470 ( .A(n_445), .B(n_399), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_377), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_457), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_423), .B(n_407), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_418), .Y(n_475) );
BUFx2_ASAP7_75t_L g476 ( .A(n_435), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_436), .B(n_408), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_423), .B(n_392), .Y(n_478) );
NOR2x1_ASAP7_75t_L g479 ( .A(n_424), .B(n_402), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_436), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_423), .B(n_392), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_411), .B(n_402), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_437), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_433), .B(n_402), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_423), .B(n_403), .Y(n_485) );
NAND2x1_ASAP7_75t_L g486 ( .A(n_445), .B(n_328), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
INVx1_ASAP7_75t_SL g488 ( .A(n_435), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_425), .B(n_391), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_411), .B(n_403), .Y(n_490) );
INVx8_ASAP7_75t_L g491 ( .A(n_410), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_441), .B(n_389), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_410), .B(n_391), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_415), .B(n_391), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_415), .B(n_391), .Y(n_495) );
INVxp67_ASAP7_75t_L g496 ( .A(n_453), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_422), .B(n_390), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_441), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_416), .B(n_389), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_422), .B(n_390), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_416), .B(n_384), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_420), .B(n_365), .Y(n_502) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_432), .A2(n_404), .B(n_384), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_452), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_430), .Y(n_505) );
INVxp67_ASAP7_75t_L g506 ( .A(n_450), .Y(n_506) );
INVxp67_ASAP7_75t_L g507 ( .A(n_450), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_430), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_420), .B(n_384), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_431), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_421), .B(n_384), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g512 ( .A1(n_449), .A2(n_307), .B(n_370), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_413), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_431), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_413), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_458), .B(n_320), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_442), .B(n_404), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_414), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_SL g519 ( .A1(n_446), .A2(n_299), .B(n_305), .C(n_328), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_484), .A2(n_429), .B1(n_442), .B2(n_443), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_505), .B(n_429), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_508), .Y(n_522) );
INVx3_ASAP7_75t_SL g523 ( .A(n_491), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_510), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_514), .B(n_421), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_468), .B(n_444), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_460), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_509), .B(n_444), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_484), .A2(n_419), .B1(n_447), .B2(n_443), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_488), .B(n_358), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_491), .A2(n_410), .B1(n_458), .B2(n_455), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_464), .B(n_439), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_486), .A2(n_458), .B(n_446), .C(n_456), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_512), .A2(n_458), .B1(n_438), .B2(n_440), .Y(n_534) );
OAI32xp33_ASAP7_75t_L g535 ( .A1(n_470), .A2(n_439), .A3(n_456), .B1(n_446), .B2(n_454), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_463), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_476), .Y(n_537) );
AOI222xp33_ASAP7_75t_L g538 ( .A1(n_499), .A2(n_438), .B1(n_440), .B2(n_455), .C1(n_454), .C2(n_451), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_482), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_464), .Y(n_540) );
INVxp67_ASAP7_75t_L g541 ( .A(n_496), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_511), .B(n_459), .Y(n_542) );
AOI222xp33_ASAP7_75t_L g543 ( .A1(n_499), .A2(n_459), .B1(n_451), .B2(n_410), .C1(n_335), .C2(n_448), .Y(n_543) );
OAI21xp5_ASAP7_75t_SL g544 ( .A1(n_493), .A2(n_456), .B(n_446), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_467), .Y(n_545) );
NOR4xp25_ASAP7_75t_SL g546 ( .A(n_493), .B(n_309), .C(n_456), .D(n_328), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_489), .A2(n_448), .B1(n_434), .B2(n_428), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_489), .A2(n_434), .B1(n_428), .B2(n_414), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_461), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_471), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_504), .B(n_404), .Y(n_551) );
OAI21xp5_ASAP7_75t_L g552 ( .A1(n_470), .A2(n_316), .B(n_335), .Y(n_552) );
AOI21xp33_ASAP7_75t_L g553 ( .A1(n_479), .A2(n_15), .B(n_404), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_475), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_462), .B(n_307), .Y(n_555) );
AOI21xp33_ASAP7_75t_SL g556 ( .A1(n_491), .A2(n_316), .B(n_312), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_474), .B(n_312), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_496), .Y(n_559) );
AOI32xp33_ASAP7_75t_L g560 ( .A1(n_494), .A2(n_314), .A3(n_296), .B1(n_286), .B2(n_293), .Y(n_560) );
AOI322xp5_ASAP7_75t_L g561 ( .A1(n_466), .A2(n_288), .A3(n_295), .B1(n_305), .B2(n_299), .C1(n_286), .C2(n_314), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_490), .B(n_307), .Y(n_562) );
A2O1A1Ixp33_ASAP7_75t_SL g563 ( .A1(n_469), .A2(n_305), .B(n_299), .C(n_25), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_497), .B(n_296), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g565 ( .A1(n_501), .A2(n_293), .B(n_299), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_506), .Y(n_566) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_469), .A2(n_256), .B1(n_303), .B2(n_294), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_516), .A2(n_295), .B1(n_288), .B2(n_254), .Y(n_568) );
OAI322xp33_ASAP7_75t_L g569 ( .A1(n_500), .A2(n_258), .A3(n_303), .B1(n_294), .B2(n_269), .C1(n_30), .C2(n_31), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_483), .B(n_498), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_487), .Y(n_571) );
NAND3xp33_ASAP7_75t_L g572 ( .A(n_503), .B(n_303), .C(n_258), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_537), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_540), .Y(n_574) );
XNOR2x1_ASAP7_75t_L g575 ( .A(n_539), .B(n_516), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_570), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_566), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_527), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_532), .Y(n_579) );
NOR2xp33_ASAP7_75t_SL g580 ( .A(n_523), .B(n_495), .Y(n_580) );
XNOR2x1_ASAP7_75t_L g581 ( .A(n_529), .B(n_472), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_530), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_538), .B(n_501), .Y(n_583) );
INVx2_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
AOI31xp33_ASAP7_75t_SL g585 ( .A1(n_543), .A2(n_517), .A3(n_503), .B(n_506), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_544), .A2(n_519), .B(n_502), .C(n_481), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_522), .B(n_473), .Y(n_587) );
BUFx2_ASAP7_75t_L g588 ( .A(n_541), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_524), .B(n_507), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_562), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_559), .A2(n_507), .B1(n_465), .B2(n_492), .C(n_478), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_545), .Y(n_592) );
AOI221xp5_ASAP7_75t_L g593 ( .A1(n_520), .A2(n_465), .B1(n_492), .B2(n_485), .C(n_477), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_550), .Y(n_594) );
OAI22xp33_ASAP7_75t_SL g595 ( .A1(n_546), .A2(n_477), .B1(n_518), .B2(n_515), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_554), .Y(n_596) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_525), .B(n_513), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_557), .Y(n_598) );
HB1xp67_ASAP7_75t_L g599 ( .A(n_542), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_571), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_549), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_521), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_528), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_555), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_526), .Y(n_605) );
CKINVDCx14_ASAP7_75t_R g606 ( .A(n_546), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_547), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_548), .Y(n_608) );
AOI21xp5_ASAP7_75t_L g609 ( .A1(n_606), .A2(n_535), .B(n_563), .Y(n_609) );
OAI211xp5_ASAP7_75t_L g610 ( .A1(n_606), .A2(n_531), .B(n_553), .C(n_534), .Y(n_610) );
INVxp67_ASAP7_75t_L g611 ( .A(n_588), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_584), .Y(n_612) );
INVxp67_ASAP7_75t_SL g613 ( .A(n_599), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_583), .A2(n_551), .B1(n_569), .B2(n_564), .C(n_558), .Y(n_614) );
AOI21xp5_ASAP7_75t_L g615 ( .A1(n_595), .A2(n_552), .B(n_569), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_586), .A2(n_533), .B1(n_568), .B2(n_561), .C(n_565), .Y(n_616) );
XNOR2xp5_ASAP7_75t_L g617 ( .A(n_575), .B(n_567), .Y(n_617) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_586), .A2(n_572), .B(n_556), .C(n_519), .Y(n_618) );
OAI211xp5_ASAP7_75t_L g619 ( .A1(n_593), .A2(n_572), .B(n_560), .C(n_301), .Y(n_619) );
AOI21xp33_ASAP7_75t_SL g620 ( .A1(n_581), .A2(n_23), .B(n_24), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_593), .B(n_303), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_607), .A2(n_288), .B(n_301), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_599), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_608), .A2(n_303), .B(n_269), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_589), .Y(n_625) );
OAI22xp5_ASAP7_75t_L g626 ( .A1(n_582), .A2(n_26), .B1(n_28), .B2(n_33), .Y(n_626) );
OAI211xp5_ASAP7_75t_L g627 ( .A1(n_573), .A2(n_34), .B(n_35), .C(n_36), .Y(n_627) );
AND5x1_ASAP7_75t_L g628 ( .A(n_580), .B(n_38), .C(n_40), .D(n_41), .E(n_42), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_591), .A2(n_45), .B(n_47), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_591), .A2(n_51), .B(n_55), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_623), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_611), .B(n_582), .Y(n_632) );
AOI221xp5_ASAP7_75t_SL g633 ( .A1(n_615), .A2(n_590), .B1(n_577), .B2(n_585), .C(n_576), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_625), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_613), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_616), .A2(n_602), .B1(n_577), .B2(n_605), .C(n_603), .Y(n_636) );
AOI21xp33_ASAP7_75t_L g637 ( .A1(n_619), .A2(n_594), .B(n_578), .Y(n_637) );
OAI21xp33_ASAP7_75t_L g638 ( .A1(n_610), .A2(n_597), .B(n_601), .Y(n_638) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_614), .A2(n_592), .B1(n_600), .B2(n_598), .C1(n_596), .C2(n_579), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_618), .A2(n_604), .B1(n_587), .B2(n_574), .C(n_61), .Y(n_640) );
OAI211xp5_ASAP7_75t_L g641 ( .A1(n_609), .A2(n_56), .B(n_59), .C(n_60), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_617), .A2(n_63), .B1(n_65), .B2(n_67), .Y(n_642) );
OAI31xp33_ASAP7_75t_L g643 ( .A1(n_629), .A2(n_69), .A3(n_70), .B(n_71), .Y(n_643) );
AOI222xp33_ASAP7_75t_L g644 ( .A1(n_636), .A2(n_621), .B1(n_612), .B2(n_626), .C1(n_624), .C2(n_622), .Y(n_644) );
OAI221xp5_ASAP7_75t_L g645 ( .A1(n_633), .A2(n_630), .B1(n_620), .B2(n_627), .C(n_626), .Y(n_645) );
NOR2xp67_ASAP7_75t_L g646 ( .A(n_635), .B(n_72), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_634), .B(n_628), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_639), .B(n_73), .Y(n_648) );
NAND3xp33_ASAP7_75t_SL g649 ( .A(n_640), .B(n_74), .C(n_75), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_631), .Y(n_650) );
NAND4xp25_ASAP7_75t_SL g651 ( .A(n_644), .B(n_637), .C(n_640), .D(n_641), .Y(n_651) );
AO22x2_ASAP7_75t_L g652 ( .A1(n_650), .A2(n_632), .B1(n_638), .B2(n_642), .Y(n_652) );
BUFx4f_ASAP7_75t_SL g653 ( .A(n_647), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_648), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_652), .Y(n_655) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_653), .Y(n_656) );
O2A1O1Ixp33_ASAP7_75t_L g657 ( .A1(n_654), .A2(n_645), .B(n_649), .C(n_646), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_656), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_655), .A2(n_651), .B1(n_643), .B2(n_80), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_658), .A2(n_657), .B1(n_79), .B2(n_85), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
BUFx3_ASAP7_75t_L g662 ( .A(n_661), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_662), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_663), .A2(n_662), .B1(n_660), .B2(n_78), .Y(n_664) );
endmodule