module real_aes_552_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_793, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_793;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_140;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_0), .B(n_121), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g487 ( .A1(n_1), .A2(n_130), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_2), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_3), .B(n_121), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_4), .B(n_137), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_5), .B(n_137), .Y(n_532) );
INVx1_ASAP7_75t_L g128 ( .A(n_6), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_7), .B(n_137), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g459 ( .A(n_8), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_9), .B(n_139), .Y(n_480) );
AND2x2_ASAP7_75t_L g157 ( .A(n_10), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g221 ( .A(n_11), .B(n_146), .Y(n_221) );
INVx2_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
AOI221x1_ASAP7_75t_L g548 ( .A1(n_13), .A2(n_24), .B1(n_121), .B2(n_130), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_14), .B(n_137), .Y(n_193) );
CKINVDCx16_ASAP7_75t_R g447 ( .A(n_15), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_16), .B(n_121), .Y(n_476) );
AO21x2_ASAP7_75t_L g474 ( .A1(n_17), .A2(n_146), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_18), .B(n_141), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_19), .B(n_137), .Y(n_498) );
AO21x1_ASAP7_75t_L g527 ( .A1(n_20), .A2(n_121), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_21), .B(n_121), .Y(n_226) );
INVx1_ASAP7_75t_L g451 ( .A(n_22), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_23), .A2(n_90), .B1(n_121), .B2(n_163), .Y(n_162) );
NAND2x1_ASAP7_75t_L g519 ( .A(n_25), .B(n_137), .Y(n_519) );
NAND2x1_ASAP7_75t_L g508 ( .A(n_26), .B(n_139), .Y(n_508) );
OR2x2_ASAP7_75t_L g144 ( .A(n_27), .B(n_87), .Y(n_144) );
OA21x2_ASAP7_75t_L g147 ( .A1(n_27), .A2(n_87), .B(n_143), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_28), .B(n_139), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_29), .B(n_137), .Y(n_479) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_30), .A2(n_158), .B(n_189), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_31), .B(n_139), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_32), .A2(n_130), .B(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_33), .B(n_137), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_34), .A2(n_130), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g127 ( .A(n_35), .B(n_128), .Y(n_127) );
AND2x2_ASAP7_75t_L g131 ( .A(n_35), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g171 ( .A(n_35), .Y(n_171) );
OR2x6_ASAP7_75t_L g449 ( .A(n_36), .B(n_450), .Y(n_449) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_37), .B(n_121), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_38), .B(n_121), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_39), .B(n_137), .Y(n_183) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_40), .A2(n_104), .B1(n_456), .B2(n_461), .C1(n_781), .C2(n_786), .Y(n_103) );
XNOR2xp5_ASAP7_75t_L g105 ( .A(n_40), .B(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_40), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_41), .B(n_139), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_42), .B(n_121), .Y(n_120) );
XNOR2xp5_ASAP7_75t_L g768 ( .A(n_43), .B(n_769), .Y(n_768) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_44), .A2(n_130), .B(n_153), .Y(n_152) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_45), .A2(n_108), .B1(n_109), .B2(n_110), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_45), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_46), .A2(n_130), .B(n_507), .Y(n_506) );
XNOR2xp5_ASAP7_75t_L g767 ( .A(n_47), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_48), .B(n_139), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_49), .B(n_139), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_50), .B(n_121), .Y(n_190) );
INVx1_ASAP7_75t_L g124 ( .A(n_51), .Y(n_124) );
INVx1_ASAP7_75t_L g134 ( .A(n_51), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_52), .B(n_137), .Y(n_155) );
AND2x2_ASAP7_75t_L g178 ( .A(n_53), .B(n_141), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_54), .B(n_139), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_55), .B(n_137), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_56), .B(n_139), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_57), .A2(n_130), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_58), .B(n_121), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_59), .B(n_121), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_60), .A2(n_130), .B(n_199), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_61), .A2(n_99), .B1(n_770), .B2(n_771), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_61), .Y(n_771) );
AND2x2_ASAP7_75t_L g232 ( .A(n_62), .B(n_142), .Y(n_232) );
AO21x1_ASAP7_75t_L g529 ( .A1(n_63), .A2(n_130), .B(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_64), .B(n_121), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_65), .B(n_139), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g110 ( .A1(n_66), .A2(n_80), .B1(n_111), .B2(n_112), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_66), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_67), .B(n_121), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_68), .B(n_139), .Y(n_194) );
AOI22xp5_ASAP7_75t_L g168 ( .A1(n_69), .A2(n_94), .B1(n_130), .B2(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_70), .B(n_137), .Y(n_229) );
AND2x2_ASAP7_75t_L g542 ( .A(n_71), .B(n_142), .Y(n_542) );
INVx1_ASAP7_75t_L g126 ( .A(n_72), .Y(n_126) );
INVx1_ASAP7_75t_L g132 ( .A(n_72), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_73), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g511 ( .A(n_74), .B(n_158), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_75), .B(n_139), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_76), .A2(n_130), .B(n_182), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g129 ( .A1(n_77), .A2(n_130), .B(n_135), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_78), .A2(n_130), .B(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g203 ( .A(n_79), .B(n_142), .Y(n_203) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_80), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_81), .B(n_141), .Y(n_160) );
INVx1_ASAP7_75t_L g452 ( .A(n_82), .Y(n_452) );
AND2x2_ASAP7_75t_L g484 ( .A(n_83), .B(n_158), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g500 ( .A(n_84), .B(n_121), .Y(n_500) );
AND2x2_ASAP7_75t_L g145 ( .A(n_85), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g528 ( .A(n_86), .B(n_185), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_88), .B(n_139), .Y(n_499) );
AND2x2_ASAP7_75t_L g522 ( .A(n_89), .B(n_158), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_91), .B(n_137), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_92), .A2(n_130), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_93), .B(n_139), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_95), .A2(n_130), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_96), .B(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_97), .B(n_137), .Y(n_489) );
BUFx2_ASAP7_75t_L g231 ( .A(n_98), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_99), .Y(n_770) );
BUFx2_ASAP7_75t_L g460 ( .A(n_100), .Y(n_460) );
BUFx2_ASAP7_75t_SL g790 ( .A(n_100), .Y(n_790) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_101), .A2(n_130), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_102), .Y(n_778) );
OAI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_443), .B(n_453), .Y(n_104) );
XNOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_113), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
OAI22xp5_ASAP7_75t_L g463 ( .A1(n_113), .A2(n_464), .B1(n_468), .B2(n_763), .Y(n_463) );
INVx3_ASAP7_75t_SL g775 ( .A(n_113), .Y(n_775) );
AND2x4_ASAP7_75t_SL g113 ( .A(n_114), .B(n_339), .Y(n_113) );
NOR3xp33_ASAP7_75t_SL g114 ( .A(n_115), .B(n_248), .C(n_280), .Y(n_114) );
OAI221xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_174), .B1(n_204), .B2(n_222), .C(n_233), .Y(n_115) );
OR2x2_ASAP7_75t_L g116 ( .A(n_117), .B(n_148), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g210 ( .A(n_118), .B(n_149), .Y(n_210) );
INVx4_ASAP7_75t_L g239 ( .A(n_118), .Y(n_239) );
AND2x4_ASAP7_75t_SL g279 ( .A(n_118), .B(n_212), .Y(n_279) );
BUFx2_ASAP7_75t_L g289 ( .A(n_118), .Y(n_289) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_118), .B(n_294), .Y(n_355) );
AND2x2_ASAP7_75t_L g364 ( .A(n_118), .B(n_292), .Y(n_364) );
OR2x2_ASAP7_75t_L g372 ( .A(n_118), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g398 ( .A(n_118), .B(n_237), .Y(n_398) );
AND2x4_ASAP7_75t_L g417 ( .A(n_118), .B(n_418), .Y(n_417) );
OR2x6_ASAP7_75t_L g118 ( .A(n_119), .B(n_145), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_129), .B(n_141), .Y(n_119) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_127), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
AND2x6_ASAP7_75t_L g139 ( .A(n_123), .B(n_132), .Y(n_139) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x4_ASAP7_75t_L g137 ( .A(n_125), .B(n_134), .Y(n_137) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx5_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
AND2x2_ASAP7_75t_L g133 ( .A(n_128), .B(n_134), .Y(n_133) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_128), .Y(n_166) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_133), .Y(n_130) );
BUFx3_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
INVx2_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
AND2x4_ASAP7_75t_L g169 ( .A(n_133), .B(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g165 ( .A(n_134), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B(n_140), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_139), .B(n_231), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_140), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_140), .A2(n_183), .B(n_184), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_140), .A2(n_193), .B(n_194), .Y(n_192) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_140), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_140), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_140), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_140), .A2(n_479), .B(n_480), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_140), .A2(n_489), .B(n_490), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_140), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_140), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_140), .A2(n_519), .B(n_520), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_140), .A2(n_531), .B(n_532), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g538 ( .A1(n_140), .A2(n_539), .B(n_540), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_140), .A2(n_550), .B(n_551), .Y(n_549) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_141), .A2(n_162), .B(n_168), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_141), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_141), .A2(n_486), .B(n_487), .Y(n_485) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_141), .A2(n_548), .B(n_552), .Y(n_547) );
OA21x2_ASAP7_75t_L g610 ( .A1(n_141), .A2(n_548), .B(n_552), .Y(n_610) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_144), .Y(n_142) );
AND2x4_ASAP7_75t_L g185 ( .A(n_143), .B(n_144), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_146), .A2(n_226), .B(n_227), .Y(n_225) );
BUFx4f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_147), .Y(n_150) );
INVx2_ASAP7_75t_SL g330 ( .A(n_148), .Y(n_330) );
OR2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_159), .Y(n_148) );
AND2x2_ASAP7_75t_L g237 ( .A(n_149), .B(n_213), .Y(n_237) );
INVx2_ASAP7_75t_L g264 ( .A(n_149), .Y(n_264) );
INVx2_ASAP7_75t_L g294 ( .A(n_149), .Y(n_294) );
AND2x2_ASAP7_75t_L g308 ( .A(n_149), .B(n_212), .Y(n_308) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_157), .Y(n_149) );
INVx4_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_156), .Y(n_151) );
INVx3_ASAP7_75t_L g196 ( .A(n_158), .Y(n_196) );
AND2x2_ASAP7_75t_L g238 ( .A(n_159), .B(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g261 ( .A(n_159), .Y(n_261) );
BUFx3_ASAP7_75t_L g275 ( .A(n_159), .Y(n_275) );
AND2x2_ASAP7_75t_L g304 ( .A(n_159), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x4_ASAP7_75t_L g208 ( .A(n_160), .B(n_161), .Y(n_208) );
AND2x4_ASAP7_75t_L g163 ( .A(n_164), .B(n_167), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_166), .Y(n_164) );
NOR2x1p5_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx1_ASAP7_75t_L g310 ( .A(n_174), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_186), .Y(n_174) );
OR2x2_ASAP7_75t_L g421 ( .A(n_175), .B(n_222), .Y(n_421) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AND2x2_ASAP7_75t_L g277 ( .A(n_176), .B(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_176), .B(n_186), .Y(n_338) );
OR2x2_ASAP7_75t_L g436 ( .A(n_176), .B(n_358), .Y(n_436) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g247 ( .A(n_177), .B(n_223), .Y(n_247) );
OR2x2_ASAP7_75t_SL g257 ( .A(n_177), .B(n_258), .Y(n_257) );
INVx4_ASAP7_75t_L g268 ( .A(n_177), .Y(n_268) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_177), .Y(n_319) );
NAND2x1_ASAP7_75t_L g325 ( .A(n_177), .B(n_224), .Y(n_325) );
AND2x2_ASAP7_75t_L g350 ( .A(n_177), .B(n_188), .Y(n_350) );
OR2x2_ASAP7_75t_L g371 ( .A(n_177), .B(n_254), .Y(n_371) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_181), .B(n_185), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_185), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_185), .A2(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_SL g494 ( .A(n_185), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_185), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g266 ( .A(n_186), .Y(n_266) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_186), .A2(n_360), .B(n_363), .C(n_365), .Y(n_359) );
AND2x2_ASAP7_75t_L g432 ( .A(n_186), .B(n_207), .Y(n_432) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
INVx1_ASAP7_75t_L g299 ( .A(n_187), .Y(n_299) );
AND2x2_ASAP7_75t_L g369 ( .A(n_187), .B(n_224), .Y(n_369) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx1_ASAP7_75t_L g243 ( .A(n_188), .Y(n_243) );
OR2x2_ASAP7_75t_L g258 ( .A(n_188), .B(n_224), .Y(n_258) );
INVx1_ASAP7_75t_L g274 ( .A(n_188), .Y(n_274) );
AND2x2_ASAP7_75t_L g286 ( .A(n_188), .B(n_195), .Y(n_286) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_188), .Y(n_392) );
NOR2x1_ASAP7_75t_SL g223 ( .A(n_195), .B(n_224), .Y(n_223) );
AO21x1_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_197), .B(n_203), .Y(n_195) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_196), .A2(n_197), .B(n_203), .Y(n_255) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_196), .A2(n_516), .B(n_522), .Y(n_515) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_196), .A2(n_536), .B(n_542), .Y(n_535) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_196), .A2(n_536), .B(n_542), .Y(n_555) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_196), .A2(n_516), .B(n_522), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
INVxp67_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_209), .Y(n_205) );
OR2x2_ASAP7_75t_L g356 ( .A(n_206), .B(n_291), .Y(n_356) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_207), .B(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g438 ( .A(n_207), .B(n_335), .Y(n_438) );
INVx3_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g283 ( .A(n_208), .B(n_264), .Y(n_283) );
AND2x2_ASAP7_75t_L g379 ( .A(n_208), .B(n_292), .Y(n_379) );
INVx1_ASAP7_75t_L g296 ( .A(n_209), .Y(n_296) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
INVx1_ASAP7_75t_L g346 ( .A(n_210), .Y(n_346) );
INVx2_ASAP7_75t_L g313 ( .A(n_211), .Y(n_313) );
HB1xp67_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g263 ( .A(n_212), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g293 ( .A(n_212), .Y(n_293) );
INVx1_ASAP7_75t_L g418 ( .A(n_212), .Y(n_418) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_213), .Y(n_375) );
AOI21x1_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_221), .Y(n_213) );
AO21x2_ASAP7_75t_L g504 ( .A1(n_214), .A2(n_505), .B(n_511), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_216), .B(n_220), .Y(n_215) );
OR2x2_ASAP7_75t_L g389 ( .A(n_222), .B(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_SL g244 ( .A(n_224), .Y(n_244) );
OR2x2_ASAP7_75t_L g267 ( .A(n_224), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g278 ( .A(n_224), .B(n_254), .Y(n_278) );
AND2x2_ASAP7_75t_L g352 ( .A(n_224), .B(n_268), .Y(n_352) );
BUFx2_ASAP7_75t_L g435 ( .A(n_224), .Y(n_435) );
OR2x6_ASAP7_75t_L g224 ( .A(n_225), .B(n_232), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_240), .B(n_245), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
AND2x2_ASAP7_75t_L g387 ( .A(n_236), .B(n_309), .Y(n_387) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g246 ( .A(n_237), .B(n_239), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_238), .B(n_308), .Y(n_409) );
INVx1_ASAP7_75t_L g439 ( .A(n_238), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g335 ( .A(n_239), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_239), .B(n_375), .Y(n_412) );
INVxp67_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
AND2x4_ASAP7_75t_SL g276 ( .A(n_242), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_242), .B(n_270), .Y(n_423) );
INVx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_243), .B(n_325), .Y(n_381) );
AND2x2_ASAP7_75t_L g399 ( .A(n_243), .B(n_352), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_244), .B(n_286), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_244), .A2(n_290), .B(n_332), .C(n_337), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_244), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g426 ( .A1(n_246), .A2(n_319), .B1(n_427), .B2(n_433), .C(n_437), .Y(n_426) );
INVx1_ASAP7_75t_SL g414 ( .A(n_247), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_259), .B1(n_265), .B2(n_269), .C(n_793), .Y(n_248) );
INVx2_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g324 ( .A(n_253), .Y(n_324) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g298 ( .A(n_254), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g329 ( .A(n_254), .B(n_274), .Y(n_329) );
INVx2_ASAP7_75t_L g362 ( .A(n_254), .Y(n_362) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI32xp33_ASAP7_75t_L g413 ( .A1(n_257), .A2(n_304), .A3(n_335), .B1(n_414), .B2(n_415), .Y(n_413) );
OR2x2_ASAP7_75t_L g384 ( .A(n_258), .B(n_371), .Y(n_384) );
INVx1_ASAP7_75t_L g394 ( .A(n_259), .Y(n_394) );
OR2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
INVx2_ASAP7_75t_L g309 ( .A(n_260), .Y(n_309) );
AND2x2_ASAP7_75t_L g380 ( .A(n_260), .B(n_355), .Y(n_380) );
OR2x2_ASAP7_75t_L g411 ( .A(n_260), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_261), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g305 ( .A(n_264), .Y(n_305) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx2_ASAP7_75t_SL g270 ( .A(n_267), .Y(n_270) );
OR2x2_ASAP7_75t_L g357 ( .A(n_267), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_268), .B(n_286), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_268), .B(n_392), .Y(n_391) );
BUFx2_ASAP7_75t_L g404 ( .A(n_268), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_271), .B(n_276), .C(n_279), .Y(n_269) );
AND2x2_ASAP7_75t_L g419 ( .A(n_271), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
BUFx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g345 ( .A(n_275), .B(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_275), .B(n_279), .Y(n_366) );
AND2x2_ASAP7_75t_L g397 ( .A(n_275), .B(n_398), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g407 ( .A1(n_277), .A2(n_408), .B(n_410), .C(n_413), .Y(n_407) );
AOI222xp33_ASAP7_75t_L g281 ( .A1(n_278), .A2(n_282), .B1(n_284), .B2(n_287), .C1(n_295), .C2(n_297), .Y(n_281) );
AND2x2_ASAP7_75t_L g349 ( .A(n_278), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g282 ( .A(n_279), .B(n_283), .Y(n_282) );
INVx2_ASAP7_75t_SL g303 ( .A(n_279), .Y(n_303) );
NAND4xp25_ASAP7_75t_L g280 ( .A(n_281), .B(n_300), .C(n_321), .D(n_331), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_283), .B(n_289), .Y(n_343) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g351 ( .A(n_286), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g358 ( .A(n_286), .Y(n_358) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g321 ( .A1(n_288), .A2(n_322), .B(n_326), .C(n_330), .Y(n_321) );
INVx2_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_289), .B(n_304), .Y(n_425) );
OR2x2_ASAP7_75t_L g429 ( .A(n_289), .B(n_315), .Y(n_429) );
INVx1_ASAP7_75t_L g402 ( .A(n_290), .Y(n_402) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_SL g336 ( .A(n_293), .Y(n_336) );
INVx1_ASAP7_75t_L g316 ( .A(n_294), .Y(n_316) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_296), .B(n_333), .Y(n_332) );
BUFx2_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
AOI322xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .A3(n_304), .B1(n_306), .B2(n_310), .C1(n_311), .C2(n_317), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_SL g382 ( .A1(n_303), .A2(n_383), .B(n_384), .C(n_385), .Y(n_382) );
INVx1_ASAP7_75t_L g405 ( .A(n_304), .Y(n_405) );
NOR2xp67_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g363 ( .A(n_309), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_314), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_315), .Y(n_385) );
INVx2_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx3_ASAP7_75t_L g328 ( .A(n_325), .Y(n_328) );
OR2x2_ASAP7_75t_L g396 ( .A(n_325), .B(n_358), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_325), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx1_ASAP7_75t_SL g428 ( .A(n_329), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_330), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND3xp33_ASAP7_75t_SL g433 ( .A(n_338), .B(n_434), .C(n_436), .Y(n_433) );
NOR3xp33_ASAP7_75t_SL g339 ( .A(n_340), .B(n_377), .C(n_406), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_341), .B(n_359), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_344), .B(n_347), .C(n_353), .Y(n_341) );
OAI31xp33_ASAP7_75t_L g386 ( .A1(n_342), .A2(n_364), .A3(n_387), .B(n_388), .Y(n_386) );
INVx1_ASAP7_75t_SL g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx2_ASAP7_75t_L g401 ( .A(n_349), .Y(n_401) );
INVx1_ASAP7_75t_L g376 ( .A(n_351), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_356), .B(n_357), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g442 ( .A(n_362), .Y(n_442) );
OAI22xp33_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_367), .B1(n_372), .B2(n_376), .Y(n_365) );
INVx3_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_371), .Y(n_383) );
OR2x2_ASAP7_75t_L g434 ( .A(n_371), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
NAND3xp33_ASAP7_75t_SL g377 ( .A(n_378), .B(n_386), .C(n_393), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_380), .B(n_381), .C(n_382), .Y(n_378) );
INVx2_ASAP7_75t_L g415 ( .A(n_379), .Y(n_415) );
INVx1_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_397), .B2(n_399), .C(n_400), .Y(n_393) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_403), .B2(n_405), .Y(n_400) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_416), .C(n_426), .Y(n_406) );
INVxp33_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_419), .B1(n_422), .B2(n_424), .Y(n_416) );
INVx2_ASAP7_75t_L g430 ( .A(n_417), .Y(n_430) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI22xp33_ASAP7_75t_SL g437 ( .A1(n_436), .A2(n_438), .B1(n_439), .B2(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g791 ( .A(n_445), .Y(n_791) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx2_ASAP7_75t_L g455 ( .A(n_446), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
OR2x6_ASAP7_75t_SL g467 ( .A(n_447), .B(n_448), .Y(n_467) );
AND2x6_ASAP7_75t_SL g766 ( .A(n_447), .B(n_449), .Y(n_766) );
OR2x2_ASAP7_75t_L g780 ( .A(n_447), .B(n_449), .Y(n_780) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g782 ( .A(n_455), .B(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_SL g457 ( .A(n_458), .B(n_460), .Y(n_457) );
INVx2_ASAP7_75t_L g785 ( .A(n_458), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_458), .A2(n_788), .B(n_791), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g784 ( .A(n_460), .B(n_785), .Y(n_784) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_767), .B(n_772), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx4f_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OAI22x1_ASAP7_75t_L g773 ( .A1(n_465), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_466), .Y(n_465) );
CKINVDCx11_ASAP7_75t_R g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g774 ( .A(n_468), .Y(n_774) );
AND2x4_ASAP7_75t_L g468 ( .A(n_469), .B(n_684), .Y(n_468) );
NOR3xp33_ASAP7_75t_SL g469 ( .A(n_470), .B(n_596), .C(n_636), .Y(n_469) );
OAI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_512), .B1(n_560), .B2(n_575), .C(n_578), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_481), .Y(n_472) );
INVx2_ASAP7_75t_L g593 ( .A(n_473), .Y(n_593) );
AND2x2_ASAP7_75t_L g623 ( .A(n_473), .B(n_624), .Y(n_623) );
BUFx3_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g561 ( .A(n_474), .B(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g568 ( .A(n_474), .B(n_503), .Y(n_568) );
INVx2_ASAP7_75t_L g574 ( .A(n_474), .Y(n_574) );
AND2x2_ASAP7_75t_L g583 ( .A(n_474), .B(n_483), .Y(n_583) );
INVx1_ASAP7_75t_L g599 ( .A(n_474), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_474), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_SL g481 ( .A(n_482), .B(n_491), .Y(n_481) );
INVx4_ASAP7_75t_L g564 ( .A(n_482), .Y(n_564) );
AND2x2_ASAP7_75t_L g595 ( .A(n_482), .B(n_504), .Y(n_595) );
AND2x2_ASAP7_75t_L g671 ( .A(n_482), .B(n_645), .Y(n_671) );
NAND2x1p5_ASAP7_75t_L g713 ( .A(n_482), .B(n_503), .Y(n_713) );
INVx5_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_483), .B(n_503), .Y(n_600) );
AND2x2_ASAP7_75t_L g624 ( .A(n_483), .B(n_504), .Y(n_624) );
BUFx2_ASAP7_75t_L g640 ( .A(n_483), .Y(n_640) );
NOR2x1_ASAP7_75t_SL g743 ( .A(n_483), .B(n_645), .Y(n_743) );
OR2x6_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g620 ( .A(n_491), .Y(n_620) );
AOI221xp5_ASAP7_75t_L g686 ( .A1(n_491), .A2(n_687), .B1(n_689), .B2(n_691), .C(n_696), .Y(n_686) );
AND2x2_ASAP7_75t_L g706 ( .A(n_491), .B(n_599), .Y(n_706) );
AND2x4_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
INVx1_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
AO21x2_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_494), .B(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g645 ( .A1(n_494), .A2(n_495), .B(n_501), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_496), .B(n_500), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_503), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g584 ( .A(n_503), .B(n_572), .Y(n_584) );
INVx2_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
AND2x2_ASAP7_75t_L g759 ( .A(n_503), .B(n_574), .Y(n_759) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_504), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .Y(n_505) );
NOR3xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_543), .C(n_558), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_523), .Y(n_513) );
INVx2_ASAP7_75t_L g673 ( .A(n_514), .Y(n_673) );
AND2x2_ASAP7_75t_L g718 ( .A(n_514), .B(n_595), .Y(n_718) );
BUFx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g663 ( .A(n_515), .Y(n_663) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_515), .B(n_590), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_517), .B(n_521), .Y(n_516) );
INVx2_ASAP7_75t_L g632 ( .A(n_523), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_523), .B(n_662), .Y(n_688) );
AND2x4_ASAP7_75t_L g721 ( .A(n_523), .B(n_668), .Y(n_721) );
AND2x4_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
AND2x2_ASAP7_75t_L g559 ( .A(n_524), .B(n_554), .Y(n_559) );
OR2x2_ASAP7_75t_L g589 ( .A(n_524), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_SL g658 ( .A(n_524), .B(n_610), .Y(n_658) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
BUFx2_ASAP7_75t_L g603 ( .A(n_525), .Y(n_603) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g577 ( .A(n_526), .Y(n_577) );
OAI21x1_ASAP7_75t_SL g526 ( .A1(n_527), .A2(n_529), .B(n_533), .Y(n_526) );
INVx1_ASAP7_75t_L g534 ( .A(n_528), .Y(n_534) );
INVx2_ASAP7_75t_L g590 ( .A(n_535), .Y(n_590) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_537), .B(n_541), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_543), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_553), .Y(n_544) );
AND2x2_ASAP7_75t_L g558 ( .A(n_545), .B(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g631 ( .A(n_545), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g716 ( .A(n_545), .Y(n_716) );
BUFx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_L g576 ( .A(n_546), .B(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g695 ( .A(n_546), .B(n_555), .Y(n_695) );
AND2x2_ASAP7_75t_L g699 ( .A(n_546), .B(n_565), .Y(n_699) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g668 ( .A(n_547), .Y(n_668) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_547), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_553), .B(n_576), .Y(n_652) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_556), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_554), .B(n_577), .Y(n_762) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g566 ( .A(n_555), .B(n_557), .Y(n_566) );
AND2x2_ASAP7_75t_L g648 ( .A(n_555), .B(n_610), .Y(n_648) );
AND2x2_ASAP7_75t_L g667 ( .A(n_555), .B(n_556), .Y(n_667) );
BUFx2_ASAP7_75t_L g588 ( .A(n_556), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_556), .B(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx3_ASAP7_75t_L g565 ( .A(n_557), .Y(n_565) );
INVxp67_ASAP7_75t_L g608 ( .A(n_557), .Y(n_608) );
INVx1_ASAP7_75t_L g581 ( .A(n_559), .Y(n_581) );
AND2x2_ASAP7_75t_L g617 ( .A(n_559), .B(n_588), .Y(n_617) );
NAND2xp33_ASAP7_75t_L g698 ( .A(n_559), .B(n_699), .Y(n_698) );
AND2x2_ASAP7_75t_L g735 ( .A(n_559), .B(n_736), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_563), .B1(n_566), .B2(n_567), .C(n_569), .Y(n_560) );
AND2x2_ASAP7_75t_L g664 ( .A(n_561), .B(n_564), .Y(n_664) );
AND2x2_ASAP7_75t_SL g683 ( .A(n_561), .B(n_624), .Y(n_683) );
AND2x2_ASAP7_75t_L g701 ( .A(n_561), .B(n_626), .Y(n_701) );
AND2x2_ASAP7_75t_L g756 ( .A(n_561), .B(n_595), .Y(n_756) );
INVx1_ASAP7_75t_L g572 ( .A(n_562), .Y(n_572) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_562), .Y(n_628) );
CKINVDCx16_ASAP7_75t_R g708 ( .A(n_563), .Y(n_708) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_564), .B(n_615), .Y(n_690) );
AND2x2_ASAP7_75t_L g657 ( .A(n_565), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g693 ( .A(n_565), .Y(n_693) );
AND2x2_ASAP7_75t_L g602 ( .A(n_566), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_566), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g744 ( .A(n_566), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_566), .B(n_668), .Y(n_754) );
AND2x4_ASAP7_75t_L g670 ( .A(n_567), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
OR2x2_ASAP7_75t_L g741 ( .A(n_568), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_573), .Y(n_570) );
OR2x2_ASAP7_75t_L g612 ( .A(n_573), .B(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g619 ( .A(n_574), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g650 ( .A(n_574), .B(n_624), .Y(n_650) );
AND2x2_ASAP7_75t_L g724 ( .A(n_574), .B(n_645), .Y(n_724) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g672 ( .A(n_576), .B(n_673), .Y(n_672) );
OAI32xp33_ASAP7_75t_L g737 ( .A1(n_576), .A2(n_738), .A3(n_740), .B1(n_741), .B2(n_744), .Y(n_737) );
AND2x4_ASAP7_75t_L g609 ( .A(n_577), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g707 ( .A(n_577), .B(n_610), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B1(n_585), .B2(n_591), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_SL g696 ( .A1(n_580), .A2(n_594), .B(n_697), .C(n_698), .Y(n_696) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g680 ( .A(n_581), .B(n_608), .Y(n_680) );
INVx1_ASAP7_75t_SL g751 ( .A(n_582), .Y(n_751) );
AND2x4_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
AND2x4_ASAP7_75t_L g654 ( .A(n_584), .B(n_593), .Y(n_654) );
AOI221xp5_ASAP7_75t_L g732 ( .A1(n_584), .A2(n_733), .B1(n_734), .B2(n_735), .C(n_737), .Y(n_732) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_587), .B(n_589), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_589), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
OAI22xp33_ASAP7_75t_L g674 ( .A1(n_592), .A2(n_622), .B1(n_675), .B2(n_676), .Y(n_674) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_593), .A2(n_711), .B(n_719), .C(n_732), .Y(n_710) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g630 ( .A(n_595), .B(n_599), .Y(n_630) );
OAI211xp5_ASAP7_75t_SL g596 ( .A1(n_597), .A2(n_601), .B(n_604), .C(n_633), .Y(n_596) );
OR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g627 ( .A(n_599), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g747 ( .A(n_599), .B(n_743), .Y(n_747) );
OAI32xp33_ASAP7_75t_L g704 ( .A1(n_600), .A2(n_705), .A3(n_707), .B1(n_708), .B2(n_709), .Y(n_704) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_SL g694 ( .A(n_603), .B(n_695), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_611), .B1(n_617), .B2(n_618), .C(n_621), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g761 ( .A(n_608), .B(n_762), .Y(n_761) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_609), .B(n_673), .Y(n_675) );
A2O1A1O1Ixp25_ASAP7_75t_L g746 ( .A1(n_609), .A2(n_678), .B(n_694), .C(n_740), .D(n_747), .Y(n_746) );
AOI31xp33_ASAP7_75t_L g748 ( .A1(n_609), .A2(n_630), .A3(n_740), .B(n_747), .Y(n_748) );
AND2x2_ASAP7_75t_L g662 ( .A(n_610), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_SL g750 ( .A(n_612), .B(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g739 ( .A(n_614), .Y(n_739) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g734 ( .A(n_615), .B(n_626), .Y(n_734) );
INVx1_ASAP7_75t_L g649 ( .A(n_617), .Y(n_649) );
AND2x2_ASAP7_75t_L g634 ( .A(n_618), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AOI31xp33_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .A3(n_629), .B(n_631), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_624), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g757 ( .A(n_624), .B(n_703), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g702 ( .A(n_626), .B(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g728 ( .A(n_626), .Y(n_728) );
INVxp67_ASAP7_75t_L g697 ( .A(n_627), .Y(n_697) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g635 ( .A(n_631), .Y(n_635) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_653), .C(n_669), .Y(n_636) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_646), .B1(n_650), .B2(n_651), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g723 ( .A(n_640), .Y(n_723) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_SL g703 ( .A(n_644), .Y(n_703) );
INVxp67_ASAP7_75t_SL g729 ( .A(n_644), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_644), .B(n_713), .Y(n_730) );
NAND2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
INVx1_ASAP7_75t_L g681 ( .A(n_648), .Y(n_681) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B1(n_664), .B2(n_665), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_662), .A2(n_667), .B1(n_701), .B2(n_702), .C(n_704), .Y(n_700) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g740 ( .A(n_667), .Y(n_740) );
AND2x2_ASAP7_75t_L g677 ( .A(n_668), .B(n_678), .Y(n_677) );
O2A1O1Ixp33_ASAP7_75t_SL g725 ( .A1(n_668), .A2(n_726), .B(n_730), .C(n_731), .Y(n_725) );
AOI211xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_672), .B(n_674), .C(n_679), .Y(n_669) );
AND2x2_ASAP7_75t_L g720 ( .A(n_673), .B(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g731 ( .A(n_678), .Y(n_731) );
AOI21xp33_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B(n_682), .Y(n_679) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
NOR3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_710), .C(n_745), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_686), .B(n_700), .Y(n_685) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g709 ( .A(n_694), .Y(n_709) );
INVxp67_ASAP7_75t_L g733 ( .A(n_698), .Y(n_733) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g717 ( .A(n_707), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B1(n_717), .B2(n_718), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
AOI21xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_722), .B(n_725), .Y(n_719) );
AND2x2_ASAP7_75t_L g722 ( .A(n_723), .B(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g758 ( .A(n_743), .B(n_759), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_748), .B1(n_749), .B2(n_752), .C(n_755), .Y(n_745) );
INVxp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI31xp33_ASAP7_75t_SL g755 ( .A1(n_756), .A2(n_757), .A3(n_758), .B(n_760), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx4_ASAP7_75t_SL g763 ( .A(n_764), .Y(n_763) );
CKINVDCx6p67_ASAP7_75t_R g776 ( .A(n_764), .Y(n_776) );
INVx3_ASAP7_75t_SL g764 ( .A(n_765), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_766), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_767), .A2(n_773), .B(n_777), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
BUFx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
BUFx4f_ASAP7_75t_SL g781 ( .A(n_782), .Y(n_781) );
INVxp67_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
CKINVDCx11_ASAP7_75t_R g788 ( .A(n_789), .Y(n_788) );
CKINVDCx8_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
endmodule