module fake_netlist_6_395_n_192 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_192);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_192;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_32;
wire n_85;
wire n_66;
wire n_130;
wire n_78;
wire n_84;
wire n_99;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_108;
wire n_94;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_30),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_10),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g58 ( 
.A(n_55),
.B(n_0),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_1),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_5),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_43),
.B(n_6),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_8),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

OR2x6_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_54),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_47),
.Y(n_77)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_73),
.B(n_32),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_52),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_52),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_51),
.B1(n_53),
.B2(n_35),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_51),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_71),
.B(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_76),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_62),
.A2(n_46),
.B1(n_34),
.B2(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

O2A1O1Ixp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_61),
.B(n_63),
.C(n_72),
.Y(n_95)
);

AOI21x1_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_61),
.B(n_63),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

NAND2x1_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_75),
.Y(n_98)
);

OAI21x1_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_60),
.B(n_72),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_60),
.B(n_70),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_64),
.B(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI21x1_ASAP7_75t_SL g105 ( 
.A1(n_77),
.A2(n_66),
.B(n_67),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_95),
.A2(n_79),
.B(n_80),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_90),
.B(n_91),
.C(n_66),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_93),
.B1(n_86),
.B2(n_78),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_88),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

AOI21x1_ASAP7_75t_SL g113 ( 
.A1(n_95),
.A2(n_80),
.B(n_88),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_111),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_92),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_76),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_91),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_101),
.B(n_107),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_115),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_117),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_123),
.B(n_117),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_111),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_118),
.Y(n_132)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_116),
.C(n_107),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_112),
.Y(n_134)
);

O2A1O1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_114),
.B(n_120),
.C(n_103),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_112),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g137 ( 
.A(n_127),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_133),
.A2(n_105),
.B(n_50),
.C(n_112),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_68),
.B1(n_69),
.B2(n_67),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_127),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_110),
.B1(n_101),
.B2(n_94),
.Y(n_143)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_143),
.Y(n_144)
);

AOI211xp5_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_135),
.B(n_136),
.C(n_126),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g146 ( 
.A1(n_139),
.A2(n_58),
.B1(n_68),
.B2(n_69),
.C(n_142),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_137),
.B(n_110),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_110),
.B1(n_101),
.B2(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_110),
.B1(n_134),
.B2(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_138),
.B(n_134),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_94),
.C(n_104),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_131),
.Y(n_152)
);

NAND4xp25_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_88),
.C(n_74),
.D(n_104),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_147),
.A2(n_8),
.B(n_9),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_152),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_149),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_131),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_145),
.B(n_10),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_153),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g165 ( 
.A(n_162),
.B(n_74),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

OAI221xp5_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_162),
.B1(n_159),
.B2(n_154),
.C(n_158),
.Y(n_169)
);

O2A1O1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_105),
.B(n_74),
.C(n_88),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

AOI221xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_161),
.B1(n_73),
.B2(n_105),
.C(n_82),
.Y(n_172)
);

OAI221xp5_ASAP7_75t_L g173 ( 
.A1(n_163),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.C(n_98),
.Y(n_173)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_165),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_98),
.C1(n_84),
.C2(n_87),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_17),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_19),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_108),
.A3(n_99),
.B1(n_24),
.B2(n_25),
.C1(n_27),
.C2(n_20),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_21),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_167),
.B(n_99),
.Y(n_179)
);

OAI221xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_106),
.B1(n_96),
.B2(n_99),
.C(n_113),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_176),
.Y(n_181)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_166),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_171),
.B(n_96),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_179),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_106),
.B(n_113),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_182),
.A2(n_174),
.B1(n_173),
.B2(n_180),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_106),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_181),
.Y(n_190)
);

OAI222xp33_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_184),
.B1(n_186),
.B2(n_183),
.C1(n_180),
.C2(n_185),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_188),
.B1(n_187),
.B2(n_190),
.Y(n_192)
);


endmodule