module fake_aes_1323_n_46 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_46);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_43;
wire n_40;
wire n_27;
wire n_39;
NAND2xp5_ASAP7_75t_L g11 ( .A(n_2), .B(n_1), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_3), .B(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_3), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_9), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
OAI21xp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_7), .B(n_8), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_17), .Y(n_20) );
NOR2xp33_ASAP7_75t_L g21 ( .A(n_17), .B(n_2), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_14), .B(n_4), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_12), .Y(n_24) );
AND2x4_ASAP7_75t_L g25 ( .A(n_15), .B(n_5), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_22), .A2(n_18), .B1(n_15), .B2(n_13), .Y(n_26) );
OAI221xp5_ASAP7_75t_L g27 ( .A1(n_21), .A2(n_18), .B1(n_13), .B2(n_11), .C(n_12), .Y(n_27) );
NAND2xp33_ASAP7_75t_R g28 ( .A(n_25), .B(n_16), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_20), .B(n_12), .Y(n_29) );
AOI22xp33_ASAP7_75t_L g30 ( .A1(n_27), .A2(n_25), .B1(n_21), .B2(n_19), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_26), .B(n_25), .Y(n_31) );
BUFx3_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_23), .Y(n_33) );
OR2x2_ASAP7_75t_L g34 ( .A(n_32), .B(n_5), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_30), .Y(n_35) );
AOI21xp5_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_30), .B(n_28), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
NAND2xp5_ASAP7_75t_L g38 ( .A(n_33), .B(n_12), .Y(n_38) );
NAND5xp2_ASAP7_75t_L g39 ( .A(n_36), .B(n_35), .C(n_28), .D(n_6), .E(n_12), .Y(n_39) );
AOI211x1_ASAP7_75t_L g40 ( .A1(n_38), .A2(n_12), .B(n_24), .C(n_10), .Y(n_40) );
INVx1_ASAP7_75t_SL g41 ( .A(n_37), .Y(n_41) );
AOI211xp5_ASAP7_75t_L g42 ( .A1(n_39), .A2(n_24), .B(n_41), .C(n_40), .Y(n_42) );
HB1xp67_ASAP7_75t_L g43 ( .A(n_40), .Y(n_43) );
HB1xp67_ASAP7_75t_L g44 ( .A(n_42), .Y(n_44) );
HB1xp67_ASAP7_75t_L g45 ( .A(n_43), .Y(n_45) );
AOI22xp33_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_24), .B1(n_45), .B2(n_39), .Y(n_46) );
endmodule