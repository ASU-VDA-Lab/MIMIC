module real_aes_8858_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g516 ( .A1(n_0), .A2(n_172), .B(n_517), .C(n_520), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_1), .B(n_467), .Y(n_521) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND3xp33_ASAP7_75t_SL g757 ( .A(n_2), .B(n_89), .C(n_750), .Y(n_757) );
INVx1_ASAP7_75t_L g184 ( .A(n_3), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_4), .B(n_144), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_5), .A2(n_440), .B(n_461), .Y(n_460) );
AO21x2_ASAP7_75t_L g469 ( .A1(n_6), .A2(n_164), .B(n_470), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g192 ( .A1(n_7), .A2(n_37), .B1(n_138), .B2(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_8), .B(n_164), .Y(n_173) );
AND2x6_ASAP7_75t_L g156 ( .A(n_9), .B(n_157), .Y(n_156) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_10), .A2(n_156), .B(n_445), .C(n_530), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_11), .B(n_38), .Y(n_111) );
INVx1_ASAP7_75t_L g134 ( .A(n_12), .Y(n_134) );
INVx1_ASAP7_75t_L g177 ( .A(n_13), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_14), .B(n_142), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_15), .B(n_144), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_16), .B(n_130), .Y(n_248) );
AO32x2_ASAP7_75t_L g190 ( .A1(n_17), .A2(n_129), .A3(n_155), .B1(n_164), .B2(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_18), .B(n_138), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_19), .B(n_130), .Y(n_186) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_20), .A2(n_52), .B1(n_138), .B2(n_193), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_21), .A2(n_80), .B1(n_138), .B2(n_142), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_22), .B(n_138), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_23), .A2(n_155), .B(n_445), .C(n_494), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g746 ( .A1(n_24), .A2(n_57), .B1(n_426), .B2(n_747), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_24), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_25), .A2(n_155), .B(n_445), .C(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_26), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_27), .B(n_159), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_28), .A2(n_440), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_29), .B(n_159), .Y(n_207) );
INVx2_ASAP7_75t_L g140 ( .A(n_30), .Y(n_140) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_31), .A2(n_443), .B(n_453), .C(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g137 ( .A(n_32), .B(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_33), .B(n_159), .Y(n_218) );
XNOR2x2_ASAP7_75t_SL g744 ( .A(n_34), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_35), .B(n_214), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_36), .A2(n_84), .B1(n_732), .B2(n_733), .Y(n_731) );
CKINVDCx20_ASAP7_75t_R g732 ( .A(n_36), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_39), .B(n_492), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_40), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_41), .B(n_144), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_42), .B(n_440), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_43), .A2(n_443), .B(n_447), .C(n_453), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_44), .B(n_138), .Y(n_167) );
INVx1_ASAP7_75t_L g518 ( .A(n_45), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_46), .A2(n_90), .B1(n_193), .B2(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g448 ( .A(n_47), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_48), .B(n_138), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_49), .B(n_138), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_50), .B(n_440), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_51), .B(n_150), .Y(n_171) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_53), .A2(n_58), .B1(n_138), .B2(n_142), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_54), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_55), .B(n_138), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_56), .B(n_138), .Y(n_211) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_57), .A2(n_122), .B1(n_426), .B2(n_427), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g426 ( .A(n_57), .Y(n_426) );
INVx1_ASAP7_75t_L g157 ( .A(n_59), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_60), .B(n_440), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_61), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_62), .A2(n_150), .B(n_180), .C(n_464), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_63), .B(n_138), .Y(n_185) );
INVx1_ASAP7_75t_L g133 ( .A(n_64), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_65), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_66), .B(n_144), .Y(n_485) );
AO32x2_ASAP7_75t_L g228 ( .A1(n_67), .A2(n_155), .A3(n_164), .B1(n_229), .B2(n_233), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_68), .B(n_145), .Y(n_531) );
INVx1_ASAP7_75t_L g148 ( .A(n_69), .Y(n_148) );
INVx1_ASAP7_75t_L g202 ( .A(n_70), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g515 ( .A(n_71), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_72), .B(n_450), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_73), .A2(n_445), .B(n_453), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_74), .B(n_142), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_75), .Y(n_462) );
INVx1_ASAP7_75t_L g752 ( .A(n_76), .Y(n_752) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_77), .A2(n_116), .B1(n_731), .B2(n_734), .C1(n_737), .C2(n_738), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_78), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_79), .B(n_449), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_81), .B(n_193), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_82), .Y(n_487) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_83), .B(n_142), .Y(n_206) );
INVx1_ASAP7_75t_L g733 ( .A(n_84), .Y(n_733) );
INVx2_ASAP7_75t_L g131 ( .A(n_85), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_86), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_87), .B(n_154), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_88), .B(n_142), .Y(n_168) );
OR2x2_ASAP7_75t_L g107 ( .A(n_89), .B(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g119 ( .A(n_89), .B(n_109), .Y(n_119) );
INVx2_ASAP7_75t_L g431 ( .A(n_89), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_91), .A2(n_101), .B1(n_142), .B2(n_143), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_92), .B(n_440), .Y(n_481) );
INVx1_ASAP7_75t_L g484 ( .A(n_93), .Y(n_484) );
INVxp67_ASAP7_75t_L g465 ( .A(n_94), .Y(n_465) );
AOI22xp33_ASAP7_75t_SL g102 ( .A1(n_95), .A2(n_103), .B1(n_753), .B2(n_758), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_96), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g506 ( .A(n_97), .Y(n_506) );
INVx1_ASAP7_75t_L g527 ( .A(n_98), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_99), .B(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g455 ( .A(n_100), .B(n_159), .Y(n_455) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_112), .B(n_750), .Y(n_103) );
NOR2xp33_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g749 ( .A(n_107), .Y(n_749) );
NOR2x2_ASAP7_75t_L g740 ( .A(n_108), .B(n_431), .Y(n_740) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g430 ( .A(n_109), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
AND2x2_ASAP7_75t_L g755 ( .A(n_111), .B(n_756), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_115), .B1(n_741), .B2(n_743), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g742 ( .A(n_114), .Y(n_742) );
OAI22x1_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_120), .B1(n_428), .B2(n_432), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g735 ( .A(n_118), .Y(n_735) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_L g734 ( .A1(n_121), .A2(n_433), .B1(n_735), .B2(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g427 ( .A(n_122), .Y(n_427) );
XNOR2xp5_ASAP7_75t_L g745 ( .A(n_122), .B(n_746), .Y(n_745) );
OR3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_354), .C(n_403), .Y(n_122) );
NAND5xp2_ASAP7_75t_L g123 ( .A(n_124), .B(n_269), .C(n_297), .D(n_327), .E(n_341), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_187), .B1(n_219), .B2(n_224), .C(n_235), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_160), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_126), .B(n_221), .Y(n_220) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g249 ( .A(n_127), .Y(n_249) );
AND2x2_ASAP7_75t_L g257 ( .A(n_127), .B(n_163), .Y(n_257) );
AND2x2_ASAP7_75t_L g280 ( .A(n_127), .B(n_162), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_127), .B(n_174), .Y(n_295) );
OR2x2_ASAP7_75t_L g304 ( .A(n_127), .B(n_242), .Y(n_304) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_127), .Y(n_307) );
AND2x2_ASAP7_75t_L g415 ( .A(n_127), .B(n_242), .Y(n_415) );
OA21x2_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_135), .B(n_158), .Y(n_127) );
OA21x2_ASAP7_75t_L g174 ( .A1(n_128), .A2(n_175), .B(n_186), .Y(n_174) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_129), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_131), .B(n_132), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI21xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_147), .B(n_155), .Y(n_135) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_141), .B(n_144), .Y(n_136) );
INVx3_ASAP7_75t_L g201 ( .A(n_138), .Y(n_201) );
HB1xp67_ASAP7_75t_L g508 ( .A(n_138), .Y(n_508) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g193 ( .A(n_139), .Y(n_193) );
BUFx3_ASAP7_75t_L g231 ( .A(n_139), .Y(n_231) );
AND2x6_ASAP7_75t_L g445 ( .A(n_139), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g143 ( .A(n_140), .Y(n_143) );
INVx1_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
INVx2_ASAP7_75t_L g178 ( .A(n_142), .Y(n_178) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_144), .A2(n_167), .B(n_168), .Y(n_166) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
O2A1O1Ixp5_ASAP7_75t_SL g200 ( .A1(n_144), .A2(n_201), .B(n_202), .C(n_203), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_144), .B(n_465), .Y(n_464) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g229 ( .A1(n_145), .A2(n_154), .B1(n_230), .B2(n_232), .Y(n_229) );
INVx3_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_146), .Y(n_154) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
INVx1_ASAP7_75t_L g214 ( .A(n_146), .Y(n_214) );
AND2x2_ASAP7_75t_L g441 ( .A(n_146), .B(n_151), .Y(n_441) );
INVx1_ASAP7_75t_L g446 ( .A(n_146), .Y(n_446) );
O2A1O1Ixp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_152), .C(n_153), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g183 ( .A1(n_149), .A2(n_172), .B(n_184), .C(n_185), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_149), .A2(n_495), .B(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_153), .A2(n_216), .B(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g191 ( .A1(n_154), .A2(n_172), .B1(n_192), .B2(n_194), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_154), .A2(n_172), .B1(n_245), .B2(n_246), .Y(n_244) );
INVx4_ASAP7_75t_L g519 ( .A(n_154), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g268 ( .A(n_155), .B(n_243), .C(n_244), .Y(n_268) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_156), .A2(n_166), .B(n_169), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g175 ( .A1(n_156), .A2(n_176), .B(n_183), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_156), .A2(n_200), .B(n_204), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g209 ( .A1(n_156), .A2(n_210), .B(n_215), .Y(n_209) );
AND2x4_ASAP7_75t_L g440 ( .A(n_156), .B(n_441), .Y(n_440) );
INVx4_ASAP7_75t_SL g454 ( .A(n_156), .Y(n_454) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_156), .B(n_441), .Y(n_528) );
OA21x2_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_199), .B(n_207), .Y(n_198) );
OA21x2_ASAP7_75t_L g208 ( .A1(n_159), .A2(n_209), .B(n_218), .Y(n_208) );
INVx2_ASAP7_75t_L g233 ( .A(n_159), .Y(n_233) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_159), .A2(n_439), .B(n_442), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_159), .A2(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g500 ( .A(n_159), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_160), .B(n_307), .Y(n_363) );
INVx2_ASAP7_75t_SL g160 ( .A(n_161), .Y(n_160) );
OAI311xp33_ASAP7_75t_L g305 ( .A1(n_161), .A2(n_306), .A3(n_307), .B1(n_308), .C1(n_323), .Y(n_305) );
AND2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_174), .Y(n_161) );
AND2x2_ASAP7_75t_L g266 ( .A(n_162), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g273 ( .A(n_162), .Y(n_273) );
AND2x2_ASAP7_75t_L g394 ( .A(n_162), .B(n_223), .Y(n_394) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_163), .B(n_223), .Y(n_222) );
AND2x2_ASAP7_75t_L g250 ( .A(n_163), .B(n_174), .Y(n_250) );
AND2x2_ASAP7_75t_L g302 ( .A(n_163), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g316 ( .A(n_163), .B(n_249), .Y(n_316) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_173), .Y(n_163) );
INVx4_ASAP7_75t_L g243 ( .A(n_164), .Y(n_243) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_164), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_164), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .Y(n_169) );
INVx2_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
AND2x2_ASAP7_75t_L g265 ( .A(n_174), .B(n_249), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .C(n_180), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_178), .A2(n_474), .B(n_475), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_178), .A2(n_531), .B(n_532), .Y(n_530) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_180), .A2(n_506), .B(n_507), .C(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_181), .A2(n_205), .B(n_206), .Y(n_204) );
INVx4_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g450 ( .A(n_182), .Y(n_450) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_195), .Y(n_187) );
OR2x2_ASAP7_75t_L g360 ( .A(n_188), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_188), .B(n_366), .Y(n_377) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_189), .B(n_373), .Y(n_372) );
BUFx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g234 ( .A(n_190), .Y(n_234) );
AND2x2_ASAP7_75t_L g301 ( .A(n_190), .B(n_228), .Y(n_301) );
AND2x2_ASAP7_75t_L g312 ( .A(n_190), .B(n_208), .Y(n_312) );
AND2x2_ASAP7_75t_L g321 ( .A(n_190), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_195), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_195), .B(n_262), .Y(n_306) );
INVx2_ASAP7_75t_SL g195 ( .A(n_196), .Y(n_195) );
OR2x2_ASAP7_75t_L g293 ( .A(n_196), .B(n_252), .Y(n_293) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_208), .Y(n_196) );
INVx2_ASAP7_75t_L g226 ( .A(n_197), .Y(n_226) );
AND2x2_ASAP7_75t_L g320 ( .A(n_197), .B(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g238 ( .A(n_198), .Y(n_238) );
OR2x2_ASAP7_75t_L g337 ( .A(n_198), .B(n_338), .Y(n_337) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_198), .Y(n_400) );
AND2x2_ASAP7_75t_L g239 ( .A(n_208), .B(n_234), .Y(n_239) );
INVx1_ASAP7_75t_L g260 ( .A(n_208), .Y(n_260) );
AND2x2_ASAP7_75t_L g281 ( .A(n_208), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g322 ( .A(n_208), .Y(n_322) );
INVx1_ASAP7_75t_L g338 ( .A(n_208), .Y(n_338) );
HB1xp67_ASAP7_75t_L g413 ( .A(n_208), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_213), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVxp67_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_221), .B(n_326), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g369 ( .A1(n_221), .A2(n_311), .B1(n_360), .B2(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
OAI211xp5_ASAP7_75t_SL g403 ( .A1(n_222), .A2(n_404), .B(n_406), .C(n_424), .Y(n_403) );
INVx2_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
AND2x2_ASAP7_75t_L g314 ( .A(n_223), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g325 ( .A(n_223), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_224), .B(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_227), .Y(n_224) );
AND2x2_ASAP7_75t_L g298 ( .A(n_225), .B(n_262), .Y(n_298) );
BUFx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_L g330 ( .A(n_226), .B(n_321), .Y(n_330) );
AND2x2_ASAP7_75t_L g349 ( .A(n_226), .B(n_263), .Y(n_349) );
AND2x4_ASAP7_75t_L g285 ( .A(n_227), .B(n_259), .Y(n_285) );
AND2x2_ASAP7_75t_L g423 ( .A(n_227), .B(n_399), .Y(n_423) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
INVx1_ASAP7_75t_L g263 ( .A(n_228), .Y(n_263) );
INVx1_ASAP7_75t_L g362 ( .A(n_228), .Y(n_362) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_231), .Y(n_452) );
INVx2_ASAP7_75t_L g520 ( .A(n_231), .Y(n_520) );
INVx1_ASAP7_75t_L g497 ( .A(n_233), .Y(n_497) );
OR2x2_ASAP7_75t_L g253 ( .A(n_234), .B(n_238), .Y(n_253) );
AND2x2_ASAP7_75t_L g262 ( .A(n_234), .B(n_263), .Y(n_262) );
NOR2xp67_ASAP7_75t_L g282 ( .A(n_234), .B(n_283), .Y(n_282) );
OAI221xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_240), .B1(n_251), .B2(n_254), .C(n_258), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_237), .A2(n_259), .B(n_261), .C(n_264), .Y(n_258) );
AND2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx1_ASAP7_75t_L g283 ( .A(n_238), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_238), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_238), .B(n_260), .Y(n_366) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_238), .Y(n_373) );
AND2x2_ASAP7_75t_L g291 ( .A(n_239), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g328 ( .A(n_239), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
INVx2_ASAP7_75t_L g319 ( .A(n_241), .Y(n_319) );
AOI222xp33_ASAP7_75t_L g368 ( .A1(n_241), .A2(n_252), .B1(n_369), .B2(n_371), .C1(n_372), .C2(n_374), .Y(n_368) );
AND2x2_ASAP7_75t_L g425 ( .A(n_241), .B(n_394), .Y(n_425) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_249), .Y(n_241) );
INVx1_ASAP7_75t_L g315 ( .A(n_242), .Y(n_315) );
AO21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_247), .Y(n_242) );
INVx3_ASAP7_75t_L g467 ( .A(n_243), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_243), .B(n_487), .Y(n_486) );
AO21x2_ASAP7_75t_L g502 ( .A1(n_243), .A2(n_503), .B(n_510), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_243), .B(n_511), .Y(n_510) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_243), .A2(n_526), .B(n_533), .Y(n_525) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x4_ASAP7_75t_L g267 ( .A(n_248), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g353 ( .A(n_250), .B(n_287), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_251), .A2(n_365), .B(n_367), .Y(n_364) );
OR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g292 ( .A(n_252), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_252), .B(n_259), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_252), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_SL g254 ( .A(n_255), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx3_ASAP7_75t_L g318 ( .A(n_256), .Y(n_318) );
OR2x2_ASAP7_75t_L g370 ( .A(n_256), .B(n_292), .Y(n_370) );
AND2x2_ASAP7_75t_L g286 ( .A(n_257), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g324 ( .A(n_257), .B(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_257), .B(n_318), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_257), .B(n_314), .Y(n_340) );
AND2x2_ASAP7_75t_L g344 ( .A(n_257), .B(n_326), .Y(n_344) );
INVxp67_ASAP7_75t_L g276 ( .A(n_259), .Y(n_276) );
BUFx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OAI22xp5_ASAP7_75t_L g333 ( .A1(n_261), .A2(n_334), .B1(n_339), .B2(n_340), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_261), .B(n_366), .Y(n_396) );
INVx1_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g382 ( .A(n_262), .B(n_373), .Y(n_382) );
AND2x2_ASAP7_75t_L g411 ( .A(n_262), .B(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g416 ( .A(n_262), .B(n_366), .Y(n_416) );
INVx1_ASAP7_75t_L g329 ( .A(n_263), .Y(n_329) );
BUFx2_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
INVx1_ASAP7_75t_L g420 ( .A(n_264), .Y(n_420) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NAND2x1p5_ASAP7_75t_L g271 ( .A(n_265), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g296 ( .A(n_266), .Y(n_296) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_267), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g279 ( .A(n_267), .B(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g288 ( .A(n_267), .Y(n_288) );
INVx3_ASAP7_75t_L g326 ( .A(n_267), .Y(n_326) );
OR2x2_ASAP7_75t_L g392 ( .A(n_267), .B(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B(n_277), .C(n_289), .Y(n_269) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_270), .A2(n_407), .B1(n_414), .B2(n_416), .C(n_417), .Y(n_406) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_278), .B(n_284), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_280), .B(n_318), .Y(n_332) );
AND2x2_ASAP7_75t_L g374 ( .A(n_280), .B(n_314), .Y(n_374) );
INVx1_ASAP7_75t_SL g387 ( .A(n_281), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_281), .B(n_335), .Y(n_390) );
INVx1_ASAP7_75t_L g408 ( .A(n_282), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_286), .A2(n_376), .B1(n_378), .B2(n_382), .C(n_383), .Y(n_375) );
AND2x2_ASAP7_75t_L g402 ( .A(n_287), .B(n_394), .Y(n_402) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g386 ( .A(n_288), .Y(n_386) );
AOI21xp33_ASAP7_75t_SL g289 ( .A1(n_290), .A2(n_293), .B(n_294), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g357 ( .A(n_292), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g343 ( .A(n_293), .Y(n_343) );
INVx1_ASAP7_75t_L g371 ( .A(n_294), .Y(n_371) );
OR2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B(n_302), .C(n_305), .Y(n_297) );
OAI31xp33_ASAP7_75t_L g424 ( .A1(n_298), .A2(n_336), .A3(n_423), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g398 ( .A(n_301), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g419 ( .A(n_301), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_303), .B(n_318), .Y(n_346) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g421 ( .A(n_304), .B(n_318), .Y(n_421) );
AOI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_313), .B1(n_317), .B2(n_320), .Y(n_308) );
NAND2xp33_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_312), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g348 ( .A(n_312), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g351 ( .A(n_312), .B(n_335), .Y(n_351) );
AND2x2_ASAP7_75t_L g405 ( .A(n_312), .B(n_400), .Y(n_405) );
AND2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_316), .Y(n_313) );
INVx1_ASAP7_75t_L g380 ( .A(n_316), .Y(n_380) );
NOR2xp67_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OAI32xp33_ASAP7_75t_L g383 ( .A1(n_318), .A2(n_352), .A3(n_384), .B1(n_386), .B2(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g358 ( .A(n_321), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_321), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g381 ( .A(n_325), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_331), .C(n_333), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_329), .B(n_366), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g341 ( .A1(n_330), .A2(n_342), .B1(n_343), .B2(n_344), .C(n_345), .Y(n_341) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g342 ( .A(n_340), .Y(n_342) );
OAI22xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND4xp25_ASAP7_75t_SL g407 ( .A(n_350), .B(n_408), .C(n_409), .D(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
NAND4xp25_ASAP7_75t_SL g354 ( .A(n_355), .B(n_368), .C(n_375), .D(n_388), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_359), .B(n_363), .C(n_364), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g385 ( .A(n_361), .Y(n_385) );
INVx2_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
OR2x2_ASAP7_75t_L g418 ( .A(n_373), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_395), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AND2x2_ASAP7_75t_L g414 ( .A(n_394), .B(n_415), .Y(n_414) );
AOI21xp33_ASAP7_75t_SL g395 ( .A1(n_396), .A2(n_397), .B(n_401), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
CKINVDCx16_ASAP7_75t_R g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B1(n_421), .B2(n_422), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g736 ( .A(n_429), .Y(n_736) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx4_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR5x1_ASAP7_75t_L g434 ( .A(n_435), .B(n_604), .C(n_682), .D(n_706), .E(n_723), .Y(n_434) );
OAI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_476), .B(n_522), .C(n_581), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_456), .Y(n_436) );
AND2x2_ASAP7_75t_L g535 ( .A(n_437), .B(n_458), .Y(n_535) );
INVx5_ASAP7_75t_SL g563 ( .A(n_437), .Y(n_563) );
AND2x2_ASAP7_75t_L g599 ( .A(n_437), .B(n_584), .Y(n_599) );
OR2x2_ASAP7_75t_L g638 ( .A(n_437), .B(n_457), .Y(n_638) );
OR2x2_ASAP7_75t_L g669 ( .A(n_437), .B(n_560), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_437), .B(n_573), .Y(n_705) );
AND2x2_ASAP7_75t_L g717 ( .A(n_437), .B(n_560), .Y(n_717) );
OR2x6_ASAP7_75t_L g437 ( .A(n_438), .B(n_455), .Y(n_437) );
BUFx2_ASAP7_75t_L g492 ( .A(n_440), .Y(n_492) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
O2A1O1Ixp33_ASAP7_75t_L g461 ( .A1(n_444), .A2(n_454), .B(n_462), .C(n_463), .Y(n_461) );
O2A1O1Ixp33_ASAP7_75t_SL g514 ( .A1(n_444), .A2(n_454), .B(n_515), .C(n_516), .Y(n_514) );
INVx5_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_451), .C(n_452), .Y(n_447) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_449), .A2(n_452), .B(n_484), .C(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g716 ( .A(n_456), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g579 ( .A(n_457), .B(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_468), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_458), .B(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_458), .Y(n_572) );
INVx3_ASAP7_75t_L g587 ( .A(n_458), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_458), .B(n_468), .Y(n_611) );
OR2x2_ASAP7_75t_L g620 ( .A(n_458), .B(n_563), .Y(n_620) );
AND2x2_ASAP7_75t_L g624 ( .A(n_458), .B(n_584), .Y(n_624) );
AND2x2_ASAP7_75t_L g630 ( .A(n_458), .B(n_631), .Y(n_630) );
INVxp67_ASAP7_75t_L g667 ( .A(n_458), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_458), .B(n_525), .Y(n_681) );
OA21x2_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_466), .Y(n_458) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_467), .A2(n_513), .B(n_521), .Y(n_512) );
OR2x2_ASAP7_75t_L g573 ( .A(n_468), .B(n_525), .Y(n_573) );
AND2x2_ASAP7_75t_L g584 ( .A(n_468), .B(n_560), .Y(n_584) );
AND2x2_ASAP7_75t_L g596 ( .A(n_468), .B(n_587), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g619 ( .A(n_468), .B(n_525), .Y(n_619) );
INVx1_ASAP7_75t_SL g631 ( .A(n_468), .Y(n_631) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x2_ASAP7_75t_L g524 ( .A(n_469), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_469), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_488), .Y(n_477) );
AND2x2_ASAP7_75t_L g544 ( .A(n_478), .B(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_478), .B(n_501), .Y(n_548) );
AND2x2_ASAP7_75t_L g551 ( .A(n_478), .B(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_478), .B(n_554), .Y(n_553) );
OR2x2_ASAP7_75t_L g576 ( .A(n_478), .B(n_567), .Y(n_576) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_478), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_478), .B(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g626 ( .A(n_478), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g672 ( .A(n_478), .B(n_555), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_478), .B(n_578), .Y(n_699) );
INVx5_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
BUFx2_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
AND2x2_ASAP7_75t_L g635 ( .A(n_479), .B(n_567), .Y(n_635) );
AND2x2_ASAP7_75t_L g719 ( .A(n_479), .B(n_587), .Y(n_719) );
OR2x6_ASAP7_75t_L g479 ( .A(n_480), .B(n_486), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_488), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g708 ( .A(n_488), .Y(n_708) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_501), .Y(n_488) );
AND2x2_ASAP7_75t_L g538 ( .A(n_489), .B(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g547 ( .A(n_489), .B(n_545), .Y(n_547) );
INVx5_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
AND2x2_ASAP7_75t_L g578 ( .A(n_489), .B(n_512), .Y(n_578) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_489), .Y(n_615) );
OR2x6_ASAP7_75t_L g489 ( .A(n_490), .B(n_498), .Y(n_489) );
AOI21xp5_ASAP7_75t_SL g490 ( .A1(n_491), .A2(n_493), .B(n_497), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
INVx1_ASAP7_75t_L g656 ( .A(n_501), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_501), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g689 ( .A(n_501), .B(n_555), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_501), .A2(n_612), .B(n_719), .C(n_720), .Y(n_718) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_512), .Y(n_501) );
BUFx2_ASAP7_75t_L g539 ( .A(n_502), .Y(n_539) );
INVx2_ASAP7_75t_L g543 ( .A(n_502), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_509), .Y(n_503) );
INVx2_ASAP7_75t_L g545 ( .A(n_512), .Y(n_545) );
AND2x2_ASAP7_75t_L g552 ( .A(n_512), .B(n_543), .Y(n_552) );
AND2x2_ASAP7_75t_L g643 ( .A(n_512), .B(n_555), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_518), .B(n_519), .Y(n_517) );
AOI211x1_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_536), .B(n_549), .C(n_574), .Y(n_522) );
INVx1_ASAP7_75t_L g640 ( .A(n_523), .Y(n_640) );
AND2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_535), .Y(n_523) );
INVx5_ASAP7_75t_SL g560 ( .A(n_525), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_525), .B(n_630), .Y(n_629) );
AOI311xp33_ASAP7_75t_L g648 ( .A1(n_525), .A2(n_649), .A3(n_651), .B(n_652), .C(n_658), .Y(n_648) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_525), .A2(n_596), .B(n_684), .C(n_687), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
INVxp67_ASAP7_75t_L g603 ( .A(n_535), .Y(n_603) );
NAND4xp25_ASAP7_75t_SL g536 ( .A(n_537), .B(n_540), .C(n_546), .D(n_548), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_537), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g594 ( .A(n_538), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_541), .B(n_547), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_541), .B(n_554), .Y(n_674) );
BUFx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_542), .B(n_555), .Y(n_692) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g567 ( .A(n_543), .Y(n_567) );
INVxp67_ASAP7_75t_L g602 ( .A(n_544), .Y(n_602) );
AND2x4_ASAP7_75t_L g554 ( .A(n_545), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g628 ( .A(n_545), .B(n_567), .Y(n_628) );
INVx1_ASAP7_75t_L g655 ( .A(n_545), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_545), .B(n_642), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_546), .B(n_616), .Y(n_636) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_547), .B(n_569), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_547), .B(n_616), .Y(n_715) );
INVx1_ASAP7_75t_L g726 ( .A(n_548), .Y(n_726) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_553), .B(n_556), .C(n_564), .Y(n_549) );
INVx1_ASAP7_75t_SL g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g568 ( .A(n_552), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g606 ( .A(n_552), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
AND2x2_ASAP7_75t_L g565 ( .A(n_554), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_554), .B(n_616), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_554), .B(n_635), .Y(n_659) );
OR2x2_ASAP7_75t_L g575 ( .A(n_555), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g607 ( .A(n_555), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_555), .B(n_567), .Y(n_622) );
AND2x2_ASAP7_75t_L g679 ( .A(n_555), .B(n_635), .Y(n_679) );
HB1xp67_ASAP7_75t_L g686 ( .A(n_555), .Y(n_686) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_557), .A2(n_569), .B1(n_691), .B2(n_693), .C(n_696), .Y(n_690) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_561), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g580 ( .A(n_560), .B(n_563), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_560), .B(n_630), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_560), .B(n_587), .Y(n_695) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
OR2x2_ASAP7_75t_L g680 ( .A(n_562), .B(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g694 ( .A(n_562), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_563), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g591 ( .A(n_563), .B(n_584), .Y(n_591) );
AND2x2_ASAP7_75t_L g661 ( .A(n_563), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_563), .B(n_610), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_563), .B(n_711), .Y(n_710) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_565), .A2(n_568), .B(n_570), .Y(n_564) );
INVx2_ASAP7_75t_L g597 ( .A(n_565), .Y(n_597) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g617 ( .A(n_567), .Y(n_617) );
OR2x2_ASAP7_75t_L g621 ( .A(n_569), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g724 ( .A(n_569), .B(n_692), .Y(n_724) );
INVx1_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_572), .B(n_573), .Y(n_571) );
AOI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_577), .B(n_579), .Y(n_574) );
INVx1_ASAP7_75t_L g728 ( .A(n_575), .Y(n_728) );
INVx2_ASAP7_75t_SL g642 ( .A(n_576), .Y(n_642) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g723 ( .A1(n_579), .A2(n_660), .B(n_724), .C(n_725), .Y(n_723) );
OAI322xp33_ASAP7_75t_SL g592 ( .A1(n_580), .A2(n_593), .A3(n_596), .B1(n_597), .B2(n_598), .C1(n_600), .C2(n_603), .Y(n_592) );
INVx2_ASAP7_75t_L g612 ( .A(n_580), .Y(n_612) );
AOI221xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_588), .B1(n_589), .B2(n_591), .C(n_592), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OAI22xp33_ASAP7_75t_SL g658 ( .A1(n_583), .A2(n_659), .B1(n_660), .B2(n_663), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_584), .B(n_587), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_584), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g657 ( .A(n_586), .B(n_619), .Y(n_657) );
INVx1_ASAP7_75t_L g647 ( .A(n_587), .Y(n_647) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_591), .A2(n_701), .B(n_703), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g625 ( .A1(n_593), .A2(n_626), .B(n_629), .Y(n_625) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp67_ASAP7_75t_SL g654 ( .A(n_595), .B(n_655), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_595), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_SL g711 ( .A(n_596), .Y(n_711) );
INVx1_ASAP7_75t_SL g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g604 ( .A(n_605), .B(n_632), .C(n_648), .D(n_664), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_608), .B(n_613), .C(n_625), .Y(n_605) );
INVx1_ASAP7_75t_L g697 ( .A(n_606), .Y(n_697) );
AND2x2_ASAP7_75t_L g645 ( .A(n_607), .B(n_628), .Y(n_645) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_612), .B(n_647), .Y(n_646) );
OAI22xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_618), .B1(n_621), .B2(n_623), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_615), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g663 ( .A(n_616), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_616), .A2(n_655), .B(n_678), .C(n_680), .Y(n_677) );
OR2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g662 ( .A(n_619), .Y(n_662) );
INVx1_ASAP7_75t_L g722 ( .A(n_620), .Y(n_722) );
NAND2xp33_ASAP7_75t_SL g712 ( .A(n_621), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g651 ( .A(n_630), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B(n_637), .C(n_639), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_641), .B1(n_644), .B2(n_646), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_642), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_647), .B(n_668), .Y(n_730) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI21xp33_ASAP7_75t_SL g652 ( .A1(n_653), .A2(n_656), .B(n_657), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g660 ( .A(n_661), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_670), .B1(n_673), .B2(n_675), .C(n_677), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVxp67_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_680), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
NAND3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_690), .C(n_700), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
CKINVDCx16_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVxp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
OAI211xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B(n_709), .C(n_718), .Y(n_706) );
INVx1_ASAP7_75t_L g727 ( .A(n_707), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_712), .B1(n_714), .B2(n_716), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g737 ( .A(n_731), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx3_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2x1p5_ASAP7_75t_L g743 ( .A(n_744), .B(n_748), .Y(n_743) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
CKINVDCx12_ASAP7_75t_R g760 ( .A(n_755), .Y(n_760) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
endmodule