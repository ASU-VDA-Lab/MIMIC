module fake_jpeg_10066_n_77 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_77);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_77;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_0),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

INVx6_ASAP7_75t_SL g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_17),
.B(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_16),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_23),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_20),
.B(n_10),
.C(n_17),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_32),
.B(n_34),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_11),
.Y(n_40)
);

OAI22x1_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_24),
.B1(n_19),
.B2(n_21),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_41),
.A2(n_25),
.B1(n_12),
.B2(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_24),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_23),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_23),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_51),
.C(n_32),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_46),
.A2(n_14),
.B1(n_15),
.B2(n_12),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_31),
.C(n_25),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_53),
.C(n_54),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_47),
.A2(n_39),
.B(n_36),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_34),
.C(n_31),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_34),
.C(n_41),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_56),
.B(n_57),
.Y(n_59)
);

AO22x1_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_36),
.B1(n_3),
.B2(n_2),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_52),
.B(n_45),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.C(n_50),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_67),
.C(n_58),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_65),
.B(n_60),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_49),
.C(n_48),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_14),
.C(n_7),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_69),
.A2(n_70),
.B1(n_11),
.B2(n_3),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

NOR2xp67_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_72),
.A2(n_73),
.B(n_7),
.Y(n_74)
);

NAND3xp33_ASAP7_75t_SL g76 ( 
.A(n_74),
.B(n_8),
.C(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);


endmodule