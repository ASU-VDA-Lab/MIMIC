module real_aes_7912_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_725;
wire n_119;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g108 ( .A(n_0), .Y(n_108) );
INVx1_ASAP7_75t_L g513 ( .A(n_1), .Y(n_513) );
INVx1_ASAP7_75t_L g193 ( .A(n_2), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_3), .A2(n_38), .B1(n_155), .B2(n_455), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_4), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g134 ( .A1(n_5), .A2(n_135), .B(n_142), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_6), .B(n_128), .Y(n_504) );
AND2x6_ASAP7_75t_L g140 ( .A(n_7), .B(n_141), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_8), .A2(n_234), .B(n_235), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_9), .B(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g152 ( .A(n_10), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_11), .B(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g133 ( .A(n_12), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_13), .B(n_165), .Y(n_450) );
INVx1_ASAP7_75t_L g240 ( .A(n_14), .Y(n_240) );
INVx1_ASAP7_75t_L g508 ( .A(n_15), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_16), .B(n_129), .Y(n_489) );
AO32x2_ASAP7_75t_L g470 ( .A1(n_17), .A2(n_128), .A3(n_162), .B1(n_471), .B2(n_475), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_18), .B(n_155), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_19), .B(n_181), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_20), .B(n_129), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_21), .A2(n_50), .B1(n_155), .B2(n_455), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g205 ( .A(n_22), .B(n_135), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g483 ( .A1(n_23), .A2(n_76), .B1(n_155), .B2(n_165), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g466 ( .A(n_24), .B(n_155), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_25), .B(n_126), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_26), .A2(n_238), .B(n_239), .C(n_241), .Y(n_237) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_27), .A2(n_74), .B1(n_724), .B2(n_725), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g725 ( .A(n_27), .Y(n_725) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_29), .B(n_158), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_30), .B(n_150), .Y(n_195) );
INVx1_ASAP7_75t_L g171 ( .A(n_31), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_32), .B(n_158), .Y(n_468) );
INVx2_ASAP7_75t_L g138 ( .A(n_33), .Y(n_138) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_34), .B(n_155), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_35), .B(n_158), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g100 ( .A1(n_36), .A2(n_101), .B1(n_113), .B2(n_735), .C(n_741), .Y(n_100) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_36), .A2(n_62), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_36), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_37), .A2(n_140), .B(n_145), .C(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g169 ( .A(n_40), .Y(n_169) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_41), .Y(n_734) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_42), .B(n_150), .Y(n_254) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_43), .B(n_155), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_44), .A2(n_86), .B1(n_212), .B2(n_455), .Y(n_482) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_45), .B(n_155), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_46), .B(n_155), .Y(n_509) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_47), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_48), .B(n_503), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_49), .B(n_135), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_51), .A2(n_60), .B1(n_155), .B2(n_165), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_52), .A2(n_145), .B1(n_165), .B2(n_167), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_53), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_54), .B(n_155), .Y(n_449) );
CKINVDCx16_ASAP7_75t_R g190 ( .A(n_55), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_56), .B(n_155), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g148 ( .A1(n_57), .A2(n_149), .B(n_151), .C(n_154), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_58), .Y(n_258) );
INVx1_ASAP7_75t_L g143 ( .A(n_59), .Y(n_143) );
INVx1_ASAP7_75t_L g141 ( .A(n_61), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_62), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_63), .B(n_155), .Y(n_514) );
INVx1_ASAP7_75t_L g132 ( .A(n_64), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_65), .Y(n_103) );
AO32x2_ASAP7_75t_L g480 ( .A1(n_66), .A2(n_128), .A3(n_220), .B1(n_475), .B2(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g525 ( .A(n_67), .Y(n_525) );
INVx1_ASAP7_75t_L g463 ( .A(n_68), .Y(n_463) );
A2O1A1Ixp33_ASAP7_75t_SL g180 ( .A1(n_69), .A2(n_154), .B(n_181), .C(n_182), .Y(n_180) );
INVxp67_ASAP7_75t_L g183 ( .A(n_70), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_71), .B(n_165), .Y(n_464) );
INVx1_ASAP7_75t_L g112 ( .A(n_72), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_73), .Y(n_175) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_74), .Y(n_724) );
INVx1_ASAP7_75t_L g251 ( .A(n_75), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_77), .A2(n_140), .B(n_145), .C(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_78), .B(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_79), .B(n_165), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_80), .B(n_194), .Y(n_208) );
INVx2_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_82), .B(n_181), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_83), .B(n_165), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_84), .A2(n_140), .B(n_145), .C(n_192), .Y(n_191) );
OR2x2_ASAP7_75t_L g105 ( .A(n_85), .B(n_106), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_85), .B(n_107), .Y(n_118) );
INVx2_ASAP7_75t_L g438 ( .A(n_85), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_87), .A2(n_99), .B1(n_165), .B2(n_166), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_88), .B(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_89), .Y(n_198) );
A2O1A1Ixp33_ASAP7_75t_L g222 ( .A1(n_90), .A2(n_140), .B(n_145), .C(n_223), .Y(n_222) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_91), .Y(n_230) );
INVx1_ASAP7_75t_L g179 ( .A(n_92), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_93), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_94), .B(n_194), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_95), .B(n_165), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_96), .B(n_128), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_97), .B(n_112), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_98), .A2(n_135), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
OA21x2_ASAP7_75t_L g102 ( .A1(n_103), .A2(n_104), .B(n_110), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g738 ( .A(n_103), .B(n_111), .Y(n_738) );
INVx1_ASAP7_75t_L g758 ( .A(n_103), .Y(n_758) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_SL g740 ( .A(n_105), .Y(n_740) );
INVx2_ASAP7_75t_L g749 ( .A(n_105), .Y(n_749) );
INVx1_ASAP7_75t_SL g754 ( .A(n_105), .Y(n_754) );
NOR2x2_ASAP7_75t_L g733 ( .A(n_106), .B(n_438), .Y(n_733) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g437 ( .A(n_107), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
AND2x2_ASAP7_75t_L g756 ( .A(n_110), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
OAI222xp33_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_722), .B1(n_723), .B2(n_726), .C1(n_730), .C2(n_734), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_119), .B1(n_436), .B2(n_439), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g727 ( .A(n_118), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_119), .A2(n_728), .B1(n_744), .B2(n_745), .Y(n_743) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g728 ( .A(n_120), .Y(n_728) );
AND3x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_358), .C(n_403), .Y(n_120) );
NOR4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_281), .C(n_322), .D(n_339), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_185), .B(n_201), .C(n_243), .Y(n_122) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_159), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_124), .B(n_186), .Y(n_185) );
NOR4xp25_ASAP7_75t_L g305 ( .A(n_124), .B(n_299), .C(n_306), .D(n_312), .Y(n_305) );
AND2x2_ASAP7_75t_L g378 ( .A(n_124), .B(n_267), .Y(n_378) );
AND2x2_ASAP7_75t_L g397 ( .A(n_124), .B(n_343), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_124), .B(n_392), .Y(n_406) );
AND2x2_ASAP7_75t_L g419 ( .A(n_124), .B(n_200), .Y(n_419) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_SL g264 ( .A(n_125), .Y(n_264) );
AND2x2_ASAP7_75t_L g271 ( .A(n_125), .B(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g321 ( .A(n_125), .B(n_160), .Y(n_321) );
AND2x2_ASAP7_75t_SL g332 ( .A(n_125), .B(n_267), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_125), .B(n_160), .Y(n_336) );
AND2x2_ASAP7_75t_L g345 ( .A(n_125), .B(n_270), .Y(n_345) );
BUFx2_ASAP7_75t_L g368 ( .A(n_125), .Y(n_368) );
AND2x2_ASAP7_75t_L g372 ( .A(n_125), .B(n_176), .Y(n_372) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_134), .B(n_157), .Y(n_125) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
NOR2xp33_ASAP7_75t_SL g214 ( .A(n_127), .B(n_215), .Y(n_214) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_127), .B(n_475), .C(n_491), .Y(n_490) );
AO21x1_ASAP7_75t_L g528 ( .A1(n_127), .A2(n_491), .B(n_529), .Y(n_528) );
INVx4_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OA21x2_ASAP7_75t_L g176 ( .A1(n_128), .A2(n_177), .B(n_184), .Y(n_176) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_128), .A2(n_496), .B(n_504), .Y(n_495) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g162 ( .A(n_129), .Y(n_162) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_130), .B(n_131), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
BUFx2_ASAP7_75t_L g234 ( .A(n_135), .Y(n_234) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_140), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g173 ( .A(n_136), .B(n_140), .Y(n_173) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_139), .Y(n_136) );
INVx1_ASAP7_75t_L g503 ( .A(n_137), .Y(n_503) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g146 ( .A(n_138), .Y(n_146) );
INVx1_ASAP7_75t_L g166 ( .A(n_138), .Y(n_166) );
INVx1_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
INVx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_139), .Y(n_168) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx4_ASAP7_75t_SL g156 ( .A(n_140), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g447 ( .A1(n_140), .A2(n_448), .B(n_452), .Y(n_447) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_140), .A2(n_462), .B(n_465), .Y(n_461) );
BUFx3_ASAP7_75t_L g475 ( .A(n_140), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_140), .A2(n_497), .B(n_500), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_140), .A2(n_507), .B(n_511), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_144), .B(n_148), .C(n_156), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_144), .A2(n_156), .B(n_179), .C(n_180), .Y(n_178) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_144), .A2(n_156), .B(n_236), .C(n_237), .Y(n_235) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_146), .Y(n_155) );
BUFx3_ASAP7_75t_L g212 ( .A(n_146), .Y(n_212) );
INVx1_ASAP7_75t_L g455 ( .A(n_146), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g452 ( .A1(n_149), .A2(n_453), .B(n_454), .Y(n_452) );
O2A1O1Ixp5_ASAP7_75t_L g524 ( .A1(n_149), .A2(n_512), .B(n_525), .C(n_526), .Y(n_524) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx4_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_150), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
OAI22xp5_ASAP7_75t_SL g481 ( .A1(n_150), .A2(n_153), .B1(n_482), .B2(n_483), .Y(n_481) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_150), .A2(n_473), .B1(n_492), .B2(n_493), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_153), .B(n_183), .Y(n_182) );
INVx5_ASAP7_75t_L g194 ( .A(n_153), .Y(n_194) );
O2A1O1Ixp5_ASAP7_75t_SL g462 ( .A1(n_154), .A2(n_194), .B(n_463), .C(n_464), .Y(n_462) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_155), .Y(n_227) );
OAI22xp33_ASAP7_75t_L g163 ( .A1(n_156), .A2(n_164), .B1(n_172), .B2(n_173), .Y(n_163) );
INVx1_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
INVx2_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
OA21x2_ASAP7_75t_L g232 ( .A1(n_158), .A2(n_233), .B(n_242), .Y(n_232) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_158), .A2(n_447), .B(n_456), .Y(n_446) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_158), .A2(n_461), .B(n_468), .Y(n_460) );
OR2x2_ASAP7_75t_L g159 ( .A(n_160), .B(n_176), .Y(n_159) );
AND2x2_ASAP7_75t_L g200 ( .A(n_160), .B(n_176), .Y(n_200) );
BUFx2_ASAP7_75t_L g274 ( .A(n_160), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_160), .A2(n_307), .B1(n_309), .B2(n_310), .Y(n_306) );
OR2x2_ASAP7_75t_L g328 ( .A(n_160), .B(n_188), .Y(n_328) );
AND2x2_ASAP7_75t_L g392 ( .A(n_160), .B(n_270), .Y(n_392) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
AND2x2_ASAP7_75t_L g260 ( .A(n_161), .B(n_188), .Y(n_260) );
AND2x2_ASAP7_75t_L g267 ( .A(n_161), .B(n_176), .Y(n_267) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_161), .Y(n_309) );
OR2x2_ASAP7_75t_L g344 ( .A(n_161), .B(n_187), .Y(n_344) );
AO21x2_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_174), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_162), .B(n_175), .Y(n_174) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_162), .A2(n_189), .B(n_197), .Y(n_188) );
INVx2_ASAP7_75t_L g213 ( .A(n_162), .Y(n_213) );
INVx2_ASAP7_75t_L g196 ( .A(n_165), .Y(n_196) );
INVx3_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI22xp5_ASAP7_75t_SL g167 ( .A1(n_168), .A2(n_169), .B1(n_170), .B2(n_171), .Y(n_167) );
INVx2_ASAP7_75t_L g170 ( .A(n_168), .Y(n_170) );
INVx4_ASAP7_75t_L g238 ( .A(n_168), .Y(n_238) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_173), .A2(n_190), .B(n_191), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_173), .A2(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g263 ( .A(n_176), .Y(n_263) );
INVx3_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
BUFx2_ASAP7_75t_L g296 ( .A(n_176), .Y(n_296) );
AND2x2_ASAP7_75t_L g329 ( .A(n_176), .B(n_264), .Y(n_329) );
INVx1_ASAP7_75t_L g451 ( .A(n_181), .Y(n_451) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_185), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_414) );
AND2x2_ASAP7_75t_L g186 ( .A(n_187), .B(n_200), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_187), .B(n_272), .Y(n_276) );
INVx1_ASAP7_75t_L g304 ( .A(n_187), .Y(n_304) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g270 ( .A(n_188), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_195), .C(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g473 ( .A(n_194), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_194), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_194), .A2(n_522), .B(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g507 ( .A1(n_196), .A2(n_508), .B(n_509), .C(n_510), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_199), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_199), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
NAND2x1_ASAP7_75t_SL g201 ( .A(n_202), .B(n_216), .Y(n_201) );
AND2x2_ASAP7_75t_L g280 ( .A(n_202), .B(n_231), .Y(n_280) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_202), .Y(n_354) );
AND2x2_ASAP7_75t_L g381 ( .A(n_202), .B(n_301), .Y(n_381) );
AND2x2_ASAP7_75t_L g389 ( .A(n_202), .B(n_351), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_202), .B(n_246), .Y(n_416) );
INVx3_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x2_ASAP7_75t_L g247 ( .A(n_203), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g265 ( .A(n_203), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g286 ( .A(n_203), .Y(n_286) );
INVx1_ASAP7_75t_L g292 ( .A(n_203), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_203), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g325 ( .A(n_203), .B(n_249), .Y(n_325) );
OR2x2_ASAP7_75t_L g363 ( .A(n_203), .B(n_318), .Y(n_363) );
AOI32xp33_ASAP7_75t_L g375 ( .A1(n_203), .A2(n_376), .A3(n_379), .B1(n_380), .B2(n_381), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_203), .B(n_351), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_203), .B(n_311), .Y(n_426) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_214), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g204 ( .A1(n_205), .A2(n_206), .B(n_213), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_209), .B(n_210), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_210), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g241 ( .A(n_212), .Y(n_241) );
INVx1_ASAP7_75t_L g256 ( .A(n_213), .Y(n_256) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_213), .A2(n_506), .B(n_515), .Y(n_505) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_213), .A2(n_520), .B(n_527), .Y(n_519) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g337 ( .A(n_217), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_231), .Y(n_217) );
INVx1_ASAP7_75t_L g299 ( .A(n_218), .Y(n_299) );
AND2x2_ASAP7_75t_L g301 ( .A(n_218), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_218), .B(n_248), .Y(n_318) );
AND2x2_ASAP7_75t_L g351 ( .A(n_218), .B(n_327), .Y(n_351) );
AND2x2_ASAP7_75t_L g388 ( .A(n_218), .B(n_249), .Y(n_388) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g246 ( .A(n_219), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_219), .B(n_248), .Y(n_278) );
AND2x2_ASAP7_75t_L g285 ( .A(n_219), .B(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g326 ( .A(n_219), .B(n_327), .Y(n_326) );
AO21x2_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_229), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_222), .B(n_228), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_227), .Y(n_223) );
INVx2_ASAP7_75t_L g302 ( .A(n_231), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_231), .B(n_248), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_231), .B(n_293), .Y(n_374) );
INVx1_ASAP7_75t_L g396 ( .A(n_231), .Y(n_396) );
INVx1_ASAP7_75t_L g413 ( .A(n_231), .Y(n_413) );
INVx2_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g266 ( .A(n_232), .B(n_248), .Y(n_266) );
AND2x2_ASAP7_75t_L g288 ( .A(n_232), .B(n_249), .Y(n_288) );
INVx1_ASAP7_75t_L g327 ( .A(n_232), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_238), .B(n_240), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_238), .A2(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g510 ( .A(n_238), .Y(n_510) );
AOI221x1_ASAP7_75t_SL g243 ( .A1(n_244), .A2(n_259), .B1(n_265), .B2(n_267), .C(n_268), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_244), .A2(n_332), .B1(n_399), .B2(n_400), .Y(n_398) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
AND2x2_ASAP7_75t_L g290 ( .A(n_245), .B(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g385 ( .A(n_245), .B(n_265), .Y(n_385) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g341 ( .A(n_246), .B(n_266), .Y(n_341) );
INVx1_ASAP7_75t_L g353 ( .A(n_247), .Y(n_353) );
AND2x2_ASAP7_75t_L g364 ( .A(n_247), .B(n_351), .Y(n_364) );
AND2x2_ASAP7_75t_L g431 ( .A(n_247), .B(n_326), .Y(n_431) );
INVx2_ASAP7_75t_L g293 ( .A(n_248), .Y(n_293) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_256), .B(n_257), .Y(n_249) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_260), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g383 ( .A(n_260), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_261), .B(n_344), .Y(n_347) );
INVx3_ASAP7_75t_SL g261 ( .A(n_262), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_262), .A2(n_383), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NOR2xp33_ASAP7_75t_SL g405 ( .A(n_265), .B(n_291), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_266), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g357 ( .A(n_266), .B(n_285), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_266), .B(n_292), .Y(n_434) );
AND2x2_ASAP7_75t_L g303 ( .A(n_267), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g370 ( .A(n_267), .Y(n_370) );
AOI21xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_273), .B(n_277), .Y(n_268) );
NAND2x1_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_270), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g319 ( .A(n_270), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_SL g331 ( .A(n_270), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g376 ( .A(n_270), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g355 ( .A(n_271), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_271), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_271), .B(n_274), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AOI211xp5_ASAP7_75t_L g342 ( .A1(n_274), .A2(n_313), .B(n_343), .C(n_345), .Y(n_342) );
AOI221xp5_ASAP7_75t_L g360 ( .A1(n_274), .A2(n_361), .B1(n_364), .B2(n_365), .C(n_369), .Y(n_360) );
AND2x2_ASAP7_75t_L g356 ( .A(n_275), .B(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g316 ( .A(n_280), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g387 ( .A(n_280), .B(n_388), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B(n_289), .C(n_314), .Y(n_281) );
NAND3xp33_ASAP7_75t_SL g400 ( .A(n_282), .B(n_401), .C(n_402), .Y(n_400) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_287), .Y(n_283) );
OR2x2_ASAP7_75t_L g373 ( .A(n_284), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B1(n_297), .B2(n_303), .C(n_305), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_291), .B(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_291), .B(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_296), .A2(n_353), .B1(n_354), .B2(n_355), .Y(n_352) );
OR2x2_ASAP7_75t_L g433 ( .A(n_296), .B(n_344), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVxp67_ASAP7_75t_L g407 ( .A(n_299), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_301), .B(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g308 ( .A(n_302), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_304), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_304), .B(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_304), .B(n_371), .Y(n_410) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_308), .Y(n_334) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g424 ( .A(n_313), .B(n_344), .Y(n_424) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_SL g402 ( .A(n_319), .Y(n_402) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
OAI322xp33_ASAP7_75t_SL g322 ( .A1(n_323), .A2(n_328), .A3(n_329), .B1(n_330), .B2(n_333), .C1(n_335), .C2(n_337), .Y(n_322) );
OAI322xp33_ASAP7_75t_L g404 ( .A1(n_323), .A2(n_405), .A3(n_406), .B1(n_407), .B2(n_408), .C1(n_409), .C2(n_411), .Y(n_404) );
CKINVDCx16_ASAP7_75t_R g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx4_ASAP7_75t_L g338 ( .A(n_325), .Y(n_338) );
AND2x2_ASAP7_75t_L g399 ( .A(n_325), .B(n_351), .Y(n_399) );
AND2x2_ASAP7_75t_L g412 ( .A(n_325), .B(n_413), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g423 ( .A(n_328), .Y(n_423) );
INVx1_ASAP7_75t_L g401 ( .A(n_329), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
OR2x2_ASAP7_75t_L g335 ( .A(n_331), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_331), .B(n_372), .Y(n_429) );
OR2x2_ASAP7_75t_L g362 ( .A(n_334), .B(n_363), .Y(n_362) );
INVxp33_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
OAI221xp5_ASAP7_75t_SL g339 ( .A1(n_338), .A2(n_340), .B1(n_342), .B2(n_346), .C(n_348), .Y(n_339) );
NOR2xp67_ASAP7_75t_L g395 ( .A(n_338), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g422 ( .A(n_338), .Y(n_422) );
INVx1_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx3_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
AOI322xp5_ASAP7_75t_L g386 ( .A1(n_345), .A2(n_370), .A3(n_387), .B1(n_389), .B2(n_390), .C1(n_393), .C2(n_397), .Y(n_386) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_352), .B1(n_356), .B2(n_357), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_359), .B(n_382), .Y(n_358) );
NAND2xp5_ASAP7_75t_SL g359 ( .A(n_360), .B(n_375), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_363), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
NAND2xp33_ASAP7_75t_SL g380 ( .A(n_366), .B(n_377), .Y(n_380) );
INVx1_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
OAI322xp33_ASAP7_75t_L g420 ( .A1(n_368), .A2(n_421), .A3(n_423), .B1(n_424), .B2(n_425), .C1(n_427), .C2(n_430), .Y(n_420) );
AOI21xp33_ASAP7_75t_SL g369 ( .A1(n_370), .A2(n_371), .B(n_373), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_378), .B(n_426), .Y(n_435) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_384), .B(n_386), .C(n_398), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
NOR4xp25_ASAP7_75t_L g403 ( .A(n_404), .B(n_414), .C(n_420), .D(n_432), .Y(n_403) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g417 ( .A(n_418), .Y(n_417) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
CKINVDCx14_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g432 ( .A1(n_433), .A2(n_434), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx6_ASAP7_75t_L g729 ( .A(n_437), .Y(n_729) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g726 ( .A1(n_440), .A2(n_727), .B1(n_728), .B2(n_729), .Y(n_726) );
OR2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_644), .Y(n_440) );
NAND5xp2_ASAP7_75t_L g441 ( .A(n_442), .B(n_563), .C(n_578), .D(n_604), .E(n_626), .Y(n_441) );
NOR2xp33_ASAP7_75t_SL g442 ( .A(n_443), .B(n_543), .Y(n_442) );
OAI221xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_484), .B1(n_516), .B2(n_532), .C(n_533), .Y(n_443) );
NOR2xp33_ASAP7_75t_SL g444 ( .A(n_445), .B(n_476), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_445), .B(n_593), .Y(n_592) );
INVx1_ASAP7_75t_SL g720 ( .A(n_445), .Y(n_720) );
AND2x2_ASAP7_75t_L g445 ( .A(n_446), .B(n_457), .Y(n_445) );
INVx1_ASAP7_75t_L g560 ( .A(n_446), .Y(n_560) );
AND2x2_ASAP7_75t_L g562 ( .A(n_446), .B(n_470), .Y(n_562) );
AND2x2_ASAP7_75t_L g572 ( .A(n_446), .B(n_469), .Y(n_572) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_446), .Y(n_590) );
INVx1_ASAP7_75t_L g600 ( .A(n_446), .Y(n_600) );
OR2x2_ASAP7_75t_L g638 ( .A(n_446), .B(n_537), .Y(n_638) );
INVx2_ASAP7_75t_L g688 ( .A(n_446), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_446), .B(n_536), .Y(n_705) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B(n_451), .Y(n_448) );
NOR2xp67_ASAP7_75t_L g457 ( .A(n_458), .B(n_469), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_459), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_459), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_SL g620 ( .A(n_459), .B(n_560), .Y(n_620) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_460), .Y(n_478) );
INVx2_ASAP7_75t_L g537 ( .A(n_460), .Y(n_537) );
OR2x2_ASAP7_75t_L g599 ( .A(n_460), .B(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g538 ( .A(n_469), .B(n_480), .Y(n_538) );
AND2x2_ASAP7_75t_L g555 ( .A(n_469), .B(n_535), .Y(n_555) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g479 ( .A(n_470), .B(n_480), .Y(n_479) );
BUFx2_ASAP7_75t_L g558 ( .A(n_470), .Y(n_558) );
AND2x2_ASAP7_75t_L g687 ( .A(n_470), .B(n_688), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_473), .A2(n_501), .B(n_502), .Y(n_500) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_473), .A2(n_512), .B(n_513), .C(n_514), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g520 ( .A1(n_475), .A2(n_521), .B(n_524), .Y(n_520) );
INVx1_ASAP7_75t_L g532 ( .A(n_476), .Y(n_532) );
AND2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_479), .Y(n_476) );
AND2x2_ASAP7_75t_L g650 ( .A(n_477), .B(n_538), .Y(n_650) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AND2x2_ASAP7_75t_L g651 ( .A(n_478), .B(n_562), .Y(n_651) );
O2A1O1Ixp33_ASAP7_75t_L g618 ( .A1(n_479), .A2(n_619), .B(n_621), .C(n_623), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_479), .B(n_619), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_479), .A2(n_549), .B1(n_692), .B2(n_693), .C(n_695), .Y(n_691) );
INVx1_ASAP7_75t_L g535 ( .A(n_480), .Y(n_535) );
INVx1_ASAP7_75t_L g571 ( .A(n_480), .Y(n_571) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_480), .Y(n_580) );
INVx1_ASAP7_75t_SL g484 ( .A(n_485), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .Y(n_485) );
AND2x2_ASAP7_75t_L g597 ( .A(n_486), .B(n_542), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_486), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_487), .B(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g689 ( .A(n_487), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g721 ( .A(n_487), .Y(n_721) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g551 ( .A(n_488), .Y(n_551) );
AND2x2_ASAP7_75t_L g577 ( .A(n_488), .B(n_531), .Y(n_577) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_488), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g593 ( .A(n_488), .B(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g529 ( .A(n_489), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_494), .B(n_633), .Y(n_668) );
INVx1_ASAP7_75t_SL g672 ( .A(n_494), .Y(n_672) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_505), .Y(n_494) );
INVx3_ASAP7_75t_L g531 ( .A(n_495), .Y(n_531) );
AND2x2_ASAP7_75t_L g542 ( .A(n_495), .B(n_519), .Y(n_542) );
AND2x2_ASAP7_75t_L g564 ( .A(n_495), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g609 ( .A(n_495), .B(n_603), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_495), .B(n_541), .Y(n_690) );
INVx2_ASAP7_75t_L g512 ( .A(n_503), .Y(n_512) );
AND2x2_ASAP7_75t_L g530 ( .A(n_505), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g541 ( .A(n_505), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_505), .B(n_519), .Y(n_566) );
AND2x2_ASAP7_75t_L g602 ( .A(n_505), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_530), .Y(n_517) );
INVx1_ASAP7_75t_L g582 ( .A(n_518), .Y(n_582) );
AND2x2_ASAP7_75t_L g624 ( .A(n_518), .B(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_518), .B(n_545), .Y(n_630) );
AOI21xp5_ASAP7_75t_SL g704 ( .A1(n_518), .A2(n_536), .B(n_559), .Y(n_704) );
AND2x2_ASAP7_75t_L g518 ( .A(n_519), .B(n_528), .Y(n_518) );
OR2x2_ASAP7_75t_L g547 ( .A(n_519), .B(n_528), .Y(n_547) );
AND2x2_ASAP7_75t_L g594 ( .A(n_519), .B(n_531), .Y(n_594) );
INVx2_ASAP7_75t_L g603 ( .A(n_519), .Y(n_603) );
INVx1_ASAP7_75t_L g709 ( .A(n_519), .Y(n_709) );
AND2x2_ASAP7_75t_L g633 ( .A(n_528), .B(n_603), .Y(n_633) );
INVx1_ASAP7_75t_L g658 ( .A(n_528), .Y(n_658) );
AND2x2_ASAP7_75t_L g567 ( .A(n_530), .B(n_551), .Y(n_567) );
AND2x2_ASAP7_75t_L g579 ( .A(n_530), .B(n_580), .Y(n_579) );
INVx2_ASAP7_75t_SL g697 ( .A(n_530), .Y(n_697) );
INVx2_ASAP7_75t_L g587 ( .A(n_531), .Y(n_587) );
AND2x2_ASAP7_75t_L g625 ( .A(n_531), .B(n_541), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_531), .B(n_709), .Y(n_708) );
OAI21xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_538), .B(n_539), .Y(n_533) );
AND2x2_ASAP7_75t_L g640 ( .A(n_534), .B(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g694 ( .A(n_534), .Y(n_694) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
INVx1_ASAP7_75t_L g614 ( .A(n_535), .Y(n_614) );
BUFx2_ASAP7_75t_L g713 ( .A(n_535), .Y(n_713) );
BUFx2_ASAP7_75t_L g584 ( .A(n_536), .Y(n_584) );
AND2x2_ASAP7_75t_L g686 ( .A(n_536), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g669 ( .A(n_537), .Y(n_669) );
AND2x4_ASAP7_75t_L g596 ( .A(n_538), .B(n_559), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_538), .B(n_620), .Y(n_632) );
AOI32xp33_ASAP7_75t_L g556 ( .A1(n_539), .A2(n_557), .A3(n_559), .B1(n_561), .B2(n_562), .Y(n_556) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
INVx3_ASAP7_75t_L g545 ( .A(n_540), .Y(n_545) );
OR2x2_ASAP7_75t_L g681 ( .A(n_540), .B(n_637), .Y(n_681) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g550 ( .A(n_541), .B(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g657 ( .A(n_541), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g549 ( .A(n_542), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g561 ( .A(n_542), .B(n_551), .Y(n_561) );
INVx1_ASAP7_75t_L g682 ( .A(n_542), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_542), .B(n_657), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_548), .B(n_552), .C(n_556), .Y(n_543) );
OAI322xp33_ASAP7_75t_L g652 ( .A1(n_544), .A2(n_589), .A3(n_653), .B1(n_655), .B2(n_659), .C1(n_660), .C2(n_664), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_546), .Y(n_544) );
INVxp67_ASAP7_75t_L g617 ( .A(n_545), .Y(n_617) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g671 ( .A(n_547), .B(n_672), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_547), .B(n_587), .Y(n_718) );
INVxp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g610 ( .A(n_550), .Y(n_610) );
OR2x2_ASAP7_75t_L g696 ( .A(n_551), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_554), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g605 ( .A(n_555), .B(n_584), .Y(n_605) );
AND2x2_ASAP7_75t_L g676 ( .A(n_555), .B(n_589), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_555), .B(n_663), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g563 ( .A1(n_557), .A2(n_564), .B1(n_567), .B2(n_568), .C(n_573), .Y(n_563) );
OR2x2_ASAP7_75t_L g574 ( .A(n_557), .B(n_570), .Y(n_574) );
AND2x2_ASAP7_75t_L g662 ( .A(n_557), .B(n_663), .Y(n_662) );
AOI32xp33_ASAP7_75t_L g701 ( .A1(n_557), .A2(n_587), .A3(n_702), .B1(n_703), .B2(n_706), .Y(n_701) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_558), .B(n_594), .C(n_617), .Y(n_635) );
AND2x2_ASAP7_75t_L g661 ( .A(n_558), .B(n_654), .Y(n_661) );
INVxp67_ASAP7_75t_L g641 ( .A(n_559), .Y(n_641) );
BUFx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_562), .B(n_614), .Y(n_670) );
INVx2_ASAP7_75t_L g680 ( .A(n_562), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_562), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g649 ( .A(n_565), .Y(n_649) );
OR2x2_ASAP7_75t_L g575 ( .A(n_566), .B(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_568), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_571), .Y(n_654) );
AND2x2_ASAP7_75t_L g613 ( .A(n_572), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g659 ( .A(n_572), .Y(n_659) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_572), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AOI21xp33_ASAP7_75t_SL g598 ( .A1(n_574), .A2(n_599), .B(n_601), .Y(n_598) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g692 ( .A(n_577), .B(n_602), .Y(n_692) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_581), .B(n_591), .C(n_598), .Y(n_578) );
AND2x2_ASAP7_75t_L g622 ( .A(n_580), .B(n_590), .Y(n_622) );
INVx2_ASAP7_75t_L g637 ( .A(n_580), .Y(n_637) );
OR2x2_ASAP7_75t_L g675 ( .A(n_580), .B(n_638), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_580), .B(n_718), .Y(n_717) );
AOI211xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_583), .B(n_585), .C(n_588), .Y(n_581) );
INVxp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_584), .B(n_622), .Y(n_621) );
OAI211xp5_ASAP7_75t_L g703 ( .A1(n_585), .A2(n_680), .B(n_704), .C(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2x1p5_ASAP7_75t_L g601 ( .A(n_586), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g643 ( .A(n_587), .B(n_633), .Y(n_643) );
INVx1_ASAP7_75t_L g648 ( .A(n_587), .Y(n_648) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVxp33_ASAP7_75t_L g699 ( .A(n_593), .Y(n_699) );
AND2x2_ASAP7_75t_L g678 ( .A(n_594), .B(n_657), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_599), .A2(n_661), .B(n_662), .Y(n_660) );
OAI322xp33_ASAP7_75t_L g679 ( .A1(n_601), .A2(n_680), .A3(n_681), .B1(n_682), .B2(n_683), .C1(n_685), .C2(n_689), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_606), .B1(n_611), .B2(n_615), .C(n_618), .Y(n_604) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g656 ( .A(n_609), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g700 ( .A(n_613), .Y(n_700) );
INVxp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_616), .B(n_636), .Y(n_702) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
INVx1_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g665 ( .A(n_625), .B(n_633), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_631), .B2(n_633), .C(n_634), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g645 ( .A1(n_629), .A2(n_646), .B1(n_650), .B2(n_651), .C(n_652), .Y(n_645) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_633), .B(n_648), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_639), .B2(n_642), .Y(n_634) );
OR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
INVx2_ASAP7_75t_SL g663 ( .A(n_638), .Y(n_663) );
INVxp67_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_645), .B(n_666), .C(n_691), .D(n_701), .E(n_711), .Y(n_644) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_647), .B(n_649), .Y(n_646) );
NOR4xp25_ASAP7_75t_L g719 ( .A(n_648), .B(n_654), .C(n_720), .D(n_721), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_651), .A2(n_712), .B1(n_714), .B2(n_716), .C(n_719), .Y(n_711) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g710 ( .A(n_657), .Y(n_710) );
OAI322xp33_ASAP7_75t_L g667 ( .A1(n_661), .A2(n_668), .A3(n_669), .B1(n_670), .B2(n_671), .C1(n_673), .C2(n_677), .Y(n_667) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_679), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_676), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g712 ( .A(n_687), .B(n_713), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_695) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
BUFx2_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp33_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_750), .B(n_755), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g742 ( .A(n_743), .B(n_748), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
endmodule