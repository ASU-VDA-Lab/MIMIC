module fake_ariane_878_n_100 (n_8, n_24, n_7, n_22, n_43, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_41, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_45, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_100);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_41;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_100;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_53;
wire n_66;
wire n_71;
wire n_96;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_72;
wire n_82;
wire n_57;
wire n_70;
wire n_85;
wire n_94;
wire n_48;
wire n_58;
wire n_65;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_81;
wire n_87;
wire n_55;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_78;
wire n_59;
wire n_63;
wire n_99;
wire n_54;

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_22),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_42),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_R g48 ( 
.A(n_18),
.B(n_6),
.Y(n_48)
);

AO21x2_ASAP7_75t_L g49 ( 
.A1(n_25),
.A2(n_24),
.B(n_14),
.Y(n_49)
);

AO21x2_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_36),
.B(n_33),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_19),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_3),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_R g55 ( 
.A(n_23),
.B(n_13),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_R g58 ( 
.A(n_0),
.B(n_5),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

NOR2x1p5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_31),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_32),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_11),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_2),
.B(n_8),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_66),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_7),
.B(n_9),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_44),
.B1(n_28),
.B2(n_37),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_61),
.B(n_43),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_62),
.B(n_59),
.C(n_69),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_SL g78 ( 
.A(n_46),
.B(n_47),
.C(n_53),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_77),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_80),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

AND2x4_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_60),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_64),
.B1(n_63),
.B2(n_52),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_49),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_86),
.Y(n_94)
);

AOI221xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_87),
.B1(n_88),
.B2(n_91),
.C(n_90),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_93),
.A2(n_72),
.B(n_48),
.C(n_50),
.Y(n_96)
);

CKINVDCx5p33_ASAP7_75t_R g97 ( 
.A(n_95),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_98),
.B1(n_68),
.B2(n_55),
.Y(n_100)
);


endmodule