module fake_jpeg_9901_n_130 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_130);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_122;
wire n_75;
wire n_121;
wire n_99;
wire n_102;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_8),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_69),
.Y(n_87)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx5_ASAP7_75t_SL g73 ( 
.A(n_63),
.Y(n_73)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_66),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_0),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_1),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_69),
.B(n_39),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_79),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_47),
.B1(n_48),
.B2(n_43),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_78),
.B1(n_80),
.B2(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_64),
.A2(n_44),
.B1(n_61),
.B2(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_2),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_54),
.B1(n_52),
.B2(n_56),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_2),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_89),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_69),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_50),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_53),
.B1(n_49),
.B2(n_4),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_5),
.B1(n_9),
.B2(n_10),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_5),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_76),
.A2(n_22),
.B1(n_6),
.B2(n_7),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_96),
.C(n_97),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_99),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_73),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_113),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_112),
.B(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_115),
.B(n_114),
.Y(n_116)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_116),
.A2(n_108),
.B(n_106),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_101),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_21),
.B(n_25),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_26),
.C(n_28),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_125),
.A2(n_102),
.B(n_75),
.Y(n_126)
);

OAI321xp33_ASAP7_75t_L g127 ( 
.A1(n_126),
.A2(n_103),
.A3(n_109),
.B1(n_111),
.B2(n_29),
.C(n_32),
.Y(n_127)
);

OAI31xp33_ASAP7_75t_SL g128 ( 
.A1(n_127),
.A2(n_111),
.A3(n_103),
.B(n_107),
.Y(n_128)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_128),
.A2(n_100),
.B(n_104),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_129),
.Y(n_130)
);


endmodule