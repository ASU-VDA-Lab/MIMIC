module real_aes_6415_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_496;
wire n_281;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_183;
wire n_266;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_1), .A2(n_138), .B(n_143), .C(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g250 ( .A(n_2), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_3), .A2(n_133), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_4), .B(n_210), .Y(n_456) );
AOI21xp33_ASAP7_75t_L g211 ( .A1(n_5), .A2(n_133), .B(n_212), .Y(n_211) );
AND2x6_ASAP7_75t_L g138 ( .A(n_6), .B(n_139), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g131 ( .A1(n_7), .A2(n_132), .B(n_140), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_40), .Y(n_116) );
INVx1_ASAP7_75t_L g545 ( .A(n_9), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g496 ( .A(n_10), .B(n_182), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_11), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g217 ( .A(n_12), .Y(n_217) );
INVx1_ASAP7_75t_L g130 ( .A(n_13), .Y(n_130) );
INVx1_ASAP7_75t_L g150 ( .A(n_14), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g504 ( .A1(n_15), .A2(n_151), .B(n_165), .C(n_505), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_16), .B(n_210), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_17), .B(n_167), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_18), .B(n_133), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_19), .B(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_20), .A2(n_198), .B(n_224), .C(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_21), .B(n_210), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_22), .B(n_182), .Y(n_478) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_23), .A2(n_147), .B(n_149), .C(n_151), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g442 ( .A(n_24), .B(n_182), .Y(n_442) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_25), .Y(n_473) );
INVx1_ASAP7_75t_L g441 ( .A(n_26), .Y(n_441) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_27), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_28), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_29), .B(n_182), .Y(n_251) );
INVx1_ASAP7_75t_L g466 ( .A(n_30), .Y(n_466) );
INVx1_ASAP7_75t_L g229 ( .A(n_31), .Y(n_229) );
INVx2_ASAP7_75t_L g136 ( .A(n_32), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_33), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_34), .A2(n_198), .B(n_218), .C(n_454), .Y(n_453) );
INVxp67_ASAP7_75t_L g467 ( .A(n_35), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_36), .A2(n_138), .B(n_143), .C(n_162), .Y(n_161) );
A2O1A1Ixp33_ASAP7_75t_L g439 ( .A1(n_37), .A2(n_143), .B(n_440), .C(n_445), .Y(n_439) );
CKINVDCx14_ASAP7_75t_R g452 ( .A(n_38), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_39), .A2(n_68), .B1(n_695), .B2(n_696), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_39), .Y(n_695) );
INVx1_ASAP7_75t_L g227 ( .A(n_41), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g543 ( .A1(n_42), .A2(n_169), .B(n_215), .C(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_43), .B(n_182), .Y(n_181) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_44), .A2(n_85), .B1(n_714), .B2(n_715), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_44), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_45), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_46), .Y(n_463) );
INVx1_ASAP7_75t_L g511 ( .A(n_47), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g230 ( .A(n_48), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_49), .B(n_133), .Y(n_201) );
OAI22xp5_ASAP7_75t_SL g693 ( .A1(n_50), .A2(n_694), .B1(n_697), .B2(n_698), .Y(n_693) );
INVx1_ASAP7_75t_L g698 ( .A(n_50), .Y(n_698) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_51), .A2(n_143), .B1(n_224), .B2(n_226), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_52), .Y(n_173) );
CKINVDCx16_ASAP7_75t_R g247 ( .A(n_53), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_54), .A2(n_215), .B(n_216), .C(n_218), .Y(n_214) );
CKINVDCx14_ASAP7_75t_R g542 ( .A(n_55), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_56), .Y(n_186) );
INVx1_ASAP7_75t_L g213 ( .A(n_57), .Y(n_213) );
INVx1_ASAP7_75t_L g139 ( .A(n_58), .Y(n_139) );
INVx1_ASAP7_75t_L g129 ( .A(n_59), .Y(n_129) );
INVx1_ASAP7_75t_SL g455 ( .A(n_60), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_61), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_62), .B(n_210), .Y(n_515) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_63), .Y(n_110) );
INVx1_ASAP7_75t_L g476 ( .A(n_64), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_SL g237 ( .A1(n_65), .A2(n_167), .B(n_218), .C(n_238), .Y(n_237) );
INVxp67_ASAP7_75t_L g239 ( .A(n_66), .Y(n_239) );
AOI22xp33_ASAP7_75t_SL g103 ( .A1(n_67), .A2(n_104), .B1(n_720), .B2(n_727), .Y(n_103) );
INVx1_ASAP7_75t_L g696 ( .A(n_68), .Y(n_696) );
INVx1_ASAP7_75t_L g725 ( .A(n_69), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_70), .A2(n_133), .B(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_71), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_72), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_73), .A2(n_133), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g177 ( .A(n_74), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_75), .A2(n_132), .B(n_462), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g438 ( .A(n_76), .Y(n_438) );
INVx1_ASAP7_75t_L g503 ( .A(n_77), .Y(n_503) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_78), .A2(n_138), .B(n_143), .C(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_79), .A2(n_133), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g506 ( .A(n_80), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_81), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g127 ( .A(n_82), .Y(n_127) );
INVx1_ASAP7_75t_L g495 ( .A(n_83), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_84), .B(n_167), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_85), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_86), .A2(n_138), .B(n_143), .C(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g112 ( .A(n_87), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g428 ( .A(n_87), .Y(n_428) );
OR2x2_ASAP7_75t_L g692 ( .A(n_87), .B(n_114), .Y(n_692) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_88), .A2(n_143), .B(n_475), .C(n_479), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g117 ( .A1(n_89), .A2(n_118), .B1(n_693), .B2(n_699), .C1(n_706), .C2(n_707), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_90), .B(n_126), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g254 ( .A(n_91), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g194 ( .A1(n_92), .A2(n_138), .B(n_143), .C(n_195), .Y(n_194) );
CKINVDCx20_ASAP7_75t_R g203 ( .A(n_93), .Y(n_203) );
OAI22xp33_ASAP7_75t_SL g711 ( .A1(n_94), .A2(n_712), .B1(n_716), .B2(n_717), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_94), .Y(n_716) );
INVx1_ASAP7_75t_L g236 ( .A(n_95), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_96), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_97), .B(n_164), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_98), .B(n_155), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_99), .B(n_155), .Y(n_154) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_100), .A2(n_133), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g514 ( .A(n_101), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_102), .B(n_725), .Y(n_724) );
AOI22x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_108), .B1(n_117), .B2(n_710), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_109), .A2(n_711), .B(n_718), .Y(n_710) );
NOR2xp33_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
BUFx2_ASAP7_75t_L g719 ( .A(n_112), .Y(n_719) );
NOR2x2_ASAP7_75t_L g709 ( .A(n_113), .B(n_428), .Y(n_709) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g427 ( .A(n_114), .B(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_427), .B1(n_429), .B2(n_692), .Y(n_118) );
INVx2_ASAP7_75t_SL g700 ( .A(n_119), .Y(n_700) );
OR4x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_323), .C(n_382), .D(n_409), .Y(n_119) );
NAND3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_265), .C(n_290), .Y(n_120) );
O2A1O1Ixp33_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_188), .B(n_208), .C(n_241), .Y(n_121) );
AOI211xp5_ASAP7_75t_SL g413 ( .A1(n_122), .A2(n_414), .B(n_416), .C(n_419), .Y(n_413) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_157), .Y(n_122) );
INVx1_ASAP7_75t_L g288 ( .A(n_123), .Y(n_288) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OR2x2_ASAP7_75t_L g263 ( .A(n_124), .B(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g295 ( .A(n_124), .Y(n_295) );
AND2x2_ASAP7_75t_L g350 ( .A(n_124), .B(n_319), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_124), .B(n_206), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_124), .B(n_207), .Y(n_408) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g269 ( .A(n_125), .Y(n_269) );
AND2x2_ASAP7_75t_L g312 ( .A(n_125), .B(n_175), .Y(n_312) );
AND2x2_ASAP7_75t_L g330 ( .A(n_125), .B(n_207), .Y(n_330) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_131), .B(n_154), .Y(n_125) );
INVx1_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
INVx2_ASAP7_75t_L g192 ( .A(n_126), .Y(n_192) );
O2A1O1Ixp33_ASAP7_75t_L g437 ( .A1(n_126), .A2(n_178), .B(n_438), .C(n_439), .Y(n_437) );
OA21x2_ASAP7_75t_L g539 ( .A1(n_126), .A2(n_540), .B(n_546), .Y(n_539) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x2_ASAP7_75t_L g156 ( .A(n_127), .B(n_128), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_130), .Y(n_128) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_138), .Y(n_133) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_134), .B(n_138), .Y(n_178) );
AND2x2_ASAP7_75t_L g134 ( .A(n_135), .B(n_137), .Y(n_134) );
INVx1_ASAP7_75t_L g444 ( .A(n_135), .Y(n_444) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
INVx1_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
INVx1_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_137), .Y(n_148) );
INVx3_ASAP7_75t_L g165 ( .A(n_137), .Y(n_165) );
INVx1_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
INVx4_ASAP7_75t_SL g153 ( .A(n_138), .Y(n_153) );
BUFx3_ASAP7_75t_L g445 ( .A(n_138), .Y(n_445) );
O2A1O1Ixp33_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_142), .B(n_146), .C(n_153), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_142), .A2(n_153), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_142), .A2(n_153), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g451 ( .A1(n_142), .A2(n_153), .B(n_452), .C(n_453), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_142), .A2(n_153), .B(n_463), .C(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_SL g502 ( .A1(n_142), .A2(n_153), .B(n_503), .C(n_504), .Y(n_502) );
O2A1O1Ixp33_ASAP7_75t_SL g510 ( .A1(n_142), .A2(n_153), .B(n_511), .C(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_SL g541 ( .A1(n_142), .A2(n_153), .B(n_542), .C(n_543), .Y(n_541) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_145), .Y(n_143) );
BUFx3_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_144), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_147), .B(n_150), .Y(n_149) );
OAI22xp33_ASAP7_75t_L g465 ( .A1(n_147), .A2(n_164), .B1(n_466), .B2(n_467), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_147), .B(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_147), .B(n_514), .Y(n_513) );
INVx4_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g226 ( .A1(n_148), .A2(n_227), .B1(n_228), .B2(n_229), .Y(n_226) );
INVx2_ASAP7_75t_L g228 ( .A(n_148), .Y(n_228) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
OAI22xp33_ASAP7_75t_L g222 ( .A1(n_153), .A2(n_178), .B1(n_223), .B2(n_230), .Y(n_222) );
INVx1_ASAP7_75t_L g479 ( .A(n_153), .Y(n_479) );
INVx4_ASAP7_75t_L g174 ( .A(n_155), .Y(n_174) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_155), .A2(n_234), .B(n_240), .Y(n_233) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_155), .Y(n_449) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g171 ( .A(n_156), .Y(n_171) );
INVx4_ASAP7_75t_L g262 ( .A(n_157), .Y(n_262) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_157), .A2(n_318), .B(n_320), .Y(n_317) );
AND2x2_ASAP7_75t_L g398 ( .A(n_157), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_175), .Y(n_157) );
INVx1_ASAP7_75t_L g205 ( .A(n_158), .Y(n_205) );
AND2x2_ASAP7_75t_L g267 ( .A(n_158), .B(n_207), .Y(n_267) );
OR2x2_ASAP7_75t_L g296 ( .A(n_158), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g310 ( .A(n_158), .Y(n_310) );
INVx3_ASAP7_75t_L g319 ( .A(n_158), .Y(n_319) );
AND2x2_ASAP7_75t_L g329 ( .A(n_158), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g362 ( .A(n_158), .B(n_268), .Y(n_362) );
AND2x2_ASAP7_75t_L g386 ( .A(n_158), .B(n_342), .Y(n_386) );
OR2x6_ASAP7_75t_L g158 ( .A(n_159), .B(n_172), .Y(n_158) );
AOI21xp5_ASAP7_75t_SL g159 ( .A1(n_160), .A2(n_161), .B(n_170), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_166), .B(n_168), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_164), .A2(n_250), .B(n_251), .C(n_252), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_164), .A2(n_441), .B(n_442), .C(n_443), .Y(n_440) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_165), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_165), .B(n_239), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_165), .B(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g180 ( .A1(n_168), .A2(n_181), .B(n_183), .Y(n_180) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_168), .A2(n_476), .B(n_477), .C(n_478), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g494 ( .A1(n_168), .A2(n_477), .B(n_495), .C(n_496), .Y(n_494) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_171), .A2(n_222), .B(n_231), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_171), .B(n_232), .Y(n_231) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_171), .A2(n_246), .B(n_253), .Y(n_245) );
NOR2xp33_ASAP7_75t_SL g172 ( .A(n_173), .B(n_174), .Y(n_172) );
INVx3_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_174), .B(n_447), .Y(n_446) );
AO21x2_ASAP7_75t_L g471 ( .A1(n_174), .A2(n_472), .B(n_480), .Y(n_471) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_174), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g207 ( .A(n_175), .Y(n_207) );
AND2x2_ASAP7_75t_L g422 ( .A(n_175), .B(n_264), .Y(n_422) );
AO21x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_184), .B(n_185), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B(n_179), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g246 ( .A1(n_178), .A2(n_247), .B(n_248), .Y(n_246) );
OAI21xp5_ASAP7_75t_L g472 ( .A1(n_178), .A2(n_473), .B(n_474), .Y(n_472) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_178), .A2(n_492), .B(n_493), .Y(n_491) );
INVx4_ASAP7_75t_L g198 ( .A(n_182), .Y(n_198) );
INVx2_ASAP7_75t_L g215 ( .A(n_182), .Y(n_215) );
INVx1_ASAP7_75t_L g460 ( .A(n_184), .Y(n_460) );
AO21x2_ASAP7_75t_L g484 ( .A1(n_184), .A2(n_485), .B(n_486), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_187), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_187), .B(n_254), .Y(n_253) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_187), .A2(n_491), .B(n_497), .Y(n_490) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_204), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_190), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g342 ( .A(n_190), .B(n_330), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_190), .B(n_319), .Y(n_404) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx2_ASAP7_75t_L g264 ( .A(n_191), .Y(n_264) );
AND2x2_ASAP7_75t_L g268 ( .A(n_191), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g309 ( .A(n_191), .B(n_310), .Y(n_309) );
AO21x2_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_193), .B(n_202), .Y(n_191) );
INVx1_ASAP7_75t_L g469 ( .A(n_192), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_192), .B(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_201), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g454 ( .A(n_198), .B(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g218 ( .A(n_200), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_204), .B(n_305), .Y(n_327) );
INVx1_ASAP7_75t_L g366 ( .A(n_204), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_204), .B(n_293), .Y(n_410) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_206), .Y(n_204) );
AND2x2_ASAP7_75t_L g273 ( .A(n_205), .B(n_268), .Y(n_273) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_207), .B(n_264), .Y(n_297) );
INVx1_ASAP7_75t_L g376 ( .A(n_207), .Y(n_376) );
AOI322xp5_ASAP7_75t_L g400 ( .A1(n_208), .A2(n_315), .A3(n_375), .B1(n_401), .B2(n_403), .C1(n_405), .C2(n_407), .Y(n_400) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_209), .B(n_220), .Y(n_208) );
AND2x2_ASAP7_75t_L g255 ( .A(n_209), .B(n_233), .Y(n_255) );
INVx1_ASAP7_75t_SL g258 ( .A(n_209), .Y(n_258) );
AND2x2_ASAP7_75t_L g260 ( .A(n_209), .B(n_221), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_209), .B(n_277), .Y(n_283) );
INVx2_ASAP7_75t_L g302 ( .A(n_209), .Y(n_302) );
AND2x2_ASAP7_75t_L g315 ( .A(n_209), .B(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g353 ( .A(n_209), .B(n_277), .Y(n_353) );
BUFx2_ASAP7_75t_L g370 ( .A(n_209), .Y(n_370) );
AND2x2_ASAP7_75t_L g384 ( .A(n_209), .B(n_244), .Y(n_384) );
OA21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_219), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_220), .B(n_272), .Y(n_299) );
AND2x2_ASAP7_75t_L g426 ( .A(n_220), .B(n_302), .Y(n_426) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_233), .Y(n_220) );
OR2x2_ASAP7_75t_L g271 ( .A(n_221), .B(n_272), .Y(n_271) );
INVx3_ASAP7_75t_L g277 ( .A(n_221), .Y(n_277) );
AND2x2_ASAP7_75t_L g322 ( .A(n_221), .B(n_245), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_221), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_221), .Y(n_406) );
INVx2_ASAP7_75t_L g252 ( .A(n_224), .Y(n_252) );
INVx3_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g477 ( .A(n_228), .Y(n_477) );
AND2x2_ASAP7_75t_L g257 ( .A(n_233), .B(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
BUFx2_ASAP7_75t_L g285 ( .A(n_233), .Y(n_285) );
AND2x2_ASAP7_75t_L g304 ( .A(n_233), .B(n_277), .Y(n_304) );
INVx3_ASAP7_75t_L g316 ( .A(n_233), .Y(n_316) );
OR2x2_ASAP7_75t_L g326 ( .A(n_233), .B(n_277), .Y(n_326) );
AOI31xp33_ASAP7_75t_SL g241 ( .A1(n_242), .A2(n_256), .A3(n_259), .B(n_261), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_255), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_243), .B(n_278), .Y(n_289) );
OR2x2_ASAP7_75t_L g313 ( .A(n_243), .B(n_283), .Y(n_313) );
INVx1_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_244), .B(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g334 ( .A(n_244), .B(n_326), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g344 ( .A(n_244), .B(n_316), .Y(n_344) );
AND2x2_ASAP7_75t_L g351 ( .A(n_244), .B(n_352), .Y(n_351) );
NAND2x1_ASAP7_75t_L g379 ( .A(n_244), .B(n_315), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_244), .B(n_370), .Y(n_380) );
AND2x2_ASAP7_75t_L g392 ( .A(n_244), .B(n_277), .Y(n_392) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g272 ( .A(n_245), .Y(n_272) );
INVx1_ASAP7_75t_L g338 ( .A(n_255), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_255), .B(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_257), .B(n_333), .Y(n_367) );
AND2x4_ASAP7_75t_L g278 ( .A(n_258), .B(n_279), .Y(n_278) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_263), .Y(n_261) );
INVx2_ASAP7_75t_L g357 ( .A(n_263), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g374 ( .A(n_263), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g305 ( .A(n_264), .B(n_295), .Y(n_305) );
AND2x2_ASAP7_75t_L g399 ( .A(n_264), .B(n_269), .Y(n_399) );
INVx1_ASAP7_75t_L g424 ( .A(n_264), .Y(n_424) );
AOI221xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_270), .B1(n_273), .B2(n_274), .C(n_280), .Y(n_265) );
CKINVDCx14_ASAP7_75t_R g286 ( .A(n_266), .Y(n_286) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_267), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_270), .B(n_321), .Y(n_340) );
INVx3_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
OR2x2_ASAP7_75t_L g389 ( .A(n_271), .B(n_285), .Y(n_389) );
AND2x2_ASAP7_75t_L g303 ( .A(n_272), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g333 ( .A(n_272), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_272), .B(n_316), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g403 ( .A(n_272), .B(n_373), .C(n_404), .Y(n_403) );
AOI211xp5_ASAP7_75t_SL g336 ( .A1(n_273), .A2(n_337), .B(n_339), .C(n_347), .Y(n_336) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_275), .A2(n_326), .B1(n_327), .B2(n_328), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_276), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_276), .B(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g418 ( .A(n_278), .B(n_392), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_286), .B1(n_287), .B2(n_289), .Y(n_280) );
NOR2xp33_ASAP7_75t_SL g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_284), .B(n_333), .Y(n_364) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_287), .A2(n_379), .B1(n_410), .B2(n_417), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_298), .B1(n_300), .B2(n_305), .C(n_306), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_296), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_296), .A2(n_307), .B1(n_313), .B2(n_314), .C(n_317), .Y(n_306) );
INVx1_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_SL g321 ( .A(n_302), .Y(n_321) );
OR2x2_ASAP7_75t_L g394 ( .A(n_302), .B(n_326), .Y(n_394) );
AND2x2_ASAP7_75t_L g396 ( .A(n_302), .B(n_304), .Y(n_396) );
INVx1_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
AOI21xp33_ASAP7_75t_SL g365 ( .A1(n_308), .A2(n_366), .B(n_367), .Y(n_365) );
OR2x2_ASAP7_75t_L g372 ( .A(n_308), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g346 ( .A(n_309), .B(n_330), .Y(n_346) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp33_ASAP7_75t_SL g363 ( .A(n_314), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_315), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_316), .B(n_352), .Y(n_415) );
O2A1O1Ixp33_ASAP7_75t_L g331 ( .A1(n_319), .A2(n_332), .B(n_334), .C(n_335), .Y(n_331) );
NAND2x1_ASAP7_75t_SL g356 ( .A(n_319), .B(n_357), .Y(n_356) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_320), .A2(n_369), .B1(n_371), .B2(n_374), .Y(n_368) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_322), .B(n_412), .Y(n_411) );
NAND5xp2_ASAP7_75t_L g323 ( .A(n_324), .B(n_336), .C(n_354), .D(n_368), .E(n_377), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_325), .B(n_331), .Y(n_324) );
INVx1_ASAP7_75t_L g381 ( .A(n_327), .Y(n_381) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_329), .A2(n_348), .B1(n_388), .B2(n_390), .C(n_393), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_330), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_333), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_333), .B(n_399), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_343), .B2(n_345), .Y(n_339) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_351), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g421 ( .A(n_350), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_362), .B2(n_363), .C(n_365), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g412 ( .A(n_370), .Y(n_412) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OAI21xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_380), .B(n_381), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_387), .C(n_400), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_385), .A2(n_410), .B(n_411), .C(n_413), .Y(n_409) );
INVx1_ASAP7_75t_SL g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_389), .B(n_391), .Y(n_390) );
AOI21xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_397), .Y(n_393) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g702 ( .A(n_427), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_429), .Y(n_703) );
XOR2xp5_ASAP7_75t_L g712 ( .A(n_429), .B(n_713), .Y(n_712) );
OR3x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_603), .C(n_650), .Y(n_429) );
NAND3xp33_ASAP7_75t_SL g430 ( .A(n_431), .B(n_549), .C(n_574), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_489), .B1(n_516), .B2(n_519), .C(n_527), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_457), .B(n_482), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_434), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_434), .B(n_532), .Y(n_647) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_448), .Y(n_434) );
AND2x2_ASAP7_75t_L g518 ( .A(n_435), .B(n_488), .Y(n_518) );
AND2x2_ASAP7_75t_L g567 ( .A(n_435), .B(n_487), .Y(n_567) );
AND2x2_ASAP7_75t_L g588 ( .A(n_435), .B(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g593 ( .A(n_435), .B(n_560), .Y(n_593) );
OR2x2_ASAP7_75t_L g601 ( .A(n_435), .B(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g673 ( .A(n_435), .B(n_470), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_435), .B(n_622), .Y(n_687) );
INVx3_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g533 ( .A(n_436), .B(n_448), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_436), .B(n_470), .Y(n_534) );
AND2x4_ASAP7_75t_L g555 ( .A(n_436), .B(n_488), .Y(n_555) );
AND2x2_ASAP7_75t_L g585 ( .A(n_436), .B(n_459), .Y(n_585) );
AND2x2_ASAP7_75t_L g594 ( .A(n_436), .B(n_584), .Y(n_594) );
AND2x2_ASAP7_75t_L g610 ( .A(n_436), .B(n_471), .Y(n_610) );
OR2x2_ASAP7_75t_L g619 ( .A(n_436), .B(n_602), .Y(n_619) );
AND2x2_ASAP7_75t_L g625 ( .A(n_436), .B(n_560), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_436), .B(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g639 ( .A(n_436), .B(n_484), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_436), .B(n_529), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_436), .B(n_589), .Y(n_678) );
OR2x6_ASAP7_75t_L g436 ( .A(n_437), .B(n_446), .Y(n_436) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_444), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
AND2x2_ASAP7_75t_L g584 ( .A(n_448), .B(n_470), .Y(n_584) );
AND2x2_ASAP7_75t_L g589 ( .A(n_448), .B(n_471), .Y(n_589) );
INVx1_ASAP7_75t_L g645 ( .A(n_448), .Y(n_645) );
OA21x2_ASAP7_75t_L g448 ( .A1(n_449), .A2(n_450), .B(n_456), .Y(n_448) );
OA21x2_ASAP7_75t_L g500 ( .A1(n_449), .A2(n_501), .B(n_507), .Y(n_500) );
OA21x2_ASAP7_75t_L g508 ( .A1(n_449), .A2(n_509), .B(n_515), .Y(n_508) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
AND2x2_ASAP7_75t_L g554 ( .A(n_458), .B(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_470), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_459), .B(n_518), .Y(n_517) );
BUFx3_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
OR2x2_ASAP7_75t_L g602 ( .A(n_459), .B(n_470), .Y(n_602) );
OR2x2_ASAP7_75t_L g663 ( .A(n_459), .B(n_570), .Y(n_663) );
OA21x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B(n_468), .Y(n_459) );
INVx1_ASAP7_75t_L g485 ( .A(n_461), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_468), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_470), .B(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g622 ( .A(n_470), .B(n_484), .Y(n_622) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g561 ( .A(n_471), .Y(n_561) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_483), .A2(n_667), .B1(n_671), .B2(n_674), .C(n_675), .Y(n_666) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_SL g530 ( .A(n_484), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_484), .B(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g661 ( .A(n_484), .B(n_518), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_487), .B(n_532), .Y(n_653) );
AND2x2_ASAP7_75t_L g560 ( .A(n_488), .B(n_561), .Y(n_560) );
INVx1_ASAP7_75t_SL g564 ( .A(n_489), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_489), .B(n_570), .Y(n_600) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
AND2x2_ASAP7_75t_L g526 ( .A(n_490), .B(n_500), .Y(n_526) );
INVx4_ASAP7_75t_L g538 ( .A(n_490), .Y(n_538) );
BUFx3_ASAP7_75t_L g580 ( .A(n_490), .Y(n_580) );
AND3x2_ASAP7_75t_L g595 ( .A(n_490), .B(n_596), .C(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g677 ( .A(n_499), .B(n_591), .Y(n_677) );
AND2x2_ASAP7_75t_L g685 ( .A(n_499), .B(n_570), .Y(n_685) );
INVx1_ASAP7_75t_SL g690 ( .A(n_499), .Y(n_690) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_508), .Y(n_499) );
INVx1_ASAP7_75t_SL g548 ( .A(n_500), .Y(n_548) );
AND2x2_ASAP7_75t_L g571 ( .A(n_500), .B(n_538), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_500), .B(n_522), .Y(n_573) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
OR2x2_ASAP7_75t_L g618 ( .A(n_500), .B(n_538), .Y(n_618) );
INVx2_ASAP7_75t_L g524 ( .A(n_508), .Y(n_524) );
AND2x2_ASAP7_75t_L g558 ( .A(n_508), .B(n_539), .Y(n_558) );
OR2x2_ASAP7_75t_L g578 ( .A(n_508), .B(n_539), .Y(n_578) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_508), .Y(n_598) );
INVx1_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
AOI21xp33_ASAP7_75t_L g648 ( .A1(n_517), .A2(n_557), .B(n_649), .Y(n_648) );
AOI322xp5_ASAP7_75t_L g684 ( .A1(n_519), .A2(n_529), .A3(n_555), .B1(n_685), .B2(n_686), .C1(n_688), .C2(n_691), .Y(n_684) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_521), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g521 ( .A(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_522), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_L g547 ( .A(n_523), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x2_ASAP7_75t_L g615 ( .A(n_524), .B(n_538), .Y(n_615) );
AND2x2_ASAP7_75t_L g682 ( .A(n_524), .B(n_539), .Y(n_682) );
INVx1_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g623 ( .A(n_526), .B(n_577), .Y(n_623) );
AOI31xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_531), .A3(n_534), .B(n_535), .Y(n_527) );
AND2x2_ASAP7_75t_L g582 ( .A(n_529), .B(n_560), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_529), .B(n_552), .Y(n_664) );
AND2x2_ASAP7_75t_L g683 ( .A(n_529), .B(n_588), .Y(n_683) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_533), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_532), .B(n_560), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_532), .B(n_589), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g609 ( .A(n_532), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_532), .B(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_533), .B(n_589), .Y(n_621) );
INVx1_ASAP7_75t_L g665 ( .A(n_533), .Y(n_665) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_547), .Y(n_536) );
INVxp67_ASAP7_75t_L g617 ( .A(n_537), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_538), .B(n_548), .Y(n_553) );
INVx1_ASAP7_75t_L g659 ( .A(n_538), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_538), .B(n_636), .Y(n_670) );
BUFx3_ASAP7_75t_L g570 ( .A(n_539), .Y(n_570) );
AND2x2_ASAP7_75t_L g596 ( .A(n_539), .B(n_548), .Y(n_596) );
INVx2_ASAP7_75t_L g636 ( .A(n_539), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g668 ( .A(n_547), .B(n_669), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B(n_556), .C(n_565), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI21xp33_ASAP7_75t_L g599 ( .A1(n_551), .A2(n_600), .B(n_601), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_552), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_552), .B(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x2_ASAP7_75t_L g632 ( .A(n_553), .B(n_578), .Y(n_632) );
INVx3_ASAP7_75t_L g563 ( .A(n_555), .Y(n_563) );
OAI22xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_559), .B1(n_562), .B2(n_564), .Y(n_556) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_558), .A2(n_582), .B(n_583), .Y(n_581) );
AND2x2_ASAP7_75t_L g607 ( .A(n_558), .B(n_571), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_558), .B(n_659), .Y(n_658) );
INVxp67_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
OR2x2_ASAP7_75t_L g562 ( .A(n_561), .B(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g631 ( .A(n_561), .Y(n_631) );
OAI21xp5_ASAP7_75t_SL g575 ( .A1(n_562), .A2(n_576), .B(n_581), .Y(n_575) );
OAI22xp33_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_568), .B1(n_572), .B2(n_573), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_567), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g591 ( .A(n_570), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_570), .B(n_613), .Y(n_612) );
NOR3xp33_ASAP7_75t_L g574 ( .A(n_575), .B(n_586), .C(n_599), .Y(n_574) );
OAI22xp5_ASAP7_75t_SL g641 ( .A1(n_576), .A2(n_642), .B1(n_646), .B2(n_647), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_577), .B(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
OR2x2_ASAP7_75t_L g646 ( .A(n_578), .B(n_579), .Y(n_646) );
AND2x2_ASAP7_75t_L g654 ( .A(n_579), .B(n_635), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
O2A1O1Ixp33_ASAP7_75t_SL g662 ( .A1(n_580), .A2(n_663), .B(n_664), .C(n_665), .Y(n_662) );
OR2x2_ASAP7_75t_L g689 ( .A(n_580), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
OAI21xp33_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_590), .B(n_592), .Y(n_586) );
INVx1_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_588), .A2(n_625), .B(n_626), .C(n_629), .Y(n_624) );
OAI21xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_594), .B(n_595), .Y(n_592) );
AND2x2_ASAP7_75t_L g657 ( .A(n_596), .B(n_615), .Y(n_657) );
INVxp67_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g635 ( .A(n_598), .B(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g640 ( .A(n_600), .Y(n_640) );
NAND3xp33_ASAP7_75t_SL g603 ( .A(n_604), .B(n_624), .C(n_637), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B(n_608), .C(n_616), .Y(n_604) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g674 ( .A(n_611), .Y(n_674) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .Y(n_611) );
INVx1_ASAP7_75t_L g634 ( .A(n_613), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_613), .B(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
A2O1A1Ixp33_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_618), .B(n_619), .C(n_620), .Y(n_616) );
INVx2_ASAP7_75t_SL g628 ( .A(n_618), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_619), .A2(n_630), .B1(n_632), .B2(n_633), .Y(n_629) );
OAI21xp33_ASAP7_75t_SL g620 ( .A1(n_621), .A2(n_622), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
AOI211xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B(n_641), .C(n_648), .Y(n_637) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVxp33_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g691 ( .A(n_645), .Y(n_691) );
NAND4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_666), .C(n_679), .D(n_684), .Y(n_650) );
AOI211xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_655), .C(n_662), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B(n_660), .Y(n_655) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_656), .A2(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g688 ( .A(n_663), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_683), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g705 ( .A(n_692), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_693), .Y(n_706) );
INVx1_ASAP7_75t_L g697 ( .A(n_694), .Y(n_697) );
OAI22xp5_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_701), .B1(n_703), .B2(n_704), .Y(n_699) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx3_ASAP7_75t_SL g726 ( .A(n_709), .Y(n_726) );
INVx1_ASAP7_75t_L g717 ( .A(n_712), .Y(n_717) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
CKINVDCx12_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g728 ( .A(n_723), .Y(n_728) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
endmodule