module fake_jpeg_18283_n_162 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_162);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_162;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx8_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_3),
.B(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_12),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_11),
.B(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_45),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_29),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_85),
.Y(n_95)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_56),
.B(n_0),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_71),
.Y(n_90)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_86),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_85),
.A2(n_58),
.B1(n_49),
.B2(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_87),
.A2(n_93),
.B1(n_94),
.B2(n_57),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_66),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_54),
.B1(n_51),
.B2(n_48),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_75),
.B1(n_48),
.B2(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_100),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_91),
.A2(n_74),
.B1(n_64),
.B2(n_81),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_82),
.B1(n_57),
.B2(n_61),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_107),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_92),
.A2(n_67),
.B1(n_55),
.B2(n_73),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_89),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_108),
.A2(n_73),
.B1(n_61),
.B2(n_6),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_102),
.B(n_66),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_112),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_60),
.A3(n_70),
.B1(n_62),
.B2(n_65),
.Y(n_112)
);

BUFx24_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_120),
.Y(n_135)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_126),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_124),
.A2(n_0),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_125),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_69),
.B(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_127),
.B(n_131),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_115),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_136),
.B1(n_139),
.B2(n_116),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_53),
.B(n_7),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_133),
.B(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_137),
.Y(n_144)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_138),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_53),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_146),
.B1(n_147),
.B2(n_133),
.Y(n_150)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_111),
.B1(n_126),
.B2(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_9),
.B1(n_10),
.B2(n_14),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_132),
.B1(n_128),
.B2(n_140),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_149),
.A2(n_150),
.B1(n_147),
.B2(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_127),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_152),
.A2(n_148),
.B1(n_141),
.B2(n_143),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_141),
.C(n_24),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_22),
.C(n_25),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_30),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_31),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_32),
.B(n_33),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_43),
.B(n_35),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_34),
.B(n_36),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_37),
.Y(n_162)
);


endmodule