module fake_jpeg_27709_n_221 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_221);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_221;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_1),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_30),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_20),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_50),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g51 ( 
.A(n_43),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_33),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_58),
.B(n_62),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_25),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_30),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_41),
.A2(n_23),
.B1(n_29),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_60),
.B1(n_53),
.B2(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_76),
.B1(n_85),
.B2(n_2),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_68),
.B(n_49),
.Y(n_97)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_51),
.A2(n_42),
.B1(n_34),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_70),
.A2(n_75),
.B1(n_86),
.B2(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_32),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_37),
.C(n_44),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_77),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_58),
.A2(n_24),
.B1(n_44),
.B2(n_16),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_37),
.C(n_44),
.Y(n_77)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_81),
.B(n_83),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_24),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_3),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_24),
.B1(n_17),
.B2(n_16),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_19),
.B1(n_31),
.B2(n_36),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_48),
.A2(n_39),
.B1(n_17),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_61),
.B1(n_56),
.B2(n_52),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_62),
.B(n_46),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_92),
.A2(n_105),
.B(n_102),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_101),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_107),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_88),
.B(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_108),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_56),
.B1(n_61),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_90),
.B1(n_71),
.B2(n_66),
.Y(n_128)
);

NOR2x1_ASAP7_75t_SL g119 ( 
.A(n_102),
.B(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_104),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_1),
.B(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_2),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_110),
.B(n_114),
.Y(n_127)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_112),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_81),
.B(n_13),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_113),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_65),
.B(n_12),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_119),
.A2(n_123),
.B(n_130),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_109),
.B(n_82),
.C(n_83),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_124),
.C(n_103),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_91),
.B(n_80),
.C(n_78),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_78),
.C(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_128),
.Y(n_142)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_133),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_66),
.B1(n_84),
.B2(n_69),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_132),
.A2(n_111),
.B1(n_104),
.B2(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_108),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_3),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_105),
.Y(n_144)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_136),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_3),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_138),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_140),
.B(n_147),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_137),
.B(n_126),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_159),
.B(n_136),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_154),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_106),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_149),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_92),
.C(n_97),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_117),
.B(n_114),
.Y(n_150)
);

AOI221xp5_ASAP7_75t_L g164 ( 
.A1(n_150),
.A2(n_127),
.B1(n_131),
.B2(n_120),
.C(n_137),
.Y(n_164)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_111),
.C(n_96),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_121),
.C(n_134),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_120),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_152),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_157),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_125),
.Y(n_156)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_99),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_123),
.A2(n_4),
.B(n_5),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_170),
.B(n_153),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_135),
.B(n_137),
.C(n_122),
.D(n_133),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_157),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_141),
.B(n_159),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_127),
.C(n_7),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_173),
.C(n_146),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_6),
.C(n_7),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_143),
.Y(n_175)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

OA21x2_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_6),
.B(n_8),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_176),
.A2(n_146),
.B1(n_153),
.B2(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_160),
.C(n_161),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_184),
.B1(n_187),
.B2(n_188),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_179),
.B(n_182),
.Y(n_194)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_150),
.CI(n_155),
.CON(n_183),
.SN(n_183)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_186),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_168),
.A2(n_158),
.B1(n_156),
.B2(n_142),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_142),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_185),
.B(n_172),
.C(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_156),
.B1(n_148),
.B2(n_10),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_191),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_192),
.C(n_195),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_180),
.C(n_177),
.Y(n_195)
);

OAI21x1_ASAP7_75t_SL g196 ( 
.A1(n_183),
.A2(n_163),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_194),
.B(n_182),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_201),
.B(n_202),
.Y(n_207)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_193),
.B(n_171),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_180),
.C(n_178),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_174),
.C(n_167),
.Y(n_210)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_191),
.B(n_183),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_170),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_206),
.B(n_210),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_204),
.A2(n_174),
.B1(n_166),
.B2(n_167),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_209),
.A2(n_202),
.B1(n_205),
.B2(n_199),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_211),
.B(n_213),
.C(n_8),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_198),
.B(n_148),
.Y(n_213)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_214),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_215),
.B(n_216),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_214),
.A2(n_206),
.B1(n_210),
.B2(n_10),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_217),
.A2(n_212),
.B(n_9),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_9),
.B(n_10),
.C(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_220),
.B(n_9),
.Y(n_221)
);


endmodule