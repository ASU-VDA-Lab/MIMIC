module fake_jpeg_11784_n_288 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_288);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_213;
wire n_153;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_30),
.B(n_0),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_57),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_26),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_70),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_62),
.Y(n_84)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_68),
.Y(n_87)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_1),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_63),
.A2(n_23),
.B1(n_39),
.B2(n_24),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_74),
.A2(n_106),
.B1(n_2),
.B2(n_3),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_79),
.B(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_57),
.B(n_32),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_86),
.Y(n_116)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_44),
.A2(n_42),
.B1(n_29),
.B2(n_39),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_104),
.B1(n_34),
.B2(n_36),
.Y(n_112)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_32),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_33),
.Y(n_119)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_103),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_42),
.B1(n_29),
.B2(n_35),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_37),
.B1(n_36),
.B2(n_28),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_107),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_74),
.A2(n_55),
.B1(n_61),
.B2(n_66),
.Y(n_109)
);

OAI21xp33_ASAP7_75t_SL g157 ( 
.A1(n_109),
.A2(n_112),
.B(n_115),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_35),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_110),
.B(n_131),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_34),
.B1(n_28),
.B2(n_37),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_67),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_118),
.C(n_78),
.Y(n_143)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_59),
.B1(n_69),
.B2(n_22),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_114),
.A2(n_95),
.B(n_99),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_90),
.B1(n_104),
.B2(n_87),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_125),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_29),
.B1(n_33),
.B2(n_4),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_77),
.B(n_91),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_94),
.A2(n_29),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_124),
.A2(n_128),
.B1(n_137),
.B2(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_18),
.Y(n_125)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_99),
.Y(n_126)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_17),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_134),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_2),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_6),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_133),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_6),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_14),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_83),
.B(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_136),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_83),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_88),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_143),
.B(n_145),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_118),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_167),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_169),
.Y(n_179)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_15),
.Y(n_155)
);

AOI322xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_120),
.A3(n_124),
.B1(n_126),
.B2(n_16),
.C1(n_129),
.C2(n_114),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_159),
.B(n_171),
.Y(n_180)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_110),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_128),
.A2(n_122),
.B(n_120),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_170),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_137),
.A2(n_100),
.B1(n_95),
.B2(n_92),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_16),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_182),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_185),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_117),
.B1(n_140),
.B2(n_123),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_184),
.A2(n_189),
.B1(n_192),
.B2(n_190),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_123),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_167),
.B(n_113),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_139),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_190),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_143),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_168),
.A2(n_139),
.B1(n_114),
.B2(n_129),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_150),
.B(n_113),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_7),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_160),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_166),
.A2(n_93),
.B1(n_97),
.B2(n_10),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_144),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_162),
.B(n_154),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_93),
.C(n_8),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_197),
.C(n_146),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_7),
.C(n_12),
.Y(n_197)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_182),
.B(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_203),
.B(n_209),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_205),
.Y(n_222)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_178),
.A2(n_152),
.B(n_170),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_214),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_183),
.A2(n_169),
.B(n_147),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_178),
.B(n_189),
.Y(n_228)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_208),
.B(n_210),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_177),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_191),
.Y(n_213)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_217),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_165),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_195),
.C(n_186),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_160),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_218),
.B(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_198),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_236),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_234),
.C(n_237),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_228),
.A2(n_215),
.B(n_211),
.Y(n_243)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_181),
.A3(n_185),
.B1(n_187),
.B2(n_194),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_231),
.A2(n_199),
.B(n_213),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_184),
.Y(n_234)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_198),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_193),
.C(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_209),
.C(n_202),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_243),
.B(n_246),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_226),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_248),
.C(n_249),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_205),
.B1(n_236),
.B2(n_228),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_227),
.B1(n_232),
.B2(n_230),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_224),
.A2(n_220),
.B(n_205),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_226),
.Y(n_247)
);

AO221x1_ASAP7_75t_L g256 ( 
.A1(n_247),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.C(n_229),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_199),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_211),
.C(n_201),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_217),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_221),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_200),
.C(n_208),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_233),
.C(n_229),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_259),
.C(n_248),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_240),
.A2(n_222),
.B(n_235),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_255),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_257),
.A2(n_258),
.B1(n_225),
.B2(n_261),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_244),
.A2(n_235),
.B(n_251),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_239),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_235),
.B(n_192),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_261),
.A2(n_249),
.B1(n_197),
.B2(n_239),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_263),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_264),
.A2(n_269),
.B1(n_174),
.B2(n_196),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_153),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_214),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_267),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_252),
.A2(n_219),
.B1(n_210),
.B2(n_180),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_253),
.B(n_155),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_193),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_269),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_265),
.B1(n_266),
.B2(n_262),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_274),
.B(n_264),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_278),
.B(n_271),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_282),
.B(n_164),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_276),
.A2(n_273),
.B(n_161),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_277),
.C(n_146),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_283),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_280),
.C(n_284),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_164),
.Y(n_288)
);


endmodule