module fake_jpeg_5429_n_32 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_32);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_32;

wire n_21;
wire n_23;
wire n_27;
wire n_22;
wire n_19;
wire n_20;
wire n_18;
wire n_30;
wire n_24;
wire n_28;
wire n_26;
wire n_25;
wire n_17;
wire n_31;
wire n_29;

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

AND2x2_ASAP7_75t_SL g18 ( 
.A(n_0),
.B(n_11),
.Y(n_18)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_7),
.B1(n_10),
.B2(n_4),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_13),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_18),
.B(n_8),
.Y(n_25)
);

NOR4xp25_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_26),
.C(n_27),
.D(n_17),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_22),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_19),
.B1(n_29),
.B2(n_23),
.Y(n_32)
);


endmodule