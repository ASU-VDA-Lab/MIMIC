module fake_jpeg_17043_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_3),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_8),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_11),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_0),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_64),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_54),
.B1(n_61),
.B2(n_57),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_80),
.A2(n_89),
.B1(n_63),
.B2(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_77),
.B(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_84),
.A2(n_92),
.B1(n_58),
.B2(n_68),
.Y(n_104)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_54),
.B1(n_61),
.B2(n_57),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_66),
.B1(n_67),
.B2(n_63),
.Y(n_92)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_55),
.Y(n_94)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_83),
.Y(n_97)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_110),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_108),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_51),
.B1(n_62),
.B2(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_59),
.B1(n_50),
.B2(n_48),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_21),
.B1(n_45),
.B2(n_44),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_112),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_19),
.B1(n_42),
.B2(n_41),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_82),
.A2(n_15),
.B1(n_39),
.B2(n_38),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_14),
.B1(n_37),
.B2(n_34),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_118),
.Y(n_133)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_105),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_128),
.A2(n_132),
.B1(n_109),
.B2(n_98),
.Y(n_136)
);

INVx2_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_136),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_126),
.A2(n_112),
.B1(n_103),
.B2(n_102),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_135),
.A2(n_139),
.B1(n_127),
.B2(n_132),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_131),
.B(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_122),
.A2(n_100),
.B1(n_118),
.B2(n_3),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_138),
.Y(n_140)
);

FAx1_ASAP7_75t_SL g139 ( 
.A(n_123),
.B(n_46),
.CI(n_33),
.CON(n_139),
.SN(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_143),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_133),
.B(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_144),
.A2(n_128),
.B(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_145),
.A2(n_147),
.B1(n_148),
.B2(n_120),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g146 ( 
.A(n_144),
.B(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_150),
.C(n_143),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_125),
.B1(n_139),
.B2(n_121),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_141),
.A2(n_139),
.B1(n_121),
.B2(n_120),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_142),
.A2(n_130),
.B(n_17),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_146),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_155),
.C(n_1),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_1),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_155),
.B1(n_29),
.B2(n_27),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_159),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_161),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_157),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_160),
.B1(n_133),
.B2(n_124),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_164),
.A2(n_124),
.B1(n_32),
.B2(n_30),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_25),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_24),
.C(n_22),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_167),
.A2(n_11),
.B(n_4),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_10),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_2),
.B(n_5),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_2),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_5),
.C(n_6),
.Y(n_172)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_6),
.B(n_7),
.Y(n_173)
);


endmodule