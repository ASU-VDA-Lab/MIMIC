module real_jpeg_703_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_0),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_0),
.A2(n_36),
.B1(n_38),
.B2(n_193),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_0),
.A2(n_69),
.B1(n_70),
.B2(n_193),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_0),
.A2(n_59),
.B1(n_64),
.B2(n_193),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_1),
.A2(n_44),
.B1(n_69),
.B2(n_70),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_1),
.A2(n_36),
.B1(n_38),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_1),
.A2(n_44),
.B1(n_59),
.B2(n_64),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_41),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_41),
.B1(n_69),
.B2(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_3),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_6),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_6),
.A2(n_36),
.B1(n_38),
.B2(n_140),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_6),
.A2(n_69),
.B1(n_70),
.B2(n_140),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_59),
.B1(n_64),
.B2(n_140),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_7),
.B(n_29),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_39),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_29),
.B(n_183),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_7),
.B(n_93),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g252 ( 
.A1(n_7),
.A2(n_38),
.B(n_253),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_7),
.B(n_59),
.C(n_73),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_7),
.A2(n_69),
.B1(n_70),
.B2(n_219),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_7),
.B(n_61),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_7),
.B(n_77),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_8),
.A2(n_36),
.B1(n_38),
.B2(n_68),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_59),
.B1(n_64),
.B2(n_68),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_9),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_9),
.A2(n_36),
.B1(n_38),
.B2(n_82),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_9),
.A2(n_69),
.B1(n_70),
.B2(n_82),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_59),
.B1(n_64),
.B2(n_82),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_14),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_14),
.A2(n_36),
.B1(n_38),
.B2(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_84),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_L g210 ( 
.A1(n_14),
.A2(n_59),
.B1(n_64),
.B2(n_84),
.Y(n_210)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_16),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_17),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_17),
.A2(n_36),
.B1(n_38),
.B2(n_174),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_17),
.A2(n_69),
.B1(n_70),
.B2(n_174),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_17),
.A2(n_59),
.B1(n_64),
.B2(n_174),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_18),
.A2(n_36),
.B1(n_38),
.B2(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_18),
.A2(n_29),
.B1(n_30),
.B2(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_18),
.A2(n_69),
.B1(n_70),
.B2(n_90),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_18),
.A2(n_59),
.B1(n_64),
.B2(n_90),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_39),
.B(n_40),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_27),
.A2(n_39),
.B1(n_139),
.B2(n_173),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_27),
.A2(n_39),
.B1(n_43),
.B2(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_34),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_30),
.A2(n_34),
.A3(n_38),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_32),
.B(n_36),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_35),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_35),
.A2(n_80),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_35),
.A2(n_80),
.B1(n_81),
.B2(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_35),
.A2(n_80),
.B1(n_103),
.B2(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_35),
.A2(n_80),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_35),
.A2(n_80),
.B1(n_192),
.B2(n_231),
.Y(n_230)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_36),
.A2(n_38),
.B1(n_94),
.B2(n_95),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_36),
.B(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g217 ( 
.A1(n_38),
.A2(n_69),
.A3(n_94),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_42),
.B(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_46),
.B(n_330),
.Y(n_329)
);

OAI21x1_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_326),
.B(n_328),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_314),
.B(n_325),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_154),
.B(n_311),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_141),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_114),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_52),
.B(n_114),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_85),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_53),
.B(n_100),
.C(n_112),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_78),
.B(n_79),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_54),
.A2(n_55),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_65),
.Y(n_55)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_56),
.A2(n_78),
.B1(n_79),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_56),
.A2(n_65),
.B1(n_66),
.B2(n_78),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_62),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_57),
.A2(n_60),
.B1(n_128),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_57),
.A2(n_60),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_57),
.A2(n_60),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_58),
.A2(n_61),
.B1(n_63),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_58),
.A2(n_61),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_58),
.A2(n_61),
.B1(n_186),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_58),
.A2(n_61),
.B1(n_223),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_58),
.A2(n_61),
.B1(n_219),
.B2(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_58),
.A2(n_61),
.B1(n_273),
.B2(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_59),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_64),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_59),
.B(n_271),
.Y(n_270)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_67),
.A2(n_71),
.B1(n_77),
.B2(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_69),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_70),
.B1(n_94),
.B2(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_69),
.B(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_70),
.B(n_95),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_77),
.B(n_99),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_71),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_71),
.A2(n_77),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_71),
.A2(n_77),
.B1(n_215),
.B2(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_71),
.A2(n_77),
.B1(n_243),
.B2(n_244),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_71),
.A2(n_77),
.B1(n_243),
.B2(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_75),
.A2(n_132),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_75),
.A2(n_167),
.B1(n_214),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_100),
.B1(n_112),
.B2(n_113),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g121 ( 
.A1(n_86),
.A2(n_87),
.B(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_98),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B1(n_93),
.B2(n_97),
.Y(n_87)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_89),
.A2(n_92),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_93),
.B1(n_97),
.B2(n_109),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_91),
.A2(n_93),
.B1(n_135),
.B2(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_91),
.A2(n_93),
.B(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_92),
.A2(n_110),
.B1(n_136),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_92),
.A2(n_136),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_92),
.A2(n_136),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_92),
.A2(n_136),
.B1(n_189),
.B2(n_205),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_92),
.A2(n_136),
.B1(n_204),
.B2(n_252),
.Y(n_251)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_96),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_102),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_102),
.B(n_106),
.C(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_102),
.B(n_145),
.C(n_152),
.Y(n_315)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_108),
.B2(n_111),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_106),
.A2(n_111),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_106),
.B(n_148),
.C(n_150),
.Y(n_324)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.C(n_122),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_133),
.C(n_137),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_124),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_137),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_141),
.A2(n_312),
.B(n_313),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_153),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_142),
.B(n_153),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_149),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g321 ( 
.A(n_151),
.Y(n_321)
);

AO21x1_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_175),
.B(n_310),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_156),
.B(n_158),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.C(n_163),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_160),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_197),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.C(n_172),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_165),
.B(n_168),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_166),
.Y(n_235)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_172),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g190 ( 
.A(n_171),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_198),
.B(n_309),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_196),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_177),
.B(n_196),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_180),
.C(n_195),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_178),
.B(n_195),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_180),
.B(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_188),
.C(n_191),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_181),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_185),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_188),
.B(n_191),
.Y(n_299)
);

AOI31xp33_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_293),
.A3(n_302),
.B(n_306),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_238),
.B(n_292),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_225),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_201),
.B(n_225),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_212),
.C(n_216),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_202),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_207),
.C(n_211),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_212),
.B(n_216),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_228),
.C(n_229),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_233),
.C(n_237),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_233),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_239),
.A2(n_287),
.B(n_291),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_256),
.B(n_286),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_248),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_246),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_242),
.B(n_245),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_247),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_267),
.B(n_285),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_265),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_265),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_279),
.B(n_284),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B(n_278),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_297),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_303),
.B(n_304),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_316),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_318),
.A2(n_320),
.B1(n_322),
.B2(n_323),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_327),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule