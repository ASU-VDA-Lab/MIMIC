module real_aes_2427_n_16 (n_13, n_4, n_0, n_3, n_5, n_2, n_15, n_7, n_8, n_6, n_9, n_12, n_1, n_14, n_10, n_11, n_16);
input n_13;
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_15;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_14;
input n_10;
input n_11;
output n_16;
wire n_17;
wire n_28;
wire n_22;
wire n_24;
wire n_41;
wire n_56;
wire n_34;
wire n_55;
wire n_19;
wire n_40;
wire n_49;
wire n_46;
wire n_53;
wire n_25;
wire n_47;
wire n_48;
wire n_43;
wire n_32;
wire n_30;
wire n_37;
wire n_51;
wire n_54;
wire n_35;
wire n_42;
wire n_39;
wire n_45;
wire n_27;
wire n_23;
wire n_38;
wire n_50;
wire n_29;
wire n_20;
wire n_52;
wire n_57;
wire n_44;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
CKINVDCx20_ASAP7_75t_R g53 ( .A(n_0), .Y(n_53) );
AOI221xp5_ASAP7_75t_SL g36 ( .A1(n_1), .A2(n_13), .B1(n_37), .B2(n_48), .C(n_51), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g26 ( .A(n_2), .Y(n_26) );
NOR3xp33_ASAP7_75t_SL g24 ( .A(n_3), .B(n_7), .C(n_25), .Y(n_24) );
CKINVDCx5p33_ASAP7_75t_R g25 ( .A(n_4), .Y(n_25) );
CKINVDCx20_ASAP7_75t_R g32 ( .A(n_5), .Y(n_32) );
NAND3xp33_ASAP7_75t_SL g28 ( .A(n_6), .B(n_29), .C(n_30), .Y(n_28) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_6), .B(n_23), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g31 ( .A(n_8), .Y(n_31) );
NOR2xp33_ASAP7_75t_R g47 ( .A(n_8), .B(n_12), .Y(n_47) );
CKINVDCx20_ASAP7_75t_R g57 ( .A(n_9), .Y(n_57) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_10), .Y(n_29) );
NOR2xp33_ASAP7_75t_R g45 ( .A(n_10), .B(n_46), .Y(n_45) );
NOR2xp33_ASAP7_75t_R g30 ( .A(n_11), .B(n_31), .Y(n_30) );
CKINVDCx20_ASAP7_75t_R g43 ( .A(n_11), .Y(n_43) );
NAND2xp33_ASAP7_75t_SL g18 ( .A(n_12), .B(n_19), .Y(n_18) );
NAND2xp33_ASAP7_75t_SL g33 ( .A(n_12), .B(n_34), .Y(n_33) );
NOR2xp33_ASAP7_75t_R g50 ( .A(n_12), .B(n_20), .Y(n_50) );
CKINVDCx20_ASAP7_75t_R g56 ( .A(n_12), .Y(n_56) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_14), .Y(n_27) );
NAND2xp33_ASAP7_75t_SL g35 ( .A(n_14), .B(n_22), .Y(n_35) );
NAND2xp33_ASAP7_75t_SL g52 ( .A(n_14), .B(n_41), .Y(n_52) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_15), .Y(n_17) );
OAI221xp5_ASAP7_75t_R g16 ( .A1(n_17), .A2(n_18), .B1(n_32), .B2(n_33), .C(n_36), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_20), .Y(n_19) );
OR2x2_ASAP7_75t_L g20 ( .A(n_21), .B(n_28), .Y(n_20) );
NAND2xp33_ASAP7_75t_SL g21 ( .A(n_22), .B(n_27), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_23), .Y(n_22) );
NAND2xp33_ASAP7_75t_SL g23 ( .A(n_24), .B(n_26), .Y(n_23) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_27), .B(n_41), .Y(n_40) );
NOR2xp33_ASAP7_75t_R g34 ( .A(n_28), .B(n_35), .Y(n_34) );
NAND2xp33_ASAP7_75t_SL g55 ( .A(n_34), .B(n_56), .Y(n_55) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_39), .B(n_42), .Y(n_38) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
CKINVDCx20_ASAP7_75t_R g54 ( .A(n_42), .Y(n_54) );
NOR2xp33_ASAP7_75t_R g42 ( .A(n_43), .B(n_44), .Y(n_42) );
CKINVDCx20_ASAP7_75t_R g44 ( .A(n_45), .Y(n_44) );
CKINVDCx14_ASAP7_75t_R g46 ( .A(n_47), .Y(n_46) );
CKINVDCx20_ASAP7_75t_R g48 ( .A(n_49), .Y(n_48) );
INVx1_ASAP7_75t_L g49 ( .A(n_50), .Y(n_49) );
OAI32xp33_ASAP7_75t_L g51 ( .A1(n_52), .A2(n_53), .A3(n_54), .B1(n_55), .B2(n_57), .Y(n_51) );
endmodule