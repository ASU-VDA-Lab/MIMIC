module real_jpeg_17916_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_0),
.Y(n_252)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_1),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_1),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_2),
.A2(n_136),
.B1(n_140),
.B2(n_141),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_2),
.Y(n_140)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_3),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_3),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_4),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_4),
.A2(n_53),
.B1(n_90),
.B2(n_93),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_53),
.B1(n_153),
.B2(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_4),
.B(n_215),
.Y(n_214)
);

OAI32xp33_ASAP7_75t_L g281 ( 
.A1(n_4),
.A2(n_282),
.A3(n_285),
.B1(n_286),
.B2(n_291),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_4),
.B(n_109),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_4),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_4),
.B(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_5),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_5),
.Y(n_204)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_5),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22x1_ASAP7_75t_L g101 ( 
.A1(n_6),
.A2(n_35),
.B1(n_102),
.B2(n_106),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_6),
.A2(n_35),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_6),
.A2(n_35),
.B1(n_307),
.B2(n_310),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_7),
.A2(n_119),
.B1(n_120),
.B2(n_124),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_7),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_7),
.B(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_7),
.A2(n_119),
.B1(n_197),
.B2(n_201),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_7),
.A2(n_119),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_10),
.Y(n_139)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_11),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_233),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_231),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_189),
.Y(n_14)
);

NOR2xp67_ASAP7_75t_L g232 ( 
.A(n_15),
.B(n_189),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_133),
.C(n_174),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_16),
.B(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_59),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_17),
.B(n_60),
.C(n_99),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_40),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_19),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x4_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_20),
.B(n_53),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_22),
.Y(n_129)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_22),
.Y(n_216)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_23),
.Y(n_132)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_23),
.Y(n_164)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_26),
.Y(n_171)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_28),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_30),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_31),
.B(n_41),
.Y(n_230)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_37),
.Y(n_229)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_52),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_46),
.B1(n_49),
.B2(n_51),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_45),
.Y(n_167)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_53),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_53),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_53),
.B(n_287),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_56),
.A2(n_161),
.B1(n_165),
.B2(n_172),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_98),
.B2(n_99),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_75),
.B(n_89),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_62),
.B(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_62),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_62),
.B(n_269),
.Y(n_299)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_70),
.B2(n_74),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_69),
.Y(n_290)
);

INVx5_ASAP7_75t_L g309 ( 
.A(n_69),
.Y(n_309)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_72),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_73),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_75),
.B(n_89),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_75),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_75),
.B(n_196),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_79),
.B1(n_82),
.B2(n_86),
.Y(n_76)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_77),
.Y(n_272)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_86),
.Y(n_270)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_87),
.Y(n_284)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_89),
.Y(n_266)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_117),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_100),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_109),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_101),
.B(n_125),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2x1p5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_109),
.B(n_118),
.Y(n_177)
);

NAND2xp33_ASAP7_75t_SL g212 ( 
.A(n_109),
.B(n_213),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_127),
.B1(n_130),
.B2(n_131),
.Y(n_126)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

O2A1O1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_119),
.A2(n_142),
.B(n_156),
.C(n_187),
.Y(n_186)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_125),
.Y(n_355)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_133),
.A2(n_174),
.B1(n_175),
.B2(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_133),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_160),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_134),
.B(n_160),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_142),
.B(n_147),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_135),
.A2(n_149),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_139),
.Y(n_312)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_145),
.Y(n_304)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_147),
.B(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_156),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_149),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_149),
.B(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_155),
.Y(n_325)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_172),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.C(n_180),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_176),
.B(n_239),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_178),
.B(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_179),
.Y(n_240)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_182),
.B(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_183),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_186),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g333 ( 
.A(n_186),
.B(n_305),
.Y(n_333)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_207),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_206),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp67_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_195),
.B(n_268),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_205),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_220),
.B2(n_221),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_213),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_217),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

OAI32xp33_ASAP7_75t_L g242 ( 
.A1(n_217),
.A2(n_243),
.A3(n_244),
.B1(n_247),
.B2(n_253),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_276),
.B(n_368),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_273),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_237),
.B(n_273),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_241),
.C(n_262),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_238),
.B(n_364),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_241),
.A2(n_262),
.B1(n_263),
.B2(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_241),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_257),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_242),
.A2(n_257),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_242),
.Y(n_358)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_257),
.Y(n_357)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_260),
.B(n_261),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AO21x1_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_302),
.B(n_305),
.Y(n_301)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_362),
.B(n_367),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_343),
.B(n_361),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_318),
.B(n_342),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_300),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_L g342 ( 
.A(n_280),
.B(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_298),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_298),
.Y(n_340)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

INVx5_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_299),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.Y(n_300)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_301),
.Y(n_360)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_303),
.B(n_306),
.Y(n_331)
);

INVx4_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_315),
.B(n_316),
.C(n_360),
.Y(n_359)
);

OAI21x1_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_337),
.B(n_341),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_332),
.B(n_336),
.Y(n_319)
);

NOR2x1_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_330),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_326),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_331),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_333),
.B(n_334),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_338),
.B(n_340),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_359),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_359),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_356),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_346),
.B(n_351),
.C(n_356),
.Y(n_366)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

NOR2x1_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_363),
.B(n_366),
.Y(n_367)
);


endmodule