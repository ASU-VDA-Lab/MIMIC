module fake_netlist_6_2932_n_1038 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1038);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1038;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_1026;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_718;
wire n_517;
wire n_1018;
wire n_852;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_842;
wire n_525;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_953;
wire n_886;
wire n_1004;
wire n_1017;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_930;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_196;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_779;
wire n_800;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_939;
wire n_819;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_1034;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_956;
wire n_960;
wire n_531;
wire n_827;
wire n_1001;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1025;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_194;
wire n_664;
wire n_949;
wire n_678;
wire n_192;
wire n_1007;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_83),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_101),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_80),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_51),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_139),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_25),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_19),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_15),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_17),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_184),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_30),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_25),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_60),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_22),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_179),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_109),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_88),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_36),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_82),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_18),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_128),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_158),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_68),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_156),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_8),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_33),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_69),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_28),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_160),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_0),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_93),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_76),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_67),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_19),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_89),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_114),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_90),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_48),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_2),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_127),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_43),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_138),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_74),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_77),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_165),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_9),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_143),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_169),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_151),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_163),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_194),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_231),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_193),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_225),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_230),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_224),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_232),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_237),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_196),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_219),
.Y(n_269)
);

BUFx2_ASAP7_75t_SL g270 ( 
.A(n_207),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_193),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_199),
.Y(n_273)
);

INVxp33_ASAP7_75t_SL g274 ( 
.A(n_201),
.Y(n_274)
);

NOR2xp67_ASAP7_75t_L g275 ( 
.A(n_190),
.B(n_0),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_205),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_226),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_229),
.Y(n_279)
);

INVxp33_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_189),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_206),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_221),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_212),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_187),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_245),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_246),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_190),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_187),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_254),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_225),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_191),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_191),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_192),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_192),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_303),
.Y(n_306)
);

OA21x2_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_218),
.B(n_202),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_305),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_242),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_294),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_294),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_197),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_302),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_270),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_261),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

OA21x2_ASAP7_75t_L g321 ( 
.A1(n_283),
.A2(n_286),
.B(n_284),
.Y(n_321)
);

CKINVDCx6p67_ASAP7_75t_R g322 ( 
.A(n_262),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_260),
.A2(n_207),
.B1(n_253),
.B2(n_220),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_253),
.B(n_200),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_288),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_265),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_291),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_198),
.Y(n_330)
);

BUFx8_ASAP7_75t_L g331 ( 
.A(n_276),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_293),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_295),
.Y(n_333)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_296),
.A2(n_208),
.B(n_204),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_289),
.Y(n_336)
);

AND2x4_ASAP7_75t_L g337 ( 
.A(n_272),
.B(n_203),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_298),
.Y(n_338)
);

AND2x4_ASAP7_75t_L g339 ( 
.A(n_275),
.B(n_203),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_258),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_268),
.A2(n_211),
.B(n_210),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_259),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_264),
.B(n_213),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_282),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_217),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_304),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_304),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

AND2x4_ASAP7_75t_L g349 ( 
.A(n_278),
.B(n_213),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_279),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_223),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_267),
.Y(n_352)
);

OAI21x1_ASAP7_75t_L g353 ( 
.A1(n_273),
.A2(n_222),
.B(n_213),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_279),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_257),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_274),
.B(n_227),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_L g358 ( 
.A(n_257),
.B(n_213),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_256),
.A2(n_222),
.B1(n_252),
.B2(n_248),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_274),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_318),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_R g362 ( 
.A(n_318),
.B(n_336),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_228),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_322),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_352),
.B(n_233),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_322),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_336),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_331),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_355),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_357),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_280),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_360),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_360),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_360),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_360),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_360),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_355),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_355),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_280),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_344),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_355),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_328),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_347),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_347),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_321),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_R g395 ( 
.A(n_348),
.B(n_260),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_347),
.Y(n_396)
);

INVx8_ASAP7_75t_L g397 ( 
.A(n_347),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_327),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_317),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_323),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_327),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_347),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_327),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_344),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_350),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_356),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_350),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_346),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_327),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_354),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_348),
.A2(n_240),
.B1(n_234),
.B2(n_235),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_316),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_346),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_356),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_359),
.A2(n_292),
.B1(n_285),
.B2(n_271),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_314),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_351),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_343),
.B(n_236),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_333),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_327),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_330),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_330),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_341),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_343),
.B(n_239),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_317),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_343),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_310),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_358),
.B(n_271),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_394),
.B(n_341),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_341),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_368),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_374),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_397),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_324),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_428),
.B(n_309),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_377),
.Y(n_441)
);

AND2x2_ASAP7_75t_SL g442 ( 
.A(n_405),
.B(n_324),
.Y(n_442)
);

BUFx4f_ASAP7_75t_L g443 ( 
.A(n_397),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_L g444 ( 
.A1(n_378),
.A2(n_342),
.B1(n_340),
.B2(n_324),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_385),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_391),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_392),
.B(n_309),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_397),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_427),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_393),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_418),
.B(n_334),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_361),
.B(n_285),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_406),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_364),
.B(n_342),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_425),
.A2(n_334),
.B1(n_307),
.B2(n_310),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_408),
.Y(n_465)
);

OAI21xp33_ASAP7_75t_L g466 ( 
.A1(n_379),
.A2(n_310),
.B(n_340),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_427),
.Y(n_467)
);

AND2x4_ASAP7_75t_SL g468 ( 
.A(n_365),
.B(n_292),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_375),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_L g471 ( 
.A1(n_425),
.A2(n_334),
.B1(n_307),
.B2(n_310),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_SL g472 ( 
.A(n_396),
.B(n_247),
.C(n_241),
.Y(n_472)
);

AND2x6_ASAP7_75t_L g473 ( 
.A(n_372),
.B(n_222),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_401),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_410),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_414),
.B(n_334),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_395),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_367),
.B(n_340),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_402),
.B(n_309),
.Y(n_479)
);

BUFx10_ASAP7_75t_L g480 ( 
.A(n_369),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_412),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_403),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_411),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_388),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_386),
.B(n_387),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_381),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_422),
.B(n_353),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_362),
.Y(n_490)
);

OR2x6_ASAP7_75t_L g491 ( 
.A(n_417),
.B(n_353),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_423),
.B(n_222),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_429),
.Y(n_493)
);

INVx4_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_424),
.B(n_335),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_420),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_384),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_370),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_415),
.B(n_421),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_413),
.B(n_337),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_431),
.B(n_339),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_371),
.B(n_255),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_416),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_407),
.B(n_320),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_407),
.B(n_321),
.Y(n_507)
);

AND2x6_ASAP7_75t_L g508 ( 
.A(n_400),
.B(n_337),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_400),
.B(n_339),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_373),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_363),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_363),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_460),
.B(n_320),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_435),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_511),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_507),
.A2(n_491),
.B1(n_460),
.B2(n_484),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_450),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_433),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_320),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_470),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_441),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_438),
.B(n_449),
.Y(n_522)
);

AND2x4_ASAP7_75t_L g523 ( 
.A(n_437),
.B(n_486),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_445),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_461),
.B(n_326),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_446),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_464),
.B(n_326),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_506),
.Y(n_529)
);

OAI221xp5_ASAP7_75t_L g530 ( 
.A1(n_507),
.A2(n_321),
.B1(n_332),
.B2(n_329),
.C(n_338),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_512),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_465),
.B(n_475),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_488),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_456),
.B(n_321),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_493),
.Y(n_535)
);

NAND2x1p5_ASAP7_75t_L g536 ( 
.A(n_449),
.B(n_453),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_439),
.B(n_332),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_476),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_499),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_476),
.A2(n_335),
.B1(n_329),
.B2(n_307),
.Y(n_541)
);

INVxp67_ASAP7_75t_L g542 ( 
.A(n_496),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_447),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_454),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_452),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_469),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_492),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_439),
.B(n_312),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_455),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_462),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_478),
.B(n_312),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_432),
.B(n_312),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_498),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_495),
.Y(n_557)
);

AO22x2_ASAP7_75t_L g558 ( 
.A1(n_492),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_481),
.B(n_477),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_490),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_457),
.B(n_313),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_455),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_457),
.B(n_313),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_467),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_458),
.A2(n_317),
.B1(n_308),
.B2(n_315),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_485),
.B(n_4),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_487),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_466),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_494),
.B(n_311),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_480),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_555),
.A2(n_443),
.B(n_453),
.Y(n_574)
);

AND3x2_ASAP7_75t_L g575 ( 
.A(n_556),
.B(n_459),
.C(n_510),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_542),
.B(n_496),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_524),
.Y(n_577)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_534),
.A2(n_434),
.B(n_432),
.Y(n_578)
);

A2O1A1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_568),
.A2(n_497),
.B(n_458),
.C(n_485),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_523),
.B(n_489),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_520),
.B(n_480),
.Y(n_581)
);

NAND3xp33_ASAP7_75t_L g582 ( 
.A(n_532),
.B(n_505),
.C(n_504),
.Y(n_582)
);

INVx1_ASAP7_75t_SL g583 ( 
.A(n_533),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_553),
.B(n_533),
.Y(n_584)
);

O2A1O1Ixp5_ASAP7_75t_L g585 ( 
.A1(n_513),
.A2(n_444),
.B(n_502),
.C(n_448),
.Y(n_585)
);

INVx6_ASAP7_75t_L g586 ( 
.A(n_523),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_536),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_557),
.B(n_562),
.Y(n_588)
);

AOI21xp5_ASAP7_75t_L g589 ( 
.A1(n_554),
.A2(n_479),
.B(n_448),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_559),
.B(n_509),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_519),
.B(n_489),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_528),
.B(n_509),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_540),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_565),
.B(n_501),
.Y(n_594)
);

BUFx8_ASAP7_75t_SL g595 ( 
.A(n_560),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g596 ( 
.A1(n_551),
.A2(n_440),
.B(n_442),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g597 ( 
.A1(n_534),
.A2(n_471),
.B(n_463),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_536),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_529),
.B(n_468),
.Y(n_599)
);

A2O1A1Ixp33_ASAP7_75t_L g600 ( 
.A1(n_570),
.A2(n_501),
.B(n_463),
.C(n_471),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g601 ( 
.A1(n_537),
.A2(n_444),
.B(n_467),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_573),
.B(n_547),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_569),
.A2(n_522),
.B(n_530),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_562),
.Y(n_604)
);

INVxp67_ASAP7_75t_SL g605 ( 
.A(n_547),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_517),
.Y(n_606)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_530),
.A2(n_467),
.B(n_472),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_514),
.B(n_508),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_564),
.B(n_508),
.Y(n_609)
);

AOI21x1_ASAP7_75t_L g610 ( 
.A1(n_549),
.A2(n_503),
.B(n_473),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_515),
.B(n_508),
.Y(n_611)
);

OAI21xp5_ASAP7_75t_L g612 ( 
.A1(n_541),
.A2(n_473),
.B(n_508),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_564),
.B(n_571),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_516),
.A2(n_473),
.B1(n_306),
.B2(n_92),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_526),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_518),
.B(n_5),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_5),
.C(n_6),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_571),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_L g619 ( 
.A1(n_525),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_527),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_552),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_531),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_546),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_590),
.B(n_535),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g626 ( 
.A1(n_601),
.A2(n_567),
.B(n_538),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_583),
.B(n_588),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_576),
.B(n_539),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_622),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_615),
.B(n_543),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_584),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_585),
.A2(n_544),
.B(n_548),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_588),
.B(n_552),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_594),
.A2(n_563),
.B1(n_561),
.B2(n_572),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_620),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_592),
.B(n_550),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_579),
.A2(n_566),
.B(n_558),
.C(n_550),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_595),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_624),
.Y(n_639)
);

INVx5_ASAP7_75t_L g640 ( 
.A(n_577),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_581),
.B(n_558),
.Y(n_641)
);

O2A1O1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_582),
.A2(n_558),
.B(n_9),
.C(n_10),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_589),
.A2(n_32),
.B(n_31),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_608),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_621),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_605),
.B(n_11),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_591),
.B(n_13),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_606),
.Y(n_648)
);

OAI22xp5_ASAP7_75t_L g649 ( 
.A1(n_611),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_SL g650 ( 
.A(n_599),
.B(n_18),
.C(n_20),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_623),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_623),
.Y(n_652)
);

O2A1O1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_619),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_653)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_600),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_593),
.A2(n_24),
.B1(n_26),
.B2(n_27),
.Y(n_655)
);

A2O1A1Ixp33_ASAP7_75t_L g656 ( 
.A1(n_596),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_656)
);

AOI21x1_ASAP7_75t_L g657 ( 
.A1(n_607),
.A2(n_183),
.B(n_103),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_578),
.A2(n_102),
.B(n_178),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_580),
.B(n_181),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_616),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_613),
.B(n_29),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_580),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_604),
.B(n_177),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_617),
.A2(n_34),
.B(n_35),
.C(n_37),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_609),
.B(n_38),
.Y(n_665)
);

O2A1O1Ixp33_ASAP7_75t_L g666 ( 
.A1(n_612),
.A2(n_40),
.B(n_41),
.C(n_44),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_604),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_667)
);

INVx4_ASAP7_75t_L g668 ( 
.A(n_577),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_602),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_SL g670 ( 
.A1(n_614),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_670)
);

OA22x2_ASAP7_75t_L g671 ( 
.A1(n_575),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_618),
.B(n_56),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_602),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_587),
.B(n_57),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_622),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_603),
.A2(n_58),
.B(n_59),
.C(n_61),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_640),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_639),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_629),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_640),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_635),
.Y(n_682)
);

BUFx6f_ASAP7_75t_SL g683 ( 
.A(n_668),
.Y(n_683)
);

BUFx4f_ASAP7_75t_SL g684 ( 
.A(n_668),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_631),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_659),
.B(n_587),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_640),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_673),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_628),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_662),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_645),
.Y(n_691)
);

BUFx4f_ASAP7_75t_SL g692 ( 
.A(n_662),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_625),
.Y(n_693)
);

CKINVDCx8_ASAP7_75t_R g694 ( 
.A(n_638),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_662),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_659),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_654),
.A2(n_597),
.B1(n_587),
.B2(n_598),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_669),
.Y(n_698)
);

INVx8_ASAP7_75t_L g699 ( 
.A(n_627),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_660),
.B(n_586),
.Y(n_700)
);

AOI22xp33_ASAP7_75t_L g701 ( 
.A1(n_655),
.A2(n_598),
.B1(n_586),
.B2(n_622),
.Y(n_701)
);

BUFx2_ASAP7_75t_SL g702 ( 
.A(n_651),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_630),
.Y(n_703)
);

BUFx4f_ASAP7_75t_SL g704 ( 
.A(n_652),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_647),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_661),
.Y(n_706)
);

INVx4_ASAP7_75t_L g707 ( 
.A(n_675),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_636),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_650),
.B(n_598),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_633),
.B(n_574),
.Y(n_710)
);

INVx4_ASAP7_75t_L g711 ( 
.A(n_671),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_646),
.B(n_610),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_626),
.Y(n_713)
);

INVx5_ASAP7_75t_SL g714 ( 
.A(n_667),
.Y(n_714)
);

INVx1_ASAP7_75t_SL g715 ( 
.A(n_665),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_657),
.Y(n_716)
);

BUFx6f_ASAP7_75t_SL g717 ( 
.A(n_663),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_672),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_634),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_632),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_641),
.B(n_62),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_644),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_674),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_642),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_656),
.Y(n_725)
);

INVx6_ASAP7_75t_L g726 ( 
.A(n_664),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_637),
.B(n_176),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_649),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_670),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_658),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_653),
.Y(n_731)
);

BUFx12f_ASAP7_75t_L g732 ( 
.A(n_666),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_676),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_643),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_718),
.B(n_63),
.Y(n_735)
);

HB1xp67_ASAP7_75t_L g736 ( 
.A(n_685),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_705),
.B(n_64),
.Y(n_737)
);

OAI21x1_ASAP7_75t_L g738 ( 
.A1(n_716),
.A2(n_734),
.B(n_710),
.Y(n_738)
);

OA21x2_ASAP7_75t_L g739 ( 
.A1(n_729),
.A2(n_66),
.B(n_70),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_693),
.B(n_71),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_696),
.B(n_690),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_696),
.B(n_72),
.Y(n_742)
);

OAI21x1_ASAP7_75t_L g743 ( 
.A1(n_710),
.A2(n_73),
.B(n_75),
.Y(n_743)
);

BUFx10_ASAP7_75t_L g744 ( 
.A(n_683),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_678),
.Y(n_745)
);

BUFx2_ASAP7_75t_L g746 ( 
.A(n_688),
.Y(n_746)
);

OAI21x1_ASAP7_75t_SL g747 ( 
.A1(n_727),
.A2(n_78),
.B(n_79),
.Y(n_747)
);

INVx3_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

NAND2x1p5_ASAP7_75t_L g749 ( 
.A(n_696),
.B(n_81),
.Y(n_749)
);

OAI221xp5_ASAP7_75t_L g750 ( 
.A1(n_701),
.A2(n_726),
.B1(n_731),
.B2(n_728),
.C(n_705),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_696),
.B(n_84),
.Y(n_751)
);

OAI21x1_ASAP7_75t_L g752 ( 
.A1(n_733),
.A2(n_85),
.B(n_86),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_679),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_677),
.Y(n_754)
);

BUFx2_ASAP7_75t_L g755 ( 
.A(n_690),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_689),
.B(n_87),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_691),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_708),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_695),
.Y(n_759)
);

OAI21xp5_ASAP7_75t_L g760 ( 
.A1(n_730),
.A2(n_94),
.B(n_95),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_701),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_682),
.Y(n_762)
);

OAI21xp5_ASAP7_75t_L g763 ( 
.A1(n_730),
.A2(n_99),
.B(n_100),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_721),
.A2(n_104),
.B(n_105),
.C(n_106),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_731),
.B(n_108),
.C(n_110),
.Y(n_765)
);

OAI21x1_ASAP7_75t_L g766 ( 
.A1(n_697),
.A2(n_111),
.B(n_112),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_715),
.B(n_113),
.Y(n_767)
);

OAI21x1_ASAP7_75t_L g768 ( 
.A1(n_697),
.A2(n_115),
.B(n_116),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_720),
.A2(n_117),
.B(n_118),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_706),
.Y(n_770)
);

INVx5_ASAP7_75t_L g771 ( 
.A(n_686),
.Y(n_771)
);

OAI21x1_ASAP7_75t_SL g772 ( 
.A1(n_711),
.A2(n_698),
.B(n_707),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_712),
.A2(n_119),
.B(n_120),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_698),
.B(n_121),
.Y(n_774)
);

BUFx12f_ASAP7_75t_SL g775 ( 
.A(n_700),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_699),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_703),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_681),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_706),
.Y(n_779)
);

AO32x2_ASAP7_75t_L g780 ( 
.A1(n_713),
.A2(n_122),
.A3(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_715),
.B(n_126),
.Y(n_781)
);

AO31x2_ASAP7_75t_L g782 ( 
.A1(n_713),
.A2(n_129),
.A3(n_130),
.B(n_131),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_711),
.B(n_132),
.Y(n_783)
);

OAI21x1_ASAP7_75t_L g784 ( 
.A1(n_680),
.A2(n_133),
.B(n_134),
.Y(n_784)
);

AOI221xp5_ASAP7_75t_L g785 ( 
.A1(n_731),
.A2(n_136),
.B1(n_137),
.B2(n_140),
.C(n_141),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_745),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_770),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_738),
.Y(n_788)
);

INVx6_ASAP7_75t_L g789 ( 
.A(n_771),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_779),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_753),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_736),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_758),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_757),
.Y(n_794)
);

CKINVDCx11_ASAP7_75t_R g795 ( 
.A(n_744),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_777),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_762),
.Y(n_797)
);

OA21x2_ASAP7_75t_L g798 ( 
.A1(n_752),
.A2(n_723),
.B(n_709),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_782),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_775),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_755),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_760),
.A2(n_732),
.B1(n_722),
.B2(n_726),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_772),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_748),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_746),
.B(n_724),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_771),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_773),
.A2(n_723),
.B(n_726),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_782),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_780),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_782),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_780),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_748),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_780),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_781),
.Y(n_814)
);

INVxp67_ASAP7_75t_SL g815 ( 
.A(n_781),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_719),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_743),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_756),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_756),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_740),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_739),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_741),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_739),
.Y(n_823)
);

CKINVDCx6p67_ASAP7_75t_R g824 ( 
.A(n_744),
.Y(n_824)
);

AOI22xp33_ASAP7_75t_L g825 ( 
.A1(n_760),
.A2(n_722),
.B1(n_724),
.B2(n_725),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_737),
.B(n_724),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_740),
.Y(n_827)
);

OR2x6_ASAP7_75t_L g828 ( 
.A(n_749),
.B(n_725),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_759),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_786),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_790),
.B(n_725),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_786),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_792),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_L g834 ( 
.A(n_802),
.B(n_825),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_787),
.B(n_776),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_800),
.B(n_750),
.C(n_763),
.Y(n_836)
);

AO31x2_ASAP7_75t_L g837 ( 
.A1(n_799),
.A2(n_761),
.A3(n_769),
.B(n_783),
.Y(n_837)
);

AOI21xp33_ASAP7_75t_L g838 ( 
.A1(n_807),
.A2(n_763),
.B(n_765),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_795),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_800),
.B(n_717),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_801),
.B(n_741),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_789),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_829),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_829),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_792),
.B(n_771),
.Y(n_845)
);

INVx6_ASAP7_75t_L g846 ( 
.A(n_828),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_821),
.A2(n_823),
.B(n_803),
.Y(n_847)
);

OR2x6_ASAP7_75t_L g848 ( 
.A(n_789),
.B(n_765),
.Y(n_848)
);

NAND2xp33_ASAP7_75t_R g849 ( 
.A(n_807),
.B(n_735),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_815),
.B(n_783),
.Y(n_850)
);

NAND2xp33_ASAP7_75t_R g851 ( 
.A(n_807),
.B(n_742),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_795),
.Y(n_852)
);

CKINVDCx16_ASAP7_75t_R g853 ( 
.A(n_826),
.Y(n_853)
);

NOR3xp33_ASAP7_75t_SL g854 ( 
.A(n_805),
.B(n_761),
.C(n_767),
.Y(n_854)
);

OR2x6_ASAP7_75t_L g855 ( 
.A(n_789),
.B(n_751),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_794),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_822),
.B(n_754),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_794),
.Y(n_858)
);

INVxp67_ASAP7_75t_L g859 ( 
.A(n_821),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_826),
.B(n_754),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_804),
.B(n_754),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_791),
.B(n_778),
.Y(n_862)
);

OR2x6_ASAP7_75t_L g863 ( 
.A(n_789),
.B(n_742),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_824),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_833),
.Y(n_865)
);

OR2x2_ASAP7_75t_L g866 ( 
.A(n_859),
.B(n_809),
.Y(n_866)
);

AO21x2_ASAP7_75t_L g867 ( 
.A1(n_838),
.A2(n_823),
.B(n_799),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_864),
.B(n_824),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_859),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_850),
.B(n_809),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_853),
.B(n_811),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_847),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_830),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_842),
.B(n_788),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_842),
.B(n_788),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_832),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_856),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_858),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_850),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_846),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_862),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_845),
.Y(n_882)
);

NAND4xp25_ASAP7_75t_L g883 ( 
.A(n_849),
.B(n_814),
.C(n_818),
.D(n_820),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_836),
.A2(n_714),
.B1(n_816),
.B2(n_828),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_831),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_841),
.B(n_811),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_835),
.Y(n_887)
);

CKINVDCx6p67_ASAP7_75t_R g888 ( 
.A(n_882),
.Y(n_888)
);

OA21x2_ASAP7_75t_L g889 ( 
.A1(n_872),
.A2(n_875),
.B(n_874),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_873),
.Y(n_890)
);

AOI211xp5_ASAP7_75t_L g891 ( 
.A1(n_883),
.A2(n_834),
.B(n_838),
.C(n_816),
.Y(n_891)
);

AO21x2_ASAP7_75t_L g892 ( 
.A1(n_872),
.A2(n_808),
.B(n_810),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_873),
.Y(n_893)
);

OAI211xp5_ASAP7_75t_L g894 ( 
.A1(n_884),
.A2(n_836),
.B(n_831),
.C(n_854),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_885),
.B(n_861),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_887),
.A2(n_848),
.B1(n_854),
.B2(n_846),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_880),
.A2(n_848),
.B1(n_714),
.B2(n_813),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_880),
.A2(n_848),
.B1(n_851),
.B2(n_828),
.Y(n_898)
);

INVx3_ASAP7_75t_L g899 ( 
.A(n_874),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_868),
.A2(n_764),
.B(n_840),
.C(n_785),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_866),
.Y(n_901)
);

OAI21xp33_ASAP7_75t_SL g902 ( 
.A1(n_871),
.A2(n_843),
.B(n_860),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_871),
.B(n_857),
.Y(n_903)
);

AND2x2_ASAP7_75t_L g904 ( 
.A(n_882),
.B(n_845),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_888),
.B(n_899),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_901),
.B(n_870),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_890),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_904),
.B(n_880),
.Y(n_908)
);

BUFx2_ASAP7_75t_L g909 ( 
.A(n_888),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_896),
.Y(n_910)
);

INVxp67_ASAP7_75t_SL g911 ( 
.A(n_889),
.Y(n_911)
);

INVx5_ASAP7_75t_SL g912 ( 
.A(n_892),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_893),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_889),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_889),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_899),
.B(n_885),
.Y(n_916)
);

INVxp67_ASAP7_75t_L g917 ( 
.A(n_894),
.Y(n_917)
);

NOR2x1_ASAP7_75t_L g918 ( 
.A(n_909),
.B(n_839),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_917),
.B(n_891),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_905),
.B(n_904),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_910),
.A2(n_898),
.B1(n_897),
.B2(n_714),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_905),
.B(n_903),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_907),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_910),
.Y(n_924)
);

NAND2x1p5_ASAP7_75t_L g925 ( 
.A(n_915),
.B(n_844),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_908),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_918),
.B(n_908),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_925),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_920),
.B(n_916),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_922),
.B(n_916),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_923),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_925),
.Y(n_932)
);

AND2x2_ASAP7_75t_SL g933 ( 
.A(n_919),
.B(n_914),
.Y(n_933)
);

AOI33xp33_ASAP7_75t_L g934 ( 
.A1(n_931),
.A2(n_924),
.A3(n_927),
.B1(n_932),
.B2(n_928),
.B3(n_929),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_928),
.B(n_924),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_929),
.B(n_930),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_933),
.A2(n_921),
.B1(n_900),
.B2(n_926),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_933),
.B(n_913),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_928),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_927),
.B(n_852),
.Y(n_940)
);

NAND2x1_ASAP7_75t_SL g941 ( 
.A(n_927),
.B(n_915),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_931),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_933),
.A2(n_900),
.B1(n_911),
.B2(n_912),
.Y(n_943)
);

HB1xp67_ASAP7_75t_L g944 ( 
.A(n_936),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_940),
.B(n_899),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_935),
.B(n_906),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_939),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_934),
.B(n_901),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_936),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_941),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_942),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_944),
.A2(n_943),
.B1(n_937),
.B2(n_938),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_946),
.Y(n_953)
);

AOI222xp33_ASAP7_75t_L g954 ( 
.A1(n_948),
.A2(n_912),
.B1(n_902),
.B2(n_869),
.C1(n_819),
.C2(n_747),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_949),
.B(n_906),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_949),
.A2(n_912),
.B1(n_870),
.B2(n_879),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_945),
.A2(n_867),
.B1(n_912),
.B2(n_892),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_950),
.A2(n_879),
.B1(n_895),
.B2(n_694),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_952),
.B(n_947),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_953),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_955),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_958),
.A2(n_951),
.B(n_954),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_956),
.Y(n_963)
);

INVxp67_ASAP7_75t_L g964 ( 
.A(n_959),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_960),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_961),
.B(n_957),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_963),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_962),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_960),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_967),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_969),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_L g972 ( 
.A(n_964),
.B(n_687),
.C(n_684),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_968),
.B(n_684),
.C(n_683),
.Y(n_973)
);

NOR3xp33_ASAP7_75t_L g974 ( 
.A(n_966),
.B(n_692),
.C(n_751),
.Y(n_974)
);

NOR2x1_ASAP7_75t_L g975 ( 
.A(n_965),
.B(n_778),
.Y(n_975)
);

AND3x4_ASAP7_75t_L g976 ( 
.A(n_974),
.B(n_692),
.C(n_774),
.Y(n_976)
);

AOI221xp5_ASAP7_75t_L g977 ( 
.A1(n_970),
.A2(n_778),
.B1(n_774),
.B2(n_702),
.C(n_867),
.Y(n_977)
);

O2A1O1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_971),
.A2(n_867),
.B(n_828),
.C(n_865),
.Y(n_978)
);

NAND4xp25_ASAP7_75t_SL g979 ( 
.A(n_972),
.B(n_866),
.C(n_704),
.D(n_878),
.Y(n_979)
);

NAND4xp75_ASAP7_75t_L g980 ( 
.A(n_975),
.B(n_704),
.C(n_798),
.D(n_878),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_977),
.B(n_973),
.Y(n_981)
);

OAI221xp5_ASAP7_75t_SL g982 ( 
.A1(n_978),
.A2(n_855),
.B1(n_863),
.B2(n_876),
.C(n_881),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_976),
.A2(n_874),
.B1(n_875),
.B2(n_881),
.Y(n_983)
);

OAI211xp5_ASAP7_75t_L g984 ( 
.A1(n_979),
.A2(n_699),
.B(n_806),
.C(n_784),
.Y(n_984)
);

AND2x4_ASAP7_75t_L g985 ( 
.A(n_980),
.B(n_875),
.Y(n_985)
);

HB1xp67_ASAP7_75t_L g986 ( 
.A(n_976),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_978),
.A2(n_766),
.B(n_768),
.C(n_876),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_976),
.B(n_699),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_986),
.B(n_877),
.Y(n_989)
);

NOR2x1_ASAP7_75t_L g990 ( 
.A(n_981),
.B(n_806),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_984),
.B(n_827),
.C(n_877),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_988),
.Y(n_992)
);

XNOR2xp5_ASAP7_75t_L g993 ( 
.A(n_985),
.B(n_142),
.Y(n_993)
);

AOI221xp5_ASAP7_75t_L g994 ( 
.A1(n_982),
.A2(n_812),
.B1(n_796),
.B2(n_886),
.C(n_793),
.Y(n_994)
);

INVx1_ASAP7_75t_SL g995 ( 
.A(n_983),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_987),
.B(n_886),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_985),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_990),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_997),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_995),
.B(n_797),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_993),
.A2(n_989),
.B1(n_992),
.B2(n_996),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_991),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_994),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_997),
.Y(n_1004)
);

NOR2x1_ASAP7_75t_L g1005 ( 
.A(n_993),
.B(n_806),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_990),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_990),
.Y(n_1007)
);

XNOR2xp5_ASAP7_75t_L g1008 ( 
.A(n_993),
.B(n_144),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_997),
.B(n_837),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_999),
.Y(n_1010)
);

INVxp33_ASAP7_75t_SL g1011 ( 
.A(n_1004),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_1001),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_998),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_1005),
.A2(n_806),
.B1(n_855),
.B2(n_863),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_1006),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1007),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_1003),
.B(n_863),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_1010),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1011),
.B(n_1002),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_1013),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_1013),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1017),
.Y(n_1022)
);

AOI21xp33_ASAP7_75t_L g1023 ( 
.A1(n_1015),
.A2(n_1012),
.B(n_1016),
.Y(n_1023)
);

OA21x2_ASAP7_75t_L g1024 ( 
.A1(n_1023),
.A2(n_1008),
.B(n_1000),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_R g1025 ( 
.A(n_1018),
.B(n_1009),
.Y(n_1025)
);

OR4x1_ASAP7_75t_L g1026 ( 
.A(n_1022),
.B(n_1014),
.C(n_146),
.D(n_147),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1026),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_1027),
.Y(n_1028)
);

AOI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_1028),
.A2(n_1019),
.B1(n_1020),
.B2(n_1021),
.Y(n_1029)
);

XNOR2xp5_ASAP7_75t_L g1030 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_1029),
.A2(n_1025),
.B(n_148),
.C(n_149),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_1030),
.A2(n_806),
.B1(n_855),
.B2(n_817),
.Y(n_1032)
);

AOI222xp33_ASAP7_75t_SL g1033 ( 
.A1(n_1031),
.A2(n_686),
.B1(n_150),
.B2(n_152),
.C1(n_153),
.C2(n_154),
.Y(n_1033)
);

AOI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1033),
.A2(n_686),
.B1(n_798),
.B2(n_827),
.Y(n_1034)
);

AOI222xp33_ASAP7_75t_L g1035 ( 
.A1(n_1032),
.A2(n_686),
.B1(n_157),
.B2(n_159),
.C1(n_166),
.C2(n_167),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_1035),
.A2(n_145),
.B(n_168),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_1036),
.A2(n_1034),
.B(n_171),
.Y(n_1037)
);

AOI211xp5_ASAP7_75t_L g1038 ( 
.A1(n_1037),
.A2(n_170),
.B(n_174),
.C(n_175),
.Y(n_1038)
);


endmodule