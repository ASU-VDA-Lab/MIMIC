module fake_ariane_2032_n_1242 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1242);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1242;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1218;
wire n_221;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_168;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_174;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

BUFx5_ASAP7_75t_L g166 ( 
.A(n_92),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_100),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_76),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_14),
.Y(n_171)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_71),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_161),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_23),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_64),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_126),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_55),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_106),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_26),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_79),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_138),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_97),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_95),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_139),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_60),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_90),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_44),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_142),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_14),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_74),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_133),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_77),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_131),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_12),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_101),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_52),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_163),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_34),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_32),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_25),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_109),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_80),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_152),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_140),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_56),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_38),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_87),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_43),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_151),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_20),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_75),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_59),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_122),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_10),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_112),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_10),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_156),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_53),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_50),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_123),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_118),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_19),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_147),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_46),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_73),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_159),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_125),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_135),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_32),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_148),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_144),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_134),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_16),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_43),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_113),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_103),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_18),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_1),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_132),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_81),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_136),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g273 ( 
.A(n_17),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_150),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_119),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_24),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_83),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_137),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_105),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_29),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_165),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_91),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_130),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_36),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_187),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_236),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g292 ( 
.A(n_195),
.B(n_0),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_187),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_236),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_173),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_173),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_171),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_195),
.B(n_2),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_211),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_266),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_185),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_176),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_167),
.B(n_2),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_192),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_215),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_171),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_217),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_218),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_175),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_171),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_175),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_232),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_171),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_171),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_171),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_238),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_220),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_202),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_220),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_252),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_226),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_172),
.B(n_3),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_265),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_273),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_199),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_227),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_273),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_269),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_210),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_273),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_228),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_231),
.B(n_3),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_177),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_242),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_181),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_227),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_248),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_243),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_182),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_268),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_239),
.B(n_4),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_281),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_282),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_243),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_226),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_186),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_226),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_209),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_208),
.B(n_5),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_189),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_207),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_170),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_193),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_170),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_194),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_179),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_179),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_169),
.B(n_6),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_174),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_178),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_197),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_207),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_208),
.Y(n_371)
);

BUFx6f_ASAP7_75t_SL g372 ( 
.A(n_199),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_183),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_184),
.B(n_6),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_204),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_188),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_297),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_297),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_366),
.B(n_204),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_306),
.Y(n_381)
);

NOR3xp33_ASAP7_75t_L g382 ( 
.A(n_347),
.B(n_200),
.C(n_198),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_203),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_219),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_244),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_310),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_319),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_316),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_327),
.B(n_221),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_168),
.Y(n_395)
);

BUFx2_ASAP7_75t_L g396 ( 
.A(n_287),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_233),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_351),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_369),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_240),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_353),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_319),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_376),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_365),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_377),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_328),
.B(n_246),
.Y(n_408)
);

INVx6_ASAP7_75t_L g409 ( 
.A(n_328),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_355),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_339),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_293),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_343),
.Y(n_415)
);

AND3x1_ASAP7_75t_L g416 ( 
.A(n_303),
.B(n_258),
.C(n_247),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_290),
.B(n_244),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_358),
.B(n_262),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_346),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_348),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_301),
.B(n_253),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_374),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_320),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_372),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_292),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_302),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_372),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_298),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_304),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_334),
.B(n_253),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_333),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_372),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_289),
.B(n_267),
.Y(n_435)
);

OAI22x1_ASAP7_75t_L g436 ( 
.A1(n_324),
.A2(n_271),
.B1(n_272),
.B2(n_275),
.Y(n_436)
);

AND2x4_ASAP7_75t_L g437 ( 
.A(n_363),
.B(n_364),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_299),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_338),
.B(n_267),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_340),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_352),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_359),
.B(n_213),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_361),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_409),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_416),
.A2(n_354),
.B1(n_322),
.B2(n_305),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_378),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_381),
.B(n_368),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_442),
.B(n_307),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_308),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g454 ( 
.A1(n_436),
.A2(n_375),
.B1(n_370),
.B2(n_357),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_378),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_442),
.B(n_312),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_381),
.B(n_166),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_378),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_168),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_441),
.B(n_317),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_436),
.A2(n_294),
.B1(n_291),
.B2(n_321),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_392),
.B(n_166),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_392),
.B(n_166),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_423),
.B(n_325),
.Y(n_468)
);

NAND3xp33_ASAP7_75t_L g469 ( 
.A(n_422),
.B(n_332),
.C(n_205),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_442),
.B(n_201),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_442),
.B(n_357),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_390),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_386),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_423),
.B(n_370),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_386),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_416),
.A2(n_354),
.B1(n_375),
.B2(n_250),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_394),
.B(n_166),
.Y(n_479)
);

OAI22xp33_ASAP7_75t_L g480 ( 
.A1(n_436),
.A2(n_300),
.B1(n_344),
.B2(n_341),
.Y(n_480)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_382),
.A2(n_256),
.B1(n_168),
.B2(n_190),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_382),
.A2(n_256),
.B1(n_168),
.B2(n_190),
.Y(n_482)
);

BUFx2_ASAP7_75t_L g483 ( 
.A(n_401),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_442),
.B(n_206),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_442),
.B(n_212),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_396),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_409),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g489 ( 
.A1(n_422),
.A2(n_256),
.B1(n_190),
.B2(n_214),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_391),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_409),
.Y(n_492)
);

INVx5_ASAP7_75t_L g493 ( 
.A(n_395),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_L g494 ( 
.A(n_442),
.B(n_216),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_386),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_423),
.B(n_295),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_SL g497 ( 
.A1(n_422),
.A2(n_309),
.B1(n_344),
.B2(n_341),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_401),
.B(n_295),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_394),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_380),
.B(n_296),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_406),
.B(n_166),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_406),
.B(n_166),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_379),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_400),
.A2(n_190),
.B1(n_256),
.B2(n_260),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_409),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_380),
.B(n_296),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_404),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_380),
.B(n_309),
.Y(n_509)
);

AO21x2_ASAP7_75t_L g510 ( 
.A1(n_393),
.A2(n_222),
.B(n_223),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_400),
.A2(n_270),
.B1(n_225),
.B2(n_229),
.Y(n_511)
);

NAND3xp33_ASAP7_75t_L g512 ( 
.A(n_406),
.B(n_224),
.C(n_230),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_379),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_379),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_425),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_400),
.A2(n_406),
.B1(n_407),
.B2(n_405),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_404),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_515),
.B(n_442),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_515),
.B(n_406),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_SL g522 ( 
.A(n_515),
.B(n_443),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_453),
.B(n_443),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_462),
.B(n_443),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_468),
.B(n_443),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_500),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_486),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_448),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_486),
.B(n_396),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_468),
.B(n_443),
.Y(n_530)
);

A2O1A1Ixp33_ASAP7_75t_L g531 ( 
.A1(n_500),
.A2(n_418),
.B(n_440),
.C(n_405),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_448),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_451),
.B(n_444),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_444),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_515),
.B(n_406),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_469),
.B(n_406),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_455),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_469),
.A2(n_444),
.B1(n_440),
.B2(n_447),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_444),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_455),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_514),
.B(n_406),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_508),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_458),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_483),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_452),
.B(n_444),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_508),
.B(n_447),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_483),
.B(n_396),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_518),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_458),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_471),
.B(n_447),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_518),
.B(n_439),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_502),
.A2(n_503),
.B(n_499),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_460),
.B(n_439),
.Y(n_553)
);

BUFx3_ASAP7_75t_L g554 ( 
.A(n_448),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_475),
.B(n_427),
.Y(n_555)
);

BUFx6f_ASAP7_75t_SL g556 ( 
.A(n_461),
.Y(n_556)
);

AOI221xp5_ASAP7_75t_L g557 ( 
.A1(n_449),
.A2(n_433),
.B1(n_418),
.B2(n_419),
.C(n_415),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_460),
.B(n_439),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_449),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_514),
.B(n_446),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_464),
.B(n_446),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_482),
.B1(n_464),
.B2(n_474),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_467),
.B(n_445),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_467),
.B(n_445),
.Y(n_565)
);

O2A1O1Ixp33_ASAP7_75t_L g566 ( 
.A1(n_456),
.A2(n_383),
.B(n_419),
.C(n_415),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_498),
.B(n_438),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_514),
.B(n_427),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_475),
.B(n_429),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_474),
.B(n_400),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_476),
.B(n_383),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_476),
.B(n_421),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_487),
.B(n_421),
.Y(n_573)
);

INVx1_ASAP7_75t_SL g574 ( 
.A(n_498),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_487),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_459),
.Y(n_576)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_431),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_501),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

O2A1O1Ixp33_ASAP7_75t_L g580 ( 
.A1(n_457),
.A2(n_420),
.B(n_412),
.C(n_398),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g581 ( 
.A(n_496),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_450),
.B(n_421),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_510),
.B(n_429),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_514),
.B(n_431),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_510),
.A2(n_437),
.B1(n_433),
.B2(n_429),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_450),
.B(n_428),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_472),
.B(n_428),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_497),
.A2(n_318),
.B1(n_311),
.B2(n_329),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_488),
.Y(n_590)
);

NAND2xp33_ASAP7_75t_L g591 ( 
.A(n_514),
.B(n_386),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_472),
.B(n_428),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_SL g594 ( 
.A(n_473),
.B(n_425),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_514),
.B(n_386),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_473),
.B(n_386),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_490),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_490),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_510),
.B(n_429),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_432),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_473),
.B(n_386),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_496),
.B(n_432),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_501),
.B(n_437),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_473),
.B(n_386),
.Y(n_604)
);

NOR2xp67_ASAP7_75t_L g605 ( 
.A(n_478),
.B(n_425),
.Y(n_605)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_510),
.A2(n_437),
.B1(n_409),
.B2(n_411),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_507),
.B(n_432),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_457),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_502),
.A2(n_398),
.B(n_393),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_477),
.B(n_389),
.Y(n_611)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_507),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_477),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_477),
.Y(n_615)
);

BUFx5_ASAP7_75t_L g616 ( 
.A(n_488),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_466),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_552),
.A2(n_503),
.B(n_499),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_526),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_520),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_525),
.B(n_417),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_541),
.A2(n_499),
.B(n_491),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_530),
.B(n_417),
.Y(n_623)
);

AOI21x1_ASAP7_75t_L g624 ( 
.A1(n_519),
.A2(n_479),
.B(n_466),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_523),
.B(n_417),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_524),
.B(n_509),
.Y(n_626)
);

AOI21xp5_ASAP7_75t_L g627 ( 
.A1(n_541),
.A2(n_504),
.B(n_491),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_554),
.Y(n_628)
);

BUFx8_ASAP7_75t_SL g629 ( 
.A(n_544),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_527),
.B(n_311),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_542),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_529),
.B(n_509),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_533),
.B(n_480),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_569),
.B(n_437),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_556),
.Y(n_635)
);

NOR2x1_ASAP7_75t_R g636 ( 
.A(n_559),
.B(n_437),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_521),
.A2(n_504),
.B(n_491),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_548),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_554),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g640 ( 
.A1(n_521),
.A2(n_513),
.B(n_504),
.Y(n_640)
);

BUFx2_ASAP7_75t_SL g641 ( 
.A(n_556),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_535),
.A2(n_534),
.B(n_519),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_536),
.A2(n_484),
.B(n_485),
.C(n_479),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_569),
.B(n_413),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_535),
.A2(n_517),
.B(n_513),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_578),
.Y(n_647)
);

OAI21xp33_ASAP7_75t_L g648 ( 
.A1(n_551),
.A2(n_511),
.B(n_454),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_547),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_574),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_555),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_610),
.A2(n_517),
.B(n_513),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_528),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_602),
.B(n_407),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_594),
.A2(n_517),
.B(n_512),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_550),
.A2(n_318),
.B1(n_329),
.B2(n_321),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_538),
.B(n_411),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_528),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_575),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_563),
.A2(n_495),
.B(n_477),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_565),
.B(n_413),
.Y(n_661)
);

INVx11_ASAP7_75t_L g662 ( 
.A(n_612),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_581),
.B(n_412),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_567),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_600),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_607),
.B(n_497),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_550),
.B(n_413),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_531),
.B(n_413),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_528),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_532),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_612),
.B(n_435),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_577),
.A2(n_350),
.B1(n_409),
.B2(n_461),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_603),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_531),
.B(n_385),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_537),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_540),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_581),
.B(n_350),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_583),
.A2(n_495),
.B(n_512),
.C(n_463),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_603),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_543),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_549),
.Y(n_683)
);

AO21x1_ASAP7_75t_L g684 ( 
.A1(n_536),
.A2(n_494),
.B(n_470),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_553),
.B(n_385),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_557),
.B(n_435),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_605),
.B(n_420),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_587),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_558),
.B(n_385),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_595),
.A2(n_495),
.B(n_506),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_598),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_595),
.A2(n_495),
.B(n_506),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_571),
.B(n_561),
.Y(n_693)
);

NOR2x1_ASAP7_75t_R g694 ( 
.A(n_568),
.B(n_291),
.Y(n_694)
);

BUFx6f_ASAP7_75t_L g695 ( 
.A(n_532),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_568),
.A2(n_461),
.B1(n_489),
.B2(n_424),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g697 ( 
.A1(n_608),
.A2(n_614),
.B(n_609),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_585),
.B(n_435),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_617),
.A2(n_506),
.B(n_389),
.Y(n_699)
);

NOR2xp67_ASAP7_75t_L g700 ( 
.A(n_545),
.B(n_408),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_572),
.A2(n_402),
.B(n_414),
.C(n_410),
.Y(n_701)
);

OAI21xp33_ASAP7_75t_L g702 ( 
.A1(n_546),
.A2(n_424),
.B(n_402),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_584),
.B(n_294),
.Y(n_703)
);

AND2x6_ASAP7_75t_SL g704 ( 
.A(n_583),
.B(n_426),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_596),
.A2(n_611),
.B(n_601),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_573),
.B(n_408),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_582),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_584),
.B(n_384),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_596),
.A2(n_389),
.B(n_488),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_539),
.B(n_599),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_576),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_599),
.B(n_384),
.Y(n_712)
);

OAI21xp5_ASAP7_75t_L g713 ( 
.A1(n_601),
.A2(n_492),
.B(n_505),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_562),
.B(n_461),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_611),
.A2(n_389),
.B(n_492),
.Y(n_715)
);

O2A1O1Ixp5_ASAP7_75t_L g716 ( 
.A1(n_684),
.A2(n_560),
.B(n_522),
.C(n_570),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_642),
.A2(n_580),
.B(n_566),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_653),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_693),
.A2(n_591),
.B(n_604),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_667),
.A2(n_589),
.B1(n_463),
.B2(n_426),
.Y(n_720)
);

OAI21xp5_ASAP7_75t_L g721 ( 
.A1(n_642),
.A2(n_606),
.B(n_560),
.Y(n_721)
);

INVx4_ASAP7_75t_L g722 ( 
.A(n_629),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_707),
.B(n_579),
.Y(n_723)
);

BUFx12f_ASAP7_75t_L g724 ( 
.A(n_635),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_651),
.B(n_430),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_712),
.B(n_593),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_679),
.A2(n_664),
.B1(n_649),
.B2(n_703),
.Y(n_727)
);

CKINVDCx20_ASAP7_75t_R g728 ( 
.A(n_650),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_630),
.B(n_613),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_SL g730 ( 
.A1(n_656),
.A2(n_430),
.B1(n_461),
.B2(n_562),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_626),
.A2(n_410),
.B(n_414),
.C(n_615),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_695),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_651),
.B(n_686),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_649),
.A2(n_532),
.B1(n_590),
.B2(n_616),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_632),
.B(n_410),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_653),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_620),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_619),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_695),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_676),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_666),
.B(n_597),
.Y(n_741)
);

O2A1O1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_634),
.A2(n_414),
.B(n_586),
.C(n_588),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_695),
.Y(n_743)
);

BUFx6f_ASAP7_75t_L g744 ( 
.A(n_658),
.Y(n_744)
);

BUFx6f_ASAP7_75t_SL g745 ( 
.A(n_647),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_662),
.B(n_592),
.Y(n_746)
);

BUFx2_ASAP7_75t_L g747 ( 
.A(n_694),
.Y(n_747)
);

O2A1O1Ixp33_ASAP7_75t_L g748 ( 
.A1(n_625),
.A2(n_689),
.B(n_685),
.C(n_633),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_697),
.A2(n_590),
.B(n_564),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_636),
.B(n_590),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_654),
.B(n_590),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_672),
.B(n_425),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_706),
.B(n_616),
.Y(n_753)
);

BUFx2_ASAP7_75t_L g754 ( 
.A(n_654),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_SL g755 ( 
.A1(n_674),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_698),
.B(n_616),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_644),
.A2(n_492),
.B(n_434),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_652),
.A2(n_434),
.B(n_425),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_641),
.Y(n_759)
);

OAI21xp33_ASAP7_75t_SL g760 ( 
.A1(n_631),
.A2(n_616),
.B(n_403),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_663),
.B(n_387),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_635),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_638),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_710),
.B(n_616),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_658),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_674),
.B(n_389),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_628),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_SL g768 ( 
.A(n_648),
.B(n_241),
.C(n_245),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_652),
.A2(n_434),
.B(n_616),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_663),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_675),
.A2(n_397),
.B1(n_387),
.B2(n_399),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_680),
.B(n_681),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_704),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_678),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_665),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_687),
.Y(n_776)
);

OAI21x1_ASAP7_75t_L g777 ( 
.A1(n_618),
.A2(n_403),
.B(n_399),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_622),
.A2(n_434),
.B(n_389),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_621),
.B(n_434),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_681),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_659),
.Y(n_781)
);

OAI22x1_ASAP7_75t_L g782 ( 
.A1(n_673),
.A2(n_249),
.B1(n_251),
.B2(n_254),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_623),
.B(n_387),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_687),
.B(n_389),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_770),
.B(n_708),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_776),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_730),
.A2(n_727),
.B1(n_772),
.B2(n_733),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_738),
.Y(n_788)
);

OAI21xp5_ASAP7_75t_L g789 ( 
.A1(n_764),
.A2(n_705),
.B(n_643),
.Y(n_789)
);

AO31x2_ASAP7_75t_L g790 ( 
.A1(n_764),
.A2(n_714),
.A3(n_699),
.B(n_669),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_772),
.A2(n_702),
.B1(n_657),
.B2(n_696),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_753),
.A2(n_699),
.B(n_701),
.Y(n_792)
);

INVx2_ASAP7_75t_R g793 ( 
.A(n_763),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_754),
.A2(n_661),
.B1(n_700),
.B2(n_639),
.Y(n_794)
);

AO31x2_ASAP7_75t_L g795 ( 
.A1(n_726),
.A2(n_622),
.A3(n_627),
.B(n_637),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_753),
.A2(n_719),
.B(n_769),
.Y(n_796)
);

AOI211x1_ASAP7_75t_L g797 ( 
.A1(n_781),
.A2(n_705),
.B(n_660),
.C(n_688),
.Y(n_797)
);

OAI22xp33_ASAP7_75t_L g798 ( 
.A1(n_773),
.A2(n_668),
.B1(n_691),
.B2(n_639),
.Y(n_798)
);

NAND3xp33_ASAP7_75t_SL g799 ( 
.A(n_746),
.B(n_701),
.C(n_259),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_717),
.A2(n_627),
.B(n_646),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_724),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_728),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_729),
.B(n_711),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_734),
.B(n_748),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_744),
.Y(n_805)
);

OAI21xp5_ASAP7_75t_L g806 ( 
.A1(n_716),
.A2(n_643),
.B(n_660),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_SL g807 ( 
.A1(n_782),
.A2(n_677),
.B1(n_671),
.B2(n_670),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_717),
.A2(n_637),
.B(n_640),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_756),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_721),
.A2(n_640),
.B(n_646),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_737),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_751),
.A2(n_725),
.B(n_721),
.C(n_768),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_735),
.B(n_682),
.Y(n_814)
);

BUFx12f_ASAP7_75t_L g815 ( 
.A(n_722),
.Y(n_815)
);

OAI21x1_ASAP7_75t_L g816 ( 
.A1(n_777),
.A2(n_655),
.B(n_624),
.Y(n_816)
);

OAI21x1_ASAP7_75t_L g817 ( 
.A1(n_778),
.A2(n_692),
.B(n_690),
.Y(n_817)
);

OA21x2_ASAP7_75t_L g818 ( 
.A1(n_758),
.A2(n_692),
.B(n_690),
.Y(n_818)
);

O2A1O1Ixp5_ASAP7_75t_L g819 ( 
.A1(n_771),
.A2(n_670),
.B(n_645),
.C(n_671),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_756),
.A2(n_628),
.B1(n_645),
.B2(n_677),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_744),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_761),
.B(n_387),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_742),
.A2(n_709),
.B(n_715),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_745),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_726),
.A2(n_709),
.B(n_715),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_740),
.Y(n_826)
);

NAND3x1_ASAP7_75t_L g827 ( 
.A(n_750),
.B(n_397),
.C(n_387),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_SL g828 ( 
.A1(n_752),
.A2(n_713),
.B(n_683),
.C(n_397),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_731),
.A2(n_397),
.B(n_280),
.C(n_279),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_720),
.B(n_397),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_775),
.B(n_7),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_780),
.B(n_7),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_749),
.A2(n_379),
.B(n_389),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_774),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_784),
.A2(n_395),
.B1(n_283),
.B2(n_278),
.Y(n_835)
);

OAI21x1_ASAP7_75t_L g836 ( 
.A1(n_757),
.A2(n_379),
.B(n_47),
.Y(n_836)
);

O2A1O1Ixp33_ASAP7_75t_L g837 ( 
.A1(n_783),
.A2(n_8),
.B(n_9),
.C(n_11),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_747),
.B(n_8),
.Y(n_838)
);

AO31x2_ASAP7_75t_L g839 ( 
.A1(n_771),
.A2(n_395),
.A3(n_493),
.B(n_94),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_766),
.A2(n_285),
.B(n_284),
.C(n_277),
.Y(n_840)
);

NAND3xp33_ASAP7_75t_SL g841 ( 
.A(n_759),
.B(n_255),
.C(n_263),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_760),
.A2(n_493),
.B(n_274),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_787),
.A2(n_723),
.B1(n_741),
.B2(n_755),
.Y(n_843)
);

BUFx3_ASAP7_75t_L g844 ( 
.A(n_786),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_803),
.B(n_723),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_788),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_807),
.A2(n_745),
.B1(n_741),
.B2(n_762),
.Y(n_847)
);

CKINVDCx20_ASAP7_75t_R g848 ( 
.A(n_824),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_826),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_805),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_811),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_834),
.Y(n_852)
);

INVx4_ASAP7_75t_L g853 ( 
.A(n_805),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_814),
.Y(n_854)
);

CKINVDCx6p67_ASAP7_75t_R g855 ( 
.A(n_815),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_SL g856 ( 
.A1(n_787),
.A2(n_718),
.B(n_736),
.Y(n_856)
);

CKINVDCx11_ASAP7_75t_R g857 ( 
.A(n_802),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_797),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_822),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_786),
.Y(n_860)
);

INVx8_ASAP7_75t_L g861 ( 
.A(n_805),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_791),
.A2(n_767),
.B1(n_722),
.B2(n_718),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_801),
.Y(n_863)
);

CKINVDCx11_ASAP7_75t_R g864 ( 
.A(n_786),
.Y(n_864)
);

INVx6_ASAP7_75t_L g865 ( 
.A(n_821),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_785),
.Y(n_866)
);

CKINVDCx11_ASAP7_75t_R g867 ( 
.A(n_821),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_797),
.Y(n_868)
);

CKINVDCx20_ASAP7_75t_R g869 ( 
.A(n_838),
.Y(n_869)
);

CKINVDCx11_ASAP7_75t_R g870 ( 
.A(n_821),
.Y(n_870)
);

INVx1_ASAP7_75t_SL g871 ( 
.A(n_832),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_812),
.Y(n_872)
);

INVx6_ASAP7_75t_L g873 ( 
.A(n_831),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_791),
.A2(n_779),
.B1(n_736),
.B2(n_744),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_809),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_798),
.A2(n_765),
.B1(n_779),
.B2(n_743),
.Y(n_876)
);

CKINVDCx16_ASAP7_75t_R g877 ( 
.A(n_841),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_830),
.A2(n_765),
.B1(n_743),
.B2(n_739),
.Y(n_878)
);

OAI21xp33_ASAP7_75t_SL g879 ( 
.A1(n_804),
.A2(n_789),
.B(n_806),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_790),
.Y(n_880)
);

INVx3_ASAP7_75t_SL g881 ( 
.A(n_812),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_SL g882 ( 
.A1(n_794),
.A2(n_765),
.B1(n_743),
.B2(n_739),
.Y(n_882)
);

OAI22xp33_ASAP7_75t_L g883 ( 
.A1(n_799),
.A2(n_739),
.B1(n_732),
.B2(n_13),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_793),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_790),
.Y(n_885)
);

CKINVDCx11_ASAP7_75t_R g886 ( 
.A(n_820),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_840),
.A2(n_732),
.B1(n_11),
.B2(n_15),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_827),
.A2(n_9),
.B1(n_15),
.B2(n_16),
.Y(n_888)
);

INVx1_ASAP7_75t_SL g889 ( 
.A(n_807),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_790),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_835),
.Y(n_891)
);

BUFx2_ASAP7_75t_SL g892 ( 
.A(n_808),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_795),
.Y(n_893)
);

CKINVDCx11_ASAP7_75t_R g894 ( 
.A(n_837),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_835),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_817),
.Y(n_896)
);

CKINVDCx6p67_ASAP7_75t_R g897 ( 
.A(n_813),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_796),
.A2(n_493),
.B(n_18),
.Y(n_898)
);

OAI21xp33_ASAP7_75t_L g899 ( 
.A1(n_800),
.A2(n_17),
.B(n_20),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_839),
.B(n_21),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_842),
.Y(n_901)
);

BUFx12f_ASAP7_75t_L g902 ( 
.A(n_819),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_839),
.B(n_21),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_858),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_875),
.B(n_810),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_880),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_868),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_885),
.Y(n_908)
);

INVx4_ASAP7_75t_L g909 ( 
.A(n_902),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_893),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_897),
.B(n_894),
.Y(n_911)
);

OR2x2_ASAP7_75t_L g912 ( 
.A(n_885),
.B(n_795),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_880),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_893),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_890),
.Y(n_915)
);

INVx1_ASAP7_75t_SL g916 ( 
.A(n_889),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_884),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_863),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_846),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_896),
.Y(n_920)
);

OAI21x1_ASAP7_75t_L g921 ( 
.A1(n_898),
.A2(n_823),
.B(n_816),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_852),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_892),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_845),
.B(n_792),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_896),
.Y(n_925)
);

OR2x2_ASAP7_75t_L g926 ( 
.A(n_859),
.B(n_795),
.Y(n_926)
);

OAI21x1_ASAP7_75t_L g927 ( 
.A1(n_874),
.A2(n_825),
.B(n_833),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_896),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_896),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_851),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_849),
.Y(n_931)
);

OAI21xp5_ASAP7_75t_L g932 ( 
.A1(n_879),
.A2(n_829),
.B(n_828),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_900),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_903),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_894),
.A2(n_818),
.B1(n_839),
.B2(n_836),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_899),
.A2(n_818),
.B(n_395),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_873),
.B(n_22),
.Y(n_937)
);

OAI21x1_ASAP7_75t_L g938 ( 
.A1(n_878),
.A2(n_395),
.B(n_98),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_872),
.Y(n_939)
);

INVx4_ASAP7_75t_SL g940 ( 
.A(n_882),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_866),
.Y(n_941)
);

AOI221xp5_ASAP7_75t_L g942 ( 
.A1(n_911),
.A2(n_933),
.B1(n_843),
.B2(n_883),
.C(n_891),
.Y(n_942)
);

AND2x4_ASAP7_75t_L g943 ( 
.A(n_923),
.B(n_844),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_934),
.B(n_873),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_934),
.B(n_873),
.Y(n_945)
);

OAI22xp33_ASAP7_75t_L g946 ( 
.A1(n_911),
.A2(n_883),
.B1(n_895),
.B2(n_862),
.Y(n_946)
);

INVx4_ASAP7_75t_L g947 ( 
.A(n_940),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_934),
.B(n_871),
.Y(n_948)
);

AOI221xp5_ASAP7_75t_L g949 ( 
.A1(n_933),
.A2(n_843),
.B1(n_887),
.B2(n_888),
.C(n_877),
.Y(n_949)
);

OR2x6_ASAP7_75t_L g950 ( 
.A(n_934),
.B(n_856),
.Y(n_950)
);

AOI21xp33_ASAP7_75t_L g951 ( 
.A1(n_923),
.A2(n_847),
.B(n_901),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_919),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_926),
.B(n_844),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_919),
.B(n_886),
.Y(n_954)
);

BUFx3_ASAP7_75t_L g955 ( 
.A(n_937),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_916),
.A2(n_869),
.B1(n_886),
.B2(n_940),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_935),
.A2(n_878),
.B(n_876),
.Y(n_957)
);

HB1xp67_ASAP7_75t_L g958 ( 
.A(n_917),
.Y(n_958)
);

AOI22xp5_ASAP7_75t_L g959 ( 
.A1(n_916),
.A2(n_864),
.B1(n_870),
.B2(n_867),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_922),
.B(n_854),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_940),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_926),
.B(n_860),
.Y(n_962)
);

OAI21x1_ASAP7_75t_L g963 ( 
.A1(n_921),
.A2(n_850),
.B(n_881),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_937),
.A2(n_881),
.B1(n_855),
.B2(n_865),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_931),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_932),
.A2(n_850),
.B(n_853),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_929),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_922),
.B(n_860),
.Y(n_968)
);

INVxp67_ASAP7_75t_L g969 ( 
.A(n_939),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_917),
.B(n_872),
.Y(n_970)
);

AO21x2_ASAP7_75t_L g971 ( 
.A1(n_936),
.A2(n_872),
.B(n_865),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_924),
.B(n_937),
.Y(n_972)
);

NOR2x1_ASAP7_75t_SL g973 ( 
.A(n_909),
.B(n_872),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_932),
.A2(n_935),
.B(n_924),
.Y(n_974)
);

BUFx10_ASAP7_75t_L g975 ( 
.A(n_939),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_918),
.B(n_857),
.Y(n_976)
);

AOI22xp33_ASAP7_75t_L g977 ( 
.A1(n_909),
.A2(n_864),
.B1(n_857),
.B2(n_870),
.Y(n_977)
);

BUFx3_ASAP7_75t_L g978 ( 
.A(n_930),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_929),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_SL g980 ( 
.A1(n_909),
.A2(n_853),
.B(n_867),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_926),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_963),
.Y(n_982)
);

INVx2_ASAP7_75t_SL g983 ( 
.A(n_975),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_978),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_958),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_978),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_944),
.B(n_920),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_972),
.B(n_912),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_944),
.B(n_920),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_965),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_947),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_952),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_965),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_952),
.Y(n_994)
);

OR2x2_ASAP7_75t_L g995 ( 
.A(n_981),
.B(n_912),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_945),
.B(n_920),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_969),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_963),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_946),
.A2(n_909),
.B1(n_940),
.B2(n_936),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_960),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_981),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_971),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_974),
.B(n_905),
.C(n_904),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_948),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_942),
.A2(n_949),
.B1(n_956),
.B2(n_954),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_976),
.B(n_918),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_945),
.B(n_920),
.Y(n_1007)
);

OAI221xp5_ASAP7_75t_SL g1008 ( 
.A1(n_1005),
.A2(n_956),
.B1(n_959),
.B2(n_950),
.C(n_977),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_990),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_992),
.Y(n_1010)
);

NOR2x1_ASAP7_75t_R g1011 ( 
.A(n_991),
.B(n_947),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_985),
.B(n_970),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_992),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_985),
.B(n_970),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_997),
.Y(n_1015)
);

AOI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_1005),
.A2(n_909),
.B1(n_957),
.B2(n_951),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_997),
.B(n_954),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_987),
.B(n_943),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_987),
.B(n_950),
.Y(n_1019)
);

OR2x2_ASAP7_75t_SL g1020 ( 
.A(n_1003),
.B(n_968),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_994),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_994),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_987),
.B(n_943),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_988),
.B(n_1000),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_989),
.B(n_943),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_995),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_989),
.B(n_943),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_988),
.B(n_905),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_989),
.B(n_967),
.Y(n_1029)
);

INVxp67_ASAP7_75t_L g1030 ( 
.A(n_1017),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_1015),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1028),
.B(n_1003),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_1019),
.B(n_991),
.Y(n_1033)
);

OR2x2_ASAP7_75t_L g1034 ( 
.A(n_1028),
.B(n_988),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1036)
);

AND2x4_ASAP7_75t_SL g1037 ( 
.A(n_1017),
.B(n_991),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1010),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_991),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1023),
.B(n_1001),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1023),
.B(n_1001),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1033),
.B(n_1025),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1033),
.B(n_1025),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1038),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1038),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_1033),
.B(n_1027),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1034),
.B(n_1020),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1032),
.B(n_1015),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1035),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1047),
.B(n_1030),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1048),
.B(n_1020),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1049),
.B(n_1034),
.Y(n_1052)
);

NAND4xp25_ASAP7_75t_L g1053 ( 
.A(n_1044),
.B(n_1031),
.C(n_1008),
.D(n_1006),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1052),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1050),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_1051),
.B(n_1042),
.Y(n_1056)
);

INVxp67_ASAP7_75t_L g1057 ( 
.A(n_1053),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1052),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_1051),
.B(n_1049),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_1051),
.B(n_1042),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_1051),
.B(n_1043),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1052),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_1051),
.A2(n_1016),
.B1(n_999),
.B2(n_959),
.Y(n_1063)
);

AOI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1051),
.A2(n_1016),
.B1(n_999),
.B2(n_957),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1060),
.B(n_1043),
.Y(n_1065)
);

OAI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1064),
.A2(n_1008),
.B1(n_1045),
.B2(n_1031),
.C(n_1024),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1055),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_1056),
.B(n_1033),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1063),
.A2(n_1046),
.B1(n_1039),
.B2(n_1037),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1057),
.B(n_1031),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_1054),
.B(n_1031),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1064),
.A2(n_1046),
.B1(n_1039),
.B2(n_1037),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1058),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_1062),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1059),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1061),
.B(n_1035),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1056),
.A2(n_848),
.B(n_980),
.Y(n_1077)
);

AOI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_1064),
.A2(n_1019),
.B1(n_948),
.B2(n_964),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1055),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1063),
.A2(n_1039),
.B1(n_1026),
.B2(n_1024),
.Y(n_1080)
);

OAI21xp33_ASAP7_75t_L g1081 ( 
.A1(n_1070),
.A2(n_1065),
.B(n_1075),
.Y(n_1081)
);

AOI22xp5_ASAP7_75t_L g1082 ( 
.A1(n_1066),
.A2(n_1039),
.B1(n_982),
.B2(n_998),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1067),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1079),
.Y(n_1084)
);

INVx1_ASAP7_75t_SL g1085 ( 
.A(n_1073),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_1078),
.A2(n_957),
.B1(n_950),
.B2(n_947),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1074),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1076),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1068),
.B(n_1040),
.Y(n_1089)
);

INVx1_ASAP7_75t_SL g1090 ( 
.A(n_1071),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1077),
.A2(n_961),
.B1(n_1026),
.B2(n_1041),
.Y(n_1091)
);

AO21x1_ASAP7_75t_L g1092 ( 
.A1(n_1072),
.A2(n_1041),
.B(n_1040),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1080),
.A2(n_998),
.B(n_982),
.C(n_950),
.Y(n_1093)
);

AOI221xp5_ASAP7_75t_L g1094 ( 
.A1(n_1069),
.A2(n_982),
.B1(n_998),
.B2(n_1000),
.C(n_1022),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1077),
.Y(n_1095)
);

OR2x2_ASAP7_75t_L g1096 ( 
.A(n_1076),
.B(n_1036),
.Y(n_1096)
);

OAI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_1066),
.A2(n_980),
.B1(n_982),
.B2(n_998),
.C(n_966),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_1075),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1067),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1096),
.Y(n_1100)
);

AOI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_1085),
.A2(n_1002),
.B(n_1009),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1098),
.Y(n_1102)
);

INVx1_ASAP7_75t_SL g1103 ( 
.A(n_1090),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1099),
.B(n_1013),
.C(n_1010),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_1085),
.B(n_1013),
.Y(n_1105)
);

NOR3x1_ASAP7_75t_L g1106 ( 
.A(n_1095),
.B(n_983),
.C(n_1021),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1090),
.B(n_1088),
.Y(n_1107)
);

AND2x2_ASAP7_75t_L g1108 ( 
.A(n_1089),
.B(n_1036),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1081),
.B(n_1012),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1083),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1084),
.B(n_1012),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1087),
.Y(n_1112)
);

AOI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1091),
.A2(n_1014),
.B1(n_983),
.B2(n_1022),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1092),
.Y(n_1114)
);

AND5x1_ASAP7_75t_L g1115 ( 
.A(n_1082),
.B(n_1011),
.C(n_961),
.D(n_940),
.E(n_973),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1094),
.B(n_1086),
.Y(n_1116)
);

OAI21xp33_ASAP7_75t_SL g1117 ( 
.A1(n_1114),
.A2(n_1097),
.B(n_1093),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1103),
.B(n_1014),
.Y(n_1118)
);

AOI211x1_ASAP7_75t_SL g1119 ( 
.A1(n_1107),
.A2(n_1105),
.B(n_1116),
.C(n_1104),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1102),
.B(n_1021),
.Y(n_1120)
);

BUFx8_ASAP7_75t_L g1121 ( 
.A(n_1112),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1111),
.A2(n_1009),
.B1(n_957),
.B2(n_961),
.Y(n_1122)
);

OAI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1100),
.A2(n_983),
.B(n_861),
.C(n_1029),
.Y(n_1123)
);

OAI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1112),
.A2(n_1009),
.B1(n_986),
.B2(n_984),
.Y(n_1124)
);

NOR3xp33_ASAP7_75t_L g1125 ( 
.A(n_1110),
.B(n_1011),
.C(n_938),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_L g1126 ( 
.A(n_1105),
.B(n_904),
.C(n_907),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1101),
.A2(n_938),
.B(n_1027),
.C(n_1002),
.Y(n_1127)
);

AOI221xp5_ASAP7_75t_L g1128 ( 
.A1(n_1111),
.A2(n_941),
.B1(n_1002),
.B2(n_936),
.C(n_907),
.Y(n_1128)
);

AOI311xp33_ASAP7_75t_L g1129 ( 
.A1(n_1106),
.A2(n_22),
.A3(n_23),
.B(n_25),
.C(n_26),
.Y(n_1129)
);

AOI211xp5_ASAP7_75t_L g1130 ( 
.A1(n_1109),
.A2(n_27),
.B(n_28),
.C(n_29),
.Y(n_1130)
);

INVx1_ASAP7_75t_SL g1131 ( 
.A(n_1108),
.Y(n_1131)
);

AND4x1_ASAP7_75t_L g1132 ( 
.A(n_1108),
.B(n_27),
.C(n_28),
.D(n_30),
.Y(n_1132)
);

AOI211xp5_ASAP7_75t_L g1133 ( 
.A1(n_1115),
.A2(n_30),
.B(n_31),
.C(n_33),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1113),
.A2(n_1029),
.B(n_861),
.Y(n_1134)
);

NAND4xp25_ASAP7_75t_L g1135 ( 
.A(n_1102),
.B(n_967),
.C(n_979),
.D(n_955),
.Y(n_1135)
);

NAND2x1_ASAP7_75t_L g1136 ( 
.A(n_1102),
.B(n_865),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1103),
.B(n_1007),
.Y(n_1137)
);

NOR4xp25_ASAP7_75t_L g1138 ( 
.A(n_1103),
.B(n_31),
.C(n_33),
.D(n_34),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1102),
.B(n_996),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1103),
.B(n_996),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1138),
.B(n_984),
.Y(n_1141)
);

AOI211xp5_ASAP7_75t_L g1142 ( 
.A1(n_1117),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1131),
.A2(n_1118),
.B1(n_1140),
.B2(n_1137),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1121),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_1121),
.Y(n_1145)
);

AOI221xp5_ASAP7_75t_L g1146 ( 
.A1(n_1125),
.A2(n_941),
.B1(n_936),
.B2(n_986),
.C(n_984),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1130),
.A2(n_986),
.B1(n_967),
.B2(n_979),
.Y(n_1147)
);

AOI221xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1120),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.C(n_39),
.Y(n_1148)
);

AOI211xp5_ASAP7_75t_L g1149 ( 
.A1(n_1119),
.A2(n_39),
.B(n_40),
.C(n_41),
.Y(n_1149)
);

XOR2x2_ASAP7_75t_L g1150 ( 
.A(n_1132),
.B(n_1133),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1123),
.A2(n_40),
.B(n_41),
.C(n_42),
.Y(n_1151)
);

AOI221x1_ASAP7_75t_L g1152 ( 
.A1(n_1135),
.A2(n_42),
.B1(n_908),
.B2(n_979),
.C(n_1007),
.Y(n_1152)
);

AOI221xp5_ASAP7_75t_L g1153 ( 
.A1(n_1127),
.A2(n_936),
.B1(n_928),
.B2(n_908),
.C(n_1007),
.Y(n_1153)
);

AOI211xp5_ASAP7_75t_L g1154 ( 
.A1(n_1139),
.A2(n_938),
.B(n_995),
.C(n_928),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1136),
.B(n_996),
.Y(n_1155)
);

AOI21xp33_ASAP7_75t_L g1156 ( 
.A1(n_1124),
.A2(n_861),
.B(n_993),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1126),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1134),
.A2(n_995),
.B(n_925),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1122),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1129),
.Y(n_1160)
);

BUFx2_ASAP7_75t_L g1161 ( 
.A(n_1128),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1121),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1125),
.A2(n_940),
.B1(n_962),
.B2(n_953),
.Y(n_1163)
);

NAND4xp25_ASAP7_75t_L g1164 ( 
.A(n_1119),
.B(n_955),
.C(n_929),
.D(n_928),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1150),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1145),
.Y(n_1166)
);

NOR2x1_ASAP7_75t_L g1167 ( 
.A(n_1144),
.B(n_929),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1141),
.Y(n_1168)
);

NAND3xp33_ASAP7_75t_L g1169 ( 
.A(n_1149),
.B(n_493),
.C(n_912),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1162),
.B(n_975),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1149),
.B(n_953),
.Y(n_1171)
);

OR2x2_ASAP7_75t_L g1172 ( 
.A(n_1160),
.B(n_990),
.Y(n_1172)
);

NOR2x1_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_929),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1143),
.B(n_975),
.Y(n_1174)
);

XOR2x1_ASAP7_75t_L g1175 ( 
.A(n_1157),
.B(n_953),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1152),
.B(n_973),
.Y(n_1176)
);

NAND2x1p5_ASAP7_75t_L g1177 ( 
.A(n_1159),
.B(n_953),
.Y(n_1177)
);

NAND4xp25_ASAP7_75t_L g1178 ( 
.A(n_1142),
.B(n_962),
.C(n_930),
.D(n_993),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1161),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1155),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1147),
.Y(n_1181)
);

NOR2x1_ASAP7_75t_L g1182 ( 
.A(n_1148),
.B(n_962),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1151),
.B(n_962),
.Y(n_1183)
);

NAND2x1p5_ASAP7_75t_L g1184 ( 
.A(n_1163),
.B(n_925),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1158),
.Y(n_1185)
);

XNOR2x1_ASAP7_75t_L g1186 ( 
.A(n_1156),
.B(n_45),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1166),
.B(n_1146),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1185),
.B(n_1170),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_SL g1189 ( 
.A(n_1165),
.B(n_1153),
.C(n_1154),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1174),
.B(n_925),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1179),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1168),
.A2(n_921),
.B(n_927),
.Y(n_1192)
);

AOI221xp5_ASAP7_75t_L g1193 ( 
.A1(n_1180),
.A2(n_993),
.B1(n_990),
.B2(n_930),
.C(n_931),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1176),
.Y(n_1194)
);

NAND3x1_ASAP7_75t_SL g1195 ( 
.A(n_1167),
.B(n_48),
.C(n_49),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1182),
.B(n_971),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1175),
.B(n_971),
.Y(n_1197)
);

INVx1_ASAP7_75t_SL g1198 ( 
.A(n_1172),
.Y(n_1198)
);

NAND3x2_ASAP7_75t_L g1199 ( 
.A(n_1181),
.B(n_921),
.C(n_57),
.Y(n_1199)
);

NOR4xp75_ASAP7_75t_L g1200 ( 
.A(n_1183),
.B(n_51),
.C(n_58),
.D(n_61),
.Y(n_1200)
);

INVxp33_ASAP7_75t_L g1201 ( 
.A(n_1177),
.Y(n_1201)
);

AOI22x1_ASAP7_75t_L g1202 ( 
.A1(n_1191),
.A2(n_1188),
.B1(n_1194),
.B2(n_1198),
.Y(n_1202)
);

OR2x6_ASAP7_75t_L g1203 ( 
.A(n_1187),
.B(n_1169),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1200),
.Y(n_1204)
);

XNOR2x1_ASAP7_75t_L g1205 ( 
.A(n_1199),
.B(n_1186),
.Y(n_1205)
);

OR2x2_ASAP7_75t_L g1206 ( 
.A(n_1201),
.B(n_1171),
.Y(n_1206)
);

AOI22xp5_ASAP7_75t_L g1207 ( 
.A1(n_1189),
.A2(n_1176),
.B1(n_1178),
.B2(n_1173),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1190),
.A2(n_1184),
.B(n_927),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1196),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1195),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1197),
.Y(n_1211)
);

NAND2x1_ASAP7_75t_L g1212 ( 
.A(n_1192),
.B(n_395),
.Y(n_1212)
);

OA211x2_ASAP7_75t_L g1213 ( 
.A1(n_1193),
.A2(n_62),
.B(n_63),
.C(n_65),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1194),
.B(n_68),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1194),
.B(n_70),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1194),
.B(n_72),
.Y(n_1216)
);

OAI22x1_ASAP7_75t_L g1217 ( 
.A1(n_1202),
.A2(n_930),
.B1(n_931),
.B2(n_493),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1206),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1210),
.A2(n_78),
.B1(n_84),
.B2(n_85),
.Y(n_1219)
);

OAI22x1_ASAP7_75t_L g1220 ( 
.A1(n_1207),
.A2(n_493),
.B1(n_914),
.B2(n_910),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1205),
.A2(n_927),
.B1(n_913),
.B2(n_915),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1204),
.A2(n_913),
.B1(n_915),
.B2(n_914),
.Y(n_1222)
);

AOI22x1_ASAP7_75t_SL g1223 ( 
.A1(n_1211),
.A2(n_86),
.B1(n_89),
.B2(n_93),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1203),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1203),
.A2(n_914),
.B1(n_910),
.B2(n_906),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1212),
.A2(n_914),
.B1(n_910),
.B2(n_395),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1224),
.Y(n_1227)
);

AO22x1_ASAP7_75t_L g1228 ( 
.A1(n_1218),
.A2(n_1216),
.B1(n_1215),
.B2(n_1214),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1217),
.A2(n_1209),
.B(n_1208),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1223),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1219),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1226),
.A2(n_1213),
.B(n_395),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1230),
.A2(n_1221),
.B1(n_1219),
.B2(n_1222),
.Y(n_1233)
);

OAI22x1_ASAP7_75t_L g1234 ( 
.A1(n_1227),
.A2(n_1220),
.B1(n_1225),
.B2(n_493),
.Y(n_1234)
);

OAI321xp33_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_910),
.A3(n_906),
.B1(n_104),
.B2(n_108),
.C(n_110),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1231),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1236),
.A2(n_1229),
.B1(n_1228),
.B2(n_906),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1237),
.B(n_1233),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1238),
.Y(n_1239)
);

AOI21xp33_ASAP7_75t_L g1240 ( 
.A1(n_1239),
.A2(n_1234),
.B(n_1235),
.Y(n_1240)
);

AOI221xp5_ASAP7_75t_L g1241 ( 
.A1(n_1240),
.A2(n_96),
.B1(n_99),
.B2(n_114),
.C(n_117),
.Y(n_1241)
);

AOI211xp5_ASAP7_75t_L g1242 ( 
.A1(n_1241),
.A2(n_121),
.B(n_124),
.C(n_128),
.Y(n_1242)
);


endmodule