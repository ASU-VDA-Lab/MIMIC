module fake_jpeg_21371_n_334 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_7),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_16),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_22),
.B(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_48),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_17),
.B1(n_16),
.B2(n_33),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_65),
.B1(n_42),
.B2(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_31),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_61),
.B(n_38),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g101 ( 
.A1(n_64),
.A2(n_50),
.B1(n_23),
.B2(n_35),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_17),
.B1(n_16),
.B2(n_33),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_67),
.A2(n_42),
.B1(n_25),
.B2(n_30),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_84),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_76),
.Y(n_124)
);

AO22x1_ASAP7_75t_SL g72 ( 
.A1(n_61),
.A2(n_42),
.B1(n_41),
.B2(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_40),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_73),
.A2(n_109),
.B1(n_113),
.B2(n_43),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_57),
.A2(n_39),
.B1(n_36),
.B2(n_48),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_74),
.A2(n_86),
.B1(n_91),
.B2(n_104),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_75),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_36),
.B1(n_48),
.B2(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_87),
.B1(n_47),
.B2(n_29),
.Y(n_143)
);

INVx5_ASAP7_75t_SL g78 ( 
.A(n_66),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_78),
.B(n_83),
.Y(n_128)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_51),
.A2(n_37),
.B1(n_42),
.B2(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_80),
.A2(n_99),
.B1(n_115),
.B2(n_43),
.Y(n_130)
);

INVxp67_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_81),
.B(n_100),
.Y(n_145)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_46),
.B1(n_25),
.B2(n_30),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_88),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_96),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_26),
.B1(n_18),
.B2(n_34),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_92),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_19),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_93),
.B(n_95),
.Y(n_132)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_19),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_102),
.Y(n_142)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_51),
.A2(n_50),
.B1(n_49),
.B2(n_26),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_68),
.B(n_18),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_23),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_35),
.B1(n_34),
.B2(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_43),
.B(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_63),
.B(n_38),
.C(n_40),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_47),
.C(n_44),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_60),
.B(n_29),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_63),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_112),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_29),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_114),
.Y(n_153)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_117),
.B(n_138),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_121),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_47),
.B1(n_44),
.B2(n_38),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_143),
.B1(n_146),
.B2(n_109),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_40),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_129),
.A2(n_82),
.B(n_90),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_113),
.A2(n_15),
.B(n_24),
.C(n_12),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_12),
.B(n_10),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_107),
.B(n_87),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_27),
.Y(n_158)
);

AOI32xp33_ASAP7_75t_L g144 ( 
.A1(n_72),
.A2(n_28),
.A3(n_27),
.B1(n_24),
.B2(n_15),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_144),
.B(n_114),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_28),
.B1(n_27),
.B2(n_31),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_101),
.A2(n_24),
.B(n_15),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_105),
.B(n_99),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_31),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_152),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_154),
.A2(n_176),
.B1(n_179),
.B2(n_139),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_108),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_155),
.B(n_158),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_156),
.A2(n_161),
.B(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_116),
.A2(n_78),
.B1(n_80),
.B2(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_159),
.B1(n_175),
.B2(n_122),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_94),
.B1(n_98),
.B2(n_79),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_145),
.B(n_132),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_160),
.B(n_164),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_135),
.B(n_115),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_150),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_165),
.A2(n_129),
.B1(n_121),
.B2(n_131),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_124),
.B(n_83),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_169),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_168),
.Y(n_188)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_135),
.B(n_90),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_112),
.B1(n_85),
.B2(n_10),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_153),
.B1(n_139),
.B2(n_134),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_181),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_141),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_180),
.Y(n_199)
);

OAI22x1_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_3),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_4),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_120),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_190),
.A2(n_202),
.B1(n_203),
.B2(n_218),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_183),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_192),
.B(n_207),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_177),
.B(n_152),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_195),
.B(n_179),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_155),
.B(n_117),
.C(n_126),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_215),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_197),
.A2(n_198),
.B(n_170),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_156),
.A2(n_129),
.B(n_149),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_157),
.A2(n_151),
.B1(n_149),
.B2(n_142),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_119),
.B1(n_153),
.B2(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_133),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_210),
.Y(n_240)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_184),
.B(n_133),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_184),
.B(n_123),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_178),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_212),
.A2(n_216),
.B1(n_159),
.B2(n_175),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_167),
.B(n_125),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_214),
.B(n_182),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_127),
.C(n_123),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_176),
.A2(n_136),
.B1(n_5),
.B2(n_6),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_220),
.A2(n_232),
.B1(n_203),
.B2(n_189),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_187),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_223),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_188),
.B(n_180),
.C(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_237),
.C(n_208),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_190),
.A2(n_170),
.B1(n_178),
.B2(n_154),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_226),
.A2(n_218),
.B1(n_196),
.B2(n_161),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_213),
.B(n_160),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_228),
.B(n_234),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_229),
.B(n_197),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_194),
.B(n_204),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_194),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_231),
.B(n_199),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_172),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_193),
.B(n_163),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_200),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_235),
.B(n_239),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_192),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_217),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_173),
.C(n_164),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_200),
.Y(n_238)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_201),
.Y(n_239)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_207),
.Y(n_241)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_242),
.B(n_243),
.Y(n_262)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_245),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_247),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_206),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_212),
.B1(n_189),
.B2(n_195),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_258),
.B1(n_240),
.B2(n_239),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_251),
.B(n_259),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_198),
.B(n_211),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_229),
.B(n_240),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_236),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_254),
.B(n_261),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_256),
.A2(n_265),
.B1(n_233),
.B2(n_232),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_266),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_210),
.B1(n_191),
.B2(n_215),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_237),
.C(n_225),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_231),
.B(n_199),
.C(n_191),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_246),
.Y(n_280)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_221),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_267),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_272),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_264),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_261),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_243),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_277),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_233),
.C(n_242),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_227),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_261),
.A2(n_220),
.B1(n_226),
.B2(n_227),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_258),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_255),
.A2(n_238),
.B1(n_219),
.B2(n_205),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_219),
.B1(n_265),
.B2(n_241),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_292),
.Y(n_309)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_290),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_272),
.A2(n_252),
.B1(n_263),
.B2(n_259),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_297),
.B1(n_283),
.B2(n_284),
.Y(n_305)
);

INVx11_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_293),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_257),
.C(n_247),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_276),
.C(n_271),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_278),
.A2(n_249),
.B1(n_266),
.B2(n_260),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_169),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_8),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_299),
.A2(n_278),
.B1(n_268),
.B2(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_285),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_305),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_306),
.C(n_298),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_268),
.B(n_275),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_7),
.C(n_8),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_297),
.Y(n_317)
);

INVx6_ASAP7_75t_L g311 ( 
.A(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_313),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_287),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_315),
.B(n_301),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_294),
.C(n_286),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_305),
.C(n_295),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_317),
.B(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_323),
.Y(n_325)
);

AOI21x1_ASAP7_75t_L g321 ( 
.A1(n_314),
.A2(n_292),
.B(n_287),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_322),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_310),
.A2(n_307),
.B1(n_288),
.B2(n_289),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_318),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_324),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_325),
.A2(n_304),
.B(n_323),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_329),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_311),
.B1(n_315),
.B2(n_316),
.Y(n_331)
);

O2A1O1Ixp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_325),
.B(n_312),
.C(n_320),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_332),
.A2(n_312),
.B1(n_295),
.B2(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_293),
.Y(n_334)
);


endmodule