module real_jpeg_6095_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_164;
wire n_48;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_1),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_2),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_4),
.Y(n_170)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_77),
.B1(n_97),
.B2(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_5),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_5),
.A2(n_100),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_6),
.Y(n_155)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_6),
.Y(n_161)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_8),
.A2(n_44),
.B1(n_90),
.B2(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_8),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_93),
.B1(n_145),
.B2(n_147),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_8),
.A2(n_93),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_9),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_9),
.A2(n_125),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_9),
.B(n_80),
.C(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_9),
.B(n_117),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_95),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_11),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_12),
.A2(n_37),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_12),
.A2(n_37),
.B1(n_44),
.B2(n_78),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_174),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_172),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_135),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_16),
.B(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.C(n_101),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_17),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_39),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_18),
.B(n_39),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_29),
.B(n_30),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_20),
.A2(n_31),
.B1(n_163),
.B2(n_169),
.Y(n_162)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_22),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_22),
.Y(n_189)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_22),
.Y(n_221)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_27),
.Y(n_196)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_27),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_28),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_30),
.A2(n_216),
.B(n_222),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_36),
.Y(n_30)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_31),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_31),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_32),
.Y(n_233)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_36),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_38),
.B(n_210),
.Y(n_209)
);

AOI32xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.A3(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_41),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_42),
.Y(n_159)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_46),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_46),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_46),
.Y(n_187)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVxp33_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_56),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_56),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_56),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_60),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_63),
.A2(n_101),
.B1(n_102),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_63),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_89),
.B1(n_94),
.B2(n_96),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_64),
.A2(n_96),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_64),
.A2(n_139),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_65),
.B(n_140),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_79),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_79),
.A2(n_89),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_85),
.B2(n_87),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_92),
.Y(n_119)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_95),
.B(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_123),
.B(n_127),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_117),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B1(n_111),
.B2(n_113),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_117),
.Y(n_134)
);

AO22x2_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_125),
.B(n_126),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_125),
.A2(n_197),
.B(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_134),
.A2(n_144),
.B(n_150),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_142),
.B2(n_171),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_142),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_152),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_162),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.Y(n_154)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_238),
.B(n_243),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_206),
.B(n_237),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_190),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_190),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_179),
.A2(n_185),
.B1(n_186),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_182),
.Y(n_184)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_200),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_191),
.B(n_201),
.C(n_205),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_197),
.B(n_198),
.Y(n_191)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_192),
.Y(n_230)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_227),
.B(n_236),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_214),
.B(n_226),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_212),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_225),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_225),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_234),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_234),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_239),
.B(n_240),
.Y(n_243)
);


endmodule