module fake_netlist_1_12584_n_33 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_8), .A2(n_0), .B1(n_5), .B2(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_3), .B(n_4), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_13), .Y(n_16) );
NOR2xp33_ASAP7_75t_L g17 ( .A(n_11), .B(n_0), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx3_ASAP7_75t_L g19 ( .A(n_16), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
INVxp67_ASAP7_75t_SL g21 ( .A(n_18), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_19), .Y(n_22) );
OR2x2_ASAP7_75t_L g23 ( .A(n_20), .B(n_19), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_22), .B(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_24), .Y(n_27) );
OAI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_20), .B1(n_19), .B2(n_14), .Y(n_28) );
OAI221xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_19), .B1(n_20), .B2(n_15), .C(n_12), .Y(n_29) );
NAND2xp5_ASAP7_75t_SL g30 ( .A(n_28), .B(n_26), .Y(n_30) );
NAND2x1_ASAP7_75t_L g31 ( .A(n_29), .B(n_9), .Y(n_31) );
OAI22xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_19), .B1(n_3), .B2(n_1), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_31), .B1(n_1), .B2(n_10), .Y(n_33) );
endmodule